//#;; Ic23fa9996925b610710d93e28c59a3e2 I10df3d67626099df882920ba6552f16d I93762d802eed04b3e1c59d1d46b35248 Ic9f869114804f0a61ce9b03def9d71f5 I9fc5887c030f7a3e19821ebec457e719
/*I816842ff6f8526885b6ad2d49236bc84*/
////////////////////////////////////////////////////////////////////////////////
//# Copyright (c) 2018 Secantec
//# No Permission to modify and distribute this program
//# even if this copyright message remains unaltered.
//#
//# Author: Secantec 27 April, 2018
//# $Id: $//#
//# Revision History
//#       MM      17  April, 2018    Initial release
//#
////////////////////////////////////////////////////////////////////////////////

// /Ic1111bd512b29e821b120b86446026b8/Id67f249b90615ca158b1258712c3a9fc -Ibea2f3fe6ec7414cdf0bf233abba7ef0 *simv* *csrc* ; If83a0aa1f9ca0f7dd5994445ba7d9e80 I21f66e7dd81ae29064c26b66d9b3e967.I288404204e3d452229308317344a285d -If83a0aa1f9ca0f7dd5994445ba7d9e80 sntc_berlekamp.1.sv > sntc_berlekamp.1.I21f66e7dd81ae29064c26b66d9b3e967.sv ; Id6bfe3ce1bf5714887f4ffbb7b94feab -sverilog -Ie1e1d3d40573127e9ee0480caf1283d6 -Ia823f97963868b5794f5a36e4dbe5dec sntc_berlekamp.1.I21f66e7dd81ae29064c26b66d9b3e967.sv -I2db95e8e1a9267b7a1188556b2013b33 sntc_berlekamp.1.I21f66e7dd81ae29064c26b66d9b3e967.sv.Idc1d71bbb5c4d2a5e936db79ef10c19f

 /*I816842ff6f8526885b6ad2d49236bc84*/

/* I0c35fcd8aa6b70a1e6a2f67174222bd1 Ifaf61c215f3a90fcc150ac387f759daf I54a78636e8c6bd0efb73150b779d5eb5 */

module  sntc_ldpc_decoder#(
// NR_2_0_4/sntc_LDPCparam.sv
parameter MM   = 'h 000a8 ,
// parameter MM =  'h  000a8  , 
parameter NN   = 'h 000d0 ,
// parameter NN =  'h  000d0  , 
parameter cmax = 'h 00017 ,
// parameter cmax =  'h  00017  , 
parameter rmax = 'h 0000a ,
// parameter rmax =  'h  0000a  , 






parameter SUM_NN         = $clog2(NN+1), // 8 : I307afb7f348272492f3cca58ef2f95d8
parameter SUM_MM         = $clog2(MM+1), // 8 : If78618843e4df2223e60ec190987c019
parameter LEN            = MM,
parameter SUM_NN_WDTH    = $clog2(SUM_NN+2),
parameter SUM_MM_WDTH    = $clog2(SUM_MM+2),
`include "NR_2_0_4/sntc_LDPC_dec_param.sv"
`include "NR_2_0_4/flogtanh/GF2_LDPC_flogtanh_param_inc.sv"
  ,
`include "NR_2_0_4/fgallag/GF2_LDPC_fgallag_param_inc.sv"
 ,
parameter MAX_SUM_WDTH_L = 24, //MAX_SUM_WDTH + 3,  // +1 for sign bit for sum0
parameter SGN_MAX_SUM_WDTH = MAX_SUM_WDTH_L - 1, //Ie86b28b55eaf8feb03e24730be892314 sign bit
parameter MAX_SUM_WDTH_L_P1 = 24, //MAX_SUM_WDTH + 3,  // +1 for sign bit for sum0
parameter SGN_MAX_SUM_WDTH_P1 = MAX_SUM_WDTH_L_P1 - 1, //Ie86b28b55eaf8feb03e24730be892314 sign bit
parameter SUM_LEN= $clog2(NN+1),
parameter HAM_LEN= 16
) (

input wire [NN-1:0]                  q0_0,
input wire [NN-1:0]                  q0_1,
output wire [NN-1:0]                 final_y_nr_dec,

input wire [MM-1:0]                  exp_syn,
input wire [31:0]                    percent_probability_int,


input wire  [SUM_LEN-1:0]            HamDist_sum_mm,
input wire  [HAM_LEN-1:0]            HamDist_loop,
input wire  [HAM_LEN-1:0]            HamDist_loop_max,
input wire  [HAM_LEN-1:0]            HamDist_loop_percentage,

output reg                           converged_loops_ended,
output reg                           converged_pass_fail,

output reg                           HamDist_cntr_inc_converged_valid,

input wire  [HAM_LEN-1:0]            HamDist_iir1,
input wire  [HAM_LEN-1:0]            HamDist_iir2,
input wire  [HAM_LEN-1:0]            HamDist_iir3,

input wire                           start_dec,
input wire                           iter_start_int,
/* I0c35fcd8aa6b70a1e6a2f67174222bd1 Ifaf61c215f3a90fcc150ac387f759daf I3bc180bd00be2c60a3a5a68e0dd49503 */
input wire                           clr,
/* I0c35fcd8aa6b70a1e6a2f67174222bd1 I18c0d99dcef0c6b3cc1cadd623fdbf9f I3bc180bd00be2c60a3a5a68e0dd49503 */
input wire                           rstn,
input wire                           clk

);

`ifdef ENCRYPT
`endif

reg [NN-1:0]                     tmp_bit;
reg [12-1:0]                     tmp_bit_msmatch_cnt;
reg [12-1:0]                     I8ff243fdce9dce8c86b33239c193d9bb;
reg [12-1:0]                     fgallag_msmatch_cnt;


wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00016;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00017;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00018;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00019;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00020;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00000_00021;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00016;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00017;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00018;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00019;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00020;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00001_00021;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00016;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00017;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00018;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00019;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00020;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00002_00021;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00016;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00017;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00018;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00019;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00020;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00003_00021;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00016;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00017;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00018;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00019;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00020;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00021;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00004_00022;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00016;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00017;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00018;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00019;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00020;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00021;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00005_00022;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00016;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00017;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00018;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00019;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00020;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00021;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00006_00022;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00016;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00017;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00018;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00019;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00020;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00021;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00007_00022;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00008_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00008_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00008_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00008_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00008_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00008_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00008_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00008_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00008_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00008_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00009_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00009_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00009_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00009_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00009_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00009_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00009_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00009_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00009_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00009_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00010_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00010_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00010_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00010_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00010_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00010_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00010_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00010_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00010_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00010_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00011_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00011_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00011_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00011_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00011_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00011_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00011_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00011_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00011_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00011_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00012_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00012_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00012_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00012_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00012_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00013_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00013_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00013_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00013_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00013_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00014_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00014_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00014_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00014_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00014_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00015_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00015_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00015_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00015_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00015_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00016_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00016_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00016_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00016_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00016_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00017_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00017_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00017_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00017_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00017_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00018_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00018_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00018_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00018_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00018_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00019_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00019_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00019_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00019_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00019_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00020_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00021_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00022_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00023_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00024_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00024_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00024_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00024_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00024_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00024_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00024_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00025_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00025_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00025_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00025_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00025_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00025_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00025_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00026_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00026_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00026_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00026_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00026_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00026_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00026_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00027_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00027_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00027_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00027_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00027_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00027_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00027_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00028_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00029_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00030_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00031_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00032_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00032_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00032_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00032_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00032_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00032_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00033_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00033_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00033_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00033_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00033_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00033_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00034_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00034_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00034_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00034_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00034_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00034_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00035_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00035_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00035_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00035_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00035_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00035_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00036_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00036_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00036_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00036_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00036_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00036_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00036_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00036_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00037_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00037_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00037_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00037_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00037_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00037_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00037_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00037_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00038_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00038_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00038_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00038_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00038_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00038_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00038_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00038_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00039_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00039_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00039_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00039_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00039_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00039_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00039_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00039_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00040_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00040_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00040_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00040_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00040_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00040_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00040_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00040_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00040_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00041_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00041_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00041_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00041_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00041_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00041_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00041_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00041_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00041_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00042_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00042_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00042_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00042_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00042_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00042_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00042_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00042_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00042_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00043_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00043_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00043_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00043_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00043_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00043_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00043_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00043_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00043_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00044_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00045_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00046_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00012;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00013;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00014;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00047_00015;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00048_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00048_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00048_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00048_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00048_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00048_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00048_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00048_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00048_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00049_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00049_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00049_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00049_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00049_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00049_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00049_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00049_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00049_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00050_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00050_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00050_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00050_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00050_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00050_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00050_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00050_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00050_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00051_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00051_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00051_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00051_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00051_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00051_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00051_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00051_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00051_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00052_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00053_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00054_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00001;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00002;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00003;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00004;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00005;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00006;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00007;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00008;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00009;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00010;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00055_00011;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00056_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00057_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00058_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00059_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00060_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00061_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00062_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00063_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00064_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00065_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00066_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00067_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00068_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00069_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00070_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00071_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00072_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00073_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00074_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00075_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00076_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00077_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00078_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00079_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00080_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00081_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00082_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00083_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00084_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00085_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00086_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00087_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00088_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00089_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00090_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00091_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00092_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00093_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00094_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00095_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00096_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00097_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00098_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00099_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00100_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00101_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00102_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00103_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00104_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00105_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00106_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00107_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00108_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00109_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00110_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00111_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00112_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00113_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00114_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00115_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00116_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00117_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00118_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00119_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00120_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00121_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00122_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00123_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00124_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00125_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00126_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00127_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00128_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00129_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00130_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00131_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00132_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00133_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00134_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00135_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00136_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00137_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00138_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00139_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00140_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00141_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00142_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00143_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00144_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00145_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00146_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00147_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00148_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00149_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00150_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00151_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00152_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00153_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00154_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00155_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00156_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00157_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00158_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00159_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00160_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00161_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00162_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00163_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00164_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00165_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00166_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00167_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00168_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00169_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00170_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00171_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00172_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00173_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00174_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00175_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00176_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00177_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00178_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00179_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00180_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00181_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00182_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00183_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00184_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00185_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00186_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00187_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00188_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00189_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00190_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00191_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00192_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00193_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00194_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00195_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00196_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00197_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00198_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00199_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00200_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00201_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00202_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00203_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00204_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00205_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00206_00000;
wire [MAX_SUM_WDTH_L-1:0]        flogtanh_00207_00000;

wire [flogtanh_WDTH -1:0]        Ia67805b59c3011bc4fc5cb1d2996f90d;
wire [MAX_SUM_WDTH_L-1:0]        I0313213a8c479f77e683ce3fa232450c;
wire [MAX_SUM_WDTH_L-1:0]        I5f68368511b59d2e365cc91b806b334e;
wire [flogtanh_WDTH -1:0]        I61fb47b07547e09c746b1fb5d7c8710d;
wire [MAX_SUM_WDTH_L-1:0]        Iad493302f9a77b86d5db79901fcf4a49;
wire [MAX_SUM_WDTH_L-1:0]        I71e4d98dca37256fcc84248a26d703e2;
wire [flogtanh_WDTH -1:0]        Ib2220549c84e87683ccf85798b2bb22f;
wire [MAX_SUM_WDTH_L-1:0]        If50382087360c9884aa683e4e94bcab8;
wire [MAX_SUM_WDTH_L-1:0]        Ib8380902ac4082f834744ddef6d0cc6a;
wire [flogtanh_WDTH -1:0]        I12f063ad18938c2ca008e1165f9119e9;
wire [MAX_SUM_WDTH_L-1:0]        I549ce8de585aa301a4e144342ed29fc6;
wire [MAX_SUM_WDTH_L-1:0]        I9570f8498d95bee230bb3c5e720bb857;
wire [flogtanh_WDTH -1:0]        Iae6b4023f9f2641ca00636181f4fb028;
wire [MAX_SUM_WDTH_L-1:0]        I8af1960c06a98594d58b64b42421b21b;
wire [MAX_SUM_WDTH_L-1:0]        I55c425102db0a6838012a165c0597680;
wire [flogtanh_WDTH -1:0]        Id11b7d1aeb413fd4920ef0e0097fc6c4;
wire [MAX_SUM_WDTH_L-1:0]        I76b14b396d6e5193cc059e68cbd400bd;
wire [MAX_SUM_WDTH_L-1:0]        Ic970a88c435a85d21ed71c6060b8a8e4;
wire [flogtanh_WDTH -1:0]        I3af03d3e0bb7e0e73e034dceda70ff3a;
wire [MAX_SUM_WDTH_L-1:0]        I8c0c834150ae5da887ab265f0f5b2982;
wire [MAX_SUM_WDTH_L-1:0]        Iec8dc328edd6cbaa2d697e05ed222746;
wire [flogtanh_WDTH -1:0]        Iba30a494dc1b66bd2862f82c16017a99;
wire [MAX_SUM_WDTH_L-1:0]        I79934362360a11c365095cfa70a112a1;
wire [MAX_SUM_WDTH_L-1:0]        I16d2084ccfb102c3bafc701872f5ef2d;
wire [flogtanh_WDTH -1:0]        Iefa075dc743d616eca65f76d2c03371c;
wire [MAX_SUM_WDTH_L-1:0]        I65d0cff1828f6d8ba153cadd058a8672;
wire [MAX_SUM_WDTH_L-1:0]        Id680a9affed622577164b3a8380494f5;
wire [flogtanh_WDTH -1:0]        Icc7a632da404a9cda7b8247706391f85;
wire [MAX_SUM_WDTH_L-1:0]        I8a4669217f831b4e42875fea28da24fd;
wire [MAX_SUM_WDTH_L-1:0]        Ifcd68be4bea38622d2d57d3a4e6fc5bb;
wire [flogtanh_WDTH -1:0]        I708c5d8d6d8f7f16c2f348c3b97b906d;
wire [MAX_SUM_WDTH_L-1:0]        Ife6c86fee255f30215fca193d9288a8e;
wire [MAX_SUM_WDTH_L-1:0]        I16deb9107193a3536979e4b5e5654b9c;
wire [flogtanh_WDTH -1:0]        I51ba1e25e01c39a77559089626bafa09;
wire [MAX_SUM_WDTH_L-1:0]        Id8e7f39e4cdcd6d7e1ee2c8f6cce1e46;
wire [MAX_SUM_WDTH_L-1:0]        I28cac65a4db3f708cc90a1b023bfe894;
wire [flogtanh_WDTH -1:0]        I2217e483aaf5124d9beb9baf5037326b;
wire [MAX_SUM_WDTH_L-1:0]        I8c394ac9f9f7e5d96afde79240c0744f;
wire [MAX_SUM_WDTH_L-1:0]        Ie763738b7faf253837e1c45de255cb5e;
wire [flogtanh_WDTH -1:0]        Ib47f8220e7a319e690649f9d6cc9f0cc;
wire [MAX_SUM_WDTH_L-1:0]        I4ab5a06a58aa9b4d293e73712d7a21e7;
wire [MAX_SUM_WDTH_L-1:0]        Icfef12499b53cd84f0aae067f30c17d0;
wire [flogtanh_WDTH -1:0]        Iffc502b536d88d080c59eb3aedd55bd1;
wire [MAX_SUM_WDTH_L-1:0]        Ib09e4bab1aeb88aa15f375adc930c9c8;
wire [MAX_SUM_WDTH_L-1:0]        I0982b8d7f99aceb8871c9c10448f54c5;
wire [flogtanh_WDTH -1:0]        Iaa823b6b13acb376f979dd52683a2231;
wire [MAX_SUM_WDTH_L-1:0]        Ifd56f5082b3fb8406b4c07761d1d61b9;
wire [MAX_SUM_WDTH_L-1:0]        I6c661048307c23c699d4b3636564de0f;
wire [flogtanh_WDTH -1:0]        Ic5f3f371b1ebfe733404b4165fe746dc;
wire [MAX_SUM_WDTH_L-1:0]        I1a7d739018ade49afeb6fbbf0315070d;
wire [MAX_SUM_WDTH_L-1:0]        I786dfcaa131b99c254aaff15bd2c2b6d;
wire [flogtanh_WDTH -1:0]        I021d991730d154218106f00e74bf9d4c;
wire [MAX_SUM_WDTH_L-1:0]        I25c7e7936b9c7b257e5766618159b29d;
wire [MAX_SUM_WDTH_L-1:0]        I2b49d74cb130542f2ca99534e2c513b1;
wire [flogtanh_WDTH -1:0]        I688e5b6520508178afdf85bb2194186d;
wire [MAX_SUM_WDTH_L-1:0]        Ie96ab4759efe3dc122ef44bfc6a90d57;
wire [MAX_SUM_WDTH_L-1:0]        I0f6cb7a5a31d6f2f6178632c0c898bc6;
wire [flogtanh_WDTH -1:0]        I658630f3cf0e86ea86c5fb78b025b0a5;
wire [MAX_SUM_WDTH_L-1:0]        I04dc248d1a638da8d295d8061c0c05af;
wire [MAX_SUM_WDTH_L-1:0]        I03bea609a189246a2375b355df47cf81;
wire [flogtanh_WDTH -1:0]        I8b17f8bae259d829b52aba173bf10b4f;
wire [MAX_SUM_WDTH_L-1:0]        I1260e022c28d8a62d5d93d3d79ddb362;
wire [MAX_SUM_WDTH_L-1:0]        If56555b7cf539750706cf678030ccdb2;
wire [flogtanh_WDTH -1:0]        I944da8181119550916eaf431c7b04c50;
wire [MAX_SUM_WDTH_L-1:0]        Ic77c9c3db51f43825807763f215fd048;
wire [MAX_SUM_WDTH_L-1:0]        I94e89b3a841f9760e3967c97e86d7160;
wire [flogtanh_WDTH -1:0]        I3aa615fa11ad382432ca658ec233f094;
wire [MAX_SUM_WDTH_L-1:0]        Ied24350a62d144813a9469693b4ebdf9;
wire [MAX_SUM_WDTH_L-1:0]        I8cab6f6faf0758f26d1a8851fae43896;
wire [flogtanh_WDTH -1:0]        Ib7c4f77c160ec436e93ca9de75b9fe42;
wire [MAX_SUM_WDTH_L-1:0]        I167e15d8d78007dec518f69156f35a5a;
wire [MAX_SUM_WDTH_L-1:0]        I6ecf7249e6151477fe74a79d0b126b21;
wire [flogtanh_WDTH -1:0]        Ic1e06942b276ee0933dc8b85dec58756;
wire [MAX_SUM_WDTH_L-1:0]        If253f429b0dfc533c619ae813c74142b;
wire [MAX_SUM_WDTH_L-1:0]        I3753b2c4ba8f1bee70def390a96586b0;
wire [flogtanh_WDTH -1:0]        Idd96d8b4e7be386203ec3ed3a81391d9;
wire [MAX_SUM_WDTH_L-1:0]        I2921abdedb74a12af95c937ddaa1b8f4;
wire [MAX_SUM_WDTH_L-1:0]        I9b919f3d4ee3f33506b87bcdaf2d43a3;
wire [flogtanh_WDTH -1:0]        I7df43eec4d78baa1e0680be2715c4495;
wire [MAX_SUM_WDTH_L-1:0]        Ia79f124f8610ca14d7c94a6bcbae2fbc;
wire [MAX_SUM_WDTH_L-1:0]        Ib3be128b6704cc04c61e0fc9814dcf20;
wire [flogtanh_WDTH -1:0]        Ief08536c38479e6bc7fe786cfaf9a10f;
wire [MAX_SUM_WDTH_L-1:0]        I3eb57d0d824ddfa6c789f4bee8a31bc9;
wire [MAX_SUM_WDTH_L-1:0]        If365a3c3ef86dca7c7315b91298c2db8;
wire [flogtanh_WDTH -1:0]        I6ef440b2077563ebbe50dde593c3875a;
wire [MAX_SUM_WDTH_L-1:0]        Ic6b78f30df38e245b28bc68cf70c2ae7;
wire [MAX_SUM_WDTH_L-1:0]        I83560e8d0f8cd37815cca6336fb2208d;
wire [flogtanh_WDTH -1:0]        I20cfad172f0a614687d72d2337ef1003;
wire [MAX_SUM_WDTH_L-1:0]        I68c4a1f713673e5cfd7d40fa2bafb2ec;
wire [MAX_SUM_WDTH_L-1:0]        I099441ae3d3dffe49b18bc578af54dc7;
wire [flogtanh_WDTH -1:0]        Icc6a92285959b25d53b452aed0718c8e;
wire [MAX_SUM_WDTH_L-1:0]        I740a82b22b7a0952639a5d85216e21a3;
wire [MAX_SUM_WDTH_L-1:0]        I58f89947eead94b5054a0fea3520ae33;
wire [flogtanh_WDTH -1:0]        I132c12f1eafbe34bca7b070354bd5f43;
wire [MAX_SUM_WDTH_L-1:0]        I09eae10c74bf18420f829c7f7370e37f;
wire [MAX_SUM_WDTH_L-1:0]        Ibf565bf1803ed43120fa54b80f6f1f29;
wire [flogtanh_WDTH -1:0]        I0f327225758bc82a67a65b8714949a91;
wire [MAX_SUM_WDTH_L-1:0]        I939101803b39bb81310da5f0e6c4a0cb;
wire [MAX_SUM_WDTH_L-1:0]        I619957528c630e7f64924a25127c93fb;
wire [flogtanh_WDTH -1:0]        Ia90d4bc44d3687e912b59e4b6ca02718;
wire [MAX_SUM_WDTH_L-1:0]        Ifea9a62f7fd17b6084afeb9d8ea50e91;
wire [MAX_SUM_WDTH_L-1:0]        If3cc31fd16469339470702045fc6d0da;
wire [flogtanh_WDTH -1:0]        I21c1757545cc2732445c7f978f7247c4;
wire [MAX_SUM_WDTH_L-1:0]        I1b740d99a82724a4bf44d320c0327ad9;
wire [MAX_SUM_WDTH_L-1:0]        I338ccc17dc6158aec0129c8b0c02c429;
wire [flogtanh_WDTH -1:0]        I096fb1aff9431ed667e5d85a6f3726a4;
wire [MAX_SUM_WDTH_L-1:0]        I2f8f6138bbd0bde03c51eafca516e891;
wire [MAX_SUM_WDTH_L-1:0]        I83d71a89f35eb73265ee3e54184e1277;
wire [flogtanh_WDTH -1:0]        Ia69d80cc1f2957ccd79cbd466dea987e;
wire [MAX_SUM_WDTH_L-1:0]        I685c70ac0a2f3404b34c778e92ed5cc7;
wire [MAX_SUM_WDTH_L-1:0]        I7362f08ed4e4ae309dfbfda112c56ad6;
wire [flogtanh_WDTH -1:0]        I2243822bb5cdbca7f2ea942c7b720da8;
wire [MAX_SUM_WDTH_L-1:0]        I759d865a49afde724f226924f73a05eb;
wire [MAX_SUM_WDTH_L-1:0]        I8be4be8471625db0749e6385f87d2dcc;
wire [flogtanh_WDTH -1:0]        Ia77953e90a0cb40984d138c2c209db01;
wire [MAX_SUM_WDTH_L-1:0]        I1917af731dc6b46486e61cf077527e99;
wire [MAX_SUM_WDTH_L-1:0]        I3d6a685a1913bd8be01fddbce1edec2e;
wire [flogtanh_WDTH -1:0]        Id0b03e6dafabbe570f2626f51c9b7121;
wire [MAX_SUM_WDTH_L-1:0]        I3a0a357e2a3b16010a236fa1390680bb;
wire [MAX_SUM_WDTH_L-1:0]        Ifd77e040c5f82790b1d5636a42fca602;
wire [flogtanh_WDTH -1:0]        I5bfac7858439b218179c95c8d8669f17;
wire [MAX_SUM_WDTH_L-1:0]        I8fc051eb8bedd8d14a81345e7f7914c1;
wire [MAX_SUM_WDTH_L-1:0]        Ifbe479e5cab3cba43444bec1e12e72a0;
wire [flogtanh_WDTH -1:0]        I52497c500164c2417f928196ddcdbf84;
wire [MAX_SUM_WDTH_L-1:0]        I9fb6f6ed170f2e914c07ca1973723f74;
wire [MAX_SUM_WDTH_L-1:0]        Ia784f35a5a46837b69eb048dabf84052;
wire [flogtanh_WDTH -1:0]        Ib499dd504da7e433bc1caa258d7e7101;
wire [MAX_SUM_WDTH_L-1:0]        Ib061c8e0e8a973cd42a1861b6f27af43;
wire [MAX_SUM_WDTH_L-1:0]        I8d0f440df332ea96e2d56eec490fbd51;
wire [flogtanh_WDTH -1:0]        I7af88e2be096e488d7269479f935d185;
wire [MAX_SUM_WDTH_L-1:0]        If746d7ebe9868d7bdf6b1884d933fbf8;
wire [MAX_SUM_WDTH_L-1:0]        I8d431a0524241fa54cf6dd1e79de4c74;
wire [flogtanh_WDTH -1:0]        Ief51cc849e0034a9a6b3ff061064ad64;
wire [MAX_SUM_WDTH_L-1:0]        I4c999268e31b807c7ebf1fcb6d0e92e0;
wire [MAX_SUM_WDTH_L-1:0]        If49f97cc0c42b23ce393b534015559a0;
wire [flogtanh_WDTH -1:0]        Ic5f096a42ae6fec933dcaf85faeeda49;
wire [MAX_SUM_WDTH_L-1:0]        If3b89280e3fb4b1526d886740bfcafa4;
wire [MAX_SUM_WDTH_L-1:0]        Ie932a22a7f1fa37087cbc9e8d73efef4;
wire [flogtanh_WDTH -1:0]        Ic9c0a2ce51d641ba7896c2c6911d0f96;
wire [MAX_SUM_WDTH_L-1:0]        I608cd3a092bac42c3f31cea0545ba5b1;
wire [MAX_SUM_WDTH_L-1:0]        I2956687a5fc2fba7149889624ef85647;
wire [flogtanh_WDTH -1:0]        Ia96b3ea2e8395671b3ac674f5a956771;
wire [MAX_SUM_WDTH_L-1:0]        I6c65ea90fb08a2fc85cd61ef7db74ad1;
wire [MAX_SUM_WDTH_L-1:0]        Iebf28886bd39c2540c90e808a9c20d3d;
wire [flogtanh_WDTH -1:0]        Ib81d241e073c97c8c8d1d0abd9a9a64f;
wire [MAX_SUM_WDTH_L-1:0]        Iac77fb31885852fa8f837806ffc0f7b5;
wire [MAX_SUM_WDTH_L-1:0]        I8d4f3e64c8e3b0710a4a6b30d27c8be8;
wire [flogtanh_WDTH -1:0]        I0fc5e49719d7132c7724ee0d406ff93e;
wire [MAX_SUM_WDTH_L-1:0]        I9b000348cc0f46026065aa4af2e5411c;
wire [MAX_SUM_WDTH_L-1:0]        I16e3f3a6802fd206654bb622fa1393fe;
wire [flogtanh_WDTH -1:0]        I4479a0c26d4fa67dee328ecae12d14a4;
wire [MAX_SUM_WDTH_L-1:0]        I9ed46b5dfd0052a65799266c17e3a6e2;
wire [MAX_SUM_WDTH_L-1:0]        I4b5713aee09999592256c407d4b8a95a;
wire [flogtanh_WDTH -1:0]        If5693e079544d04478ec3da9a0ba28d7;
wire [MAX_SUM_WDTH_L-1:0]        Ie1cc391df396e85d4eb86799697a10f5;
wire [MAX_SUM_WDTH_L-1:0]        Ieb1dbb98d5e5bda5b9ce803857f2ca26;
wire [flogtanh_WDTH -1:0]        I701a0ec899c88feef97aeb45fe19e639;
wire [MAX_SUM_WDTH_L-1:0]        I4d60c396c543011e7df7eeb9c9a97137;
wire [MAX_SUM_WDTH_L-1:0]        Ife1c8d014675240a94f1133a78703ed5;
wire [flogtanh_WDTH -1:0]        I6e9d61b111a45e4ea92ff12d33801755;
wire [MAX_SUM_WDTH_L-1:0]        I2ceb0debcadefafcbf0243be5f88f1a0;
wire [MAX_SUM_WDTH_L-1:0]        I94d9412a7b43fa0bd4b9a6d32d313fc7;
wire [flogtanh_WDTH -1:0]        Ief65b0dab6ce1c2fc23cd297a21ac8de;
wire [MAX_SUM_WDTH_L-1:0]        Ieeb8646e8e988cd3e9af56d6aeb23bc1;
wire [MAX_SUM_WDTH_L-1:0]        If13e359e530823319046ce20027445dd;
wire [flogtanh_WDTH -1:0]        Ibb843c4198a06c8e46bc954663c52a28;
wire [MAX_SUM_WDTH_L-1:0]        Ibcadabc2f0ee0f0666a36571bf34a329;
wire [MAX_SUM_WDTH_L-1:0]        I221777352b48c4e228c6637410113854;
wire [flogtanh_WDTH -1:0]        I0c043ef5daa388e93fb3cf6465c217b5;
wire [MAX_SUM_WDTH_L-1:0]        Ic762049ed90ead4c601316c55b05f9fc;
wire [MAX_SUM_WDTH_L-1:0]        I1ee46fec2b82cf8e5142f8e2ac5d9d8a;
wire [flogtanh_WDTH -1:0]        Ife3f07ad3ad5228f10da7020a01e7069;
wire [MAX_SUM_WDTH_L-1:0]        I8c490934df0e2ca56338854686dec05d;
wire [MAX_SUM_WDTH_L-1:0]        Ie45aaf966aa0a94803050b5f43d69e6c;
wire [flogtanh_WDTH -1:0]        I2dacd37cecd93c6e9134cb55ed917d78;
wire [MAX_SUM_WDTH_L-1:0]        I16d19d1f42cf6f0bb1a4f67256aa2d75;
wire [MAX_SUM_WDTH_L-1:0]        I88aedd7f52399f5fd435c3415f2218ca;
wire [flogtanh_WDTH -1:0]        I2419bc316181acd41e29ad005241d812;
wire [MAX_SUM_WDTH_L-1:0]        I5f703ca84e25e921f2d39aae0e1ce236;
wire [MAX_SUM_WDTH_L-1:0]        I7651176b0a74846108fbaabc5cc4900a;
wire [flogtanh_WDTH -1:0]        I35faf0af91f4972ae843883993fc84f4;
wire [MAX_SUM_WDTH_L-1:0]        Ib9de52ec38d9894c339f0d2222da3392;
wire [MAX_SUM_WDTH_L-1:0]        I57ac487adc18165136e9b3c7c50f95ad;
wire [flogtanh_WDTH -1:0]        I4dd2e7b6a685958d7aac77a38354e05f;
wire [MAX_SUM_WDTH_L-1:0]        Ida9dc9ab7922a658c11f40e95543380e;
wire [MAX_SUM_WDTH_L-1:0]        Ic95668328a2121027436f682bac50b9c;
wire [flogtanh_WDTH -1:0]        Ib27460a2e2b13abc54f5ba37f32c8653;
wire [MAX_SUM_WDTH_L-1:0]        I37405a9f44d2155c4e3ecbb317d4b460;
wire [MAX_SUM_WDTH_L-1:0]        I118726375ca9381e45f001965fcefc5b;
wire [flogtanh_WDTH -1:0]        Ia3fa91387788798672eb6199a2eaa389;
wire [MAX_SUM_WDTH_L-1:0]        I47527b41185c39cf18b85e38e3b870de;
wire [MAX_SUM_WDTH_L-1:0]        Ic8d47ff5d6c31601a57df868da78c2d4;
wire [flogtanh_WDTH -1:0]        Ieecd194ccc5698a2ba16efd969cfd621;
wire [MAX_SUM_WDTH_L-1:0]        I995e084dd500652af249f8362d318a97;
wire [MAX_SUM_WDTH_L-1:0]        I7cdc5ada6fc68ee31fd4062e2ff004d3;
wire [flogtanh_WDTH -1:0]        Ifb09fa1840c5a1ddbfc81cda21c11f1e;
wire [MAX_SUM_WDTH_L-1:0]        Id844e291780b20b6e8fd26f9e45fa605;
wire [MAX_SUM_WDTH_L-1:0]        I59547aacdcfde31dc016ec2acbb2f4b4;
wire [flogtanh_WDTH -1:0]        I4ce505ae2025bab3abcf5a44e0ed5034;
wire [MAX_SUM_WDTH_L-1:0]        If47a892c09147f3013077bf8ecf88619;
wire [MAX_SUM_WDTH_L-1:0]        Ia7f53f0cd86055da72c13ac474f052a1;
wire [flogtanh_WDTH -1:0]        Id40a7ca1cde7a70cc13e752e19132808;
wire [MAX_SUM_WDTH_L-1:0]        I41d2ac3db0c604f72f048017b3e8c5cb;
wire [MAX_SUM_WDTH_L-1:0]        I915054f2fbb8b93516d8748a3e3e29e2;
wire [flogtanh_WDTH -1:0]        If7274be2bcc8b2a235c3538db5506d90;
wire [MAX_SUM_WDTH_L-1:0]        I9a54d4d4c2c34cc7807874b016d7c4e2;
wire [MAX_SUM_WDTH_L-1:0]        If257757fa31c2f4cc9ec322e4ecccf83;
wire [flogtanh_WDTH -1:0]        I3e611982ec9ff6437f22e11b2552693a;
wire [MAX_SUM_WDTH_L-1:0]        Ica6b595e3f7d1227e3e90d111d4d7585;
wire [MAX_SUM_WDTH_L-1:0]        If91268e2b84df18785cd6a53e53eb4e9;
wire [flogtanh_WDTH -1:0]        I8fcf0a468234f365c33059e26b9f5821;
wire [MAX_SUM_WDTH_L-1:0]        Icb87e0bd4997398dfb11b851e85e5d50;
wire [MAX_SUM_WDTH_L-1:0]        Ia072f1d679429d3c3180f8eb67fc7dd7;
wire [flogtanh_WDTH -1:0]        I3f80250ee19e8250898f2bcc055c2e5b;
wire [MAX_SUM_WDTH_L-1:0]        Ia1d6b8a34f2f4b6b3495ae760183f9b3;
wire [MAX_SUM_WDTH_L-1:0]        I91a8168d3b087ab3891cd6d479427b95;
wire [flogtanh_WDTH -1:0]        I06b3652935db14aaa057f0cf3cffef66;
wire [MAX_SUM_WDTH_L-1:0]        Ib74566da453368c9846342fdeafcee15;
wire [MAX_SUM_WDTH_L-1:0]        Id1dce8c1542f1279badb381aca3c9b51;
wire [flogtanh_WDTH -1:0]        Ib01d30e88a3a1fcb204246baafeb47c8;
wire [MAX_SUM_WDTH_L-1:0]        If2cfb11905db55514942ab73b9db82aa;
wire [MAX_SUM_WDTH_L-1:0]        I8983f003c30a218543f39f5bbcd9a25c;
wire [flogtanh_WDTH -1:0]        I9f688c58878405d1d2865ddc40659c2b;
wire [MAX_SUM_WDTH_L-1:0]        I60da6c145c6e2723bf4ff550f857a977;
wire [MAX_SUM_WDTH_L-1:0]        Id1b5c33bc63f75561b7cce6fc0981c69;
wire [flogtanh_WDTH -1:0]        Ic9c77123914f831cee5bc4586b6a2a8b;
wire [MAX_SUM_WDTH_L-1:0]        I0f3219717265b7d82d487dea1a63cb62;
wire [MAX_SUM_WDTH_L-1:0]        I003f95fb8f2027efa41a1936e8b53986;
wire [flogtanh_WDTH -1:0]        Ifd42760504e0f106eb9061d9b9a2d18a;
wire [MAX_SUM_WDTH_L-1:0]        I9a4db851c1d6935ab3dfdae9fb85680e;
wire [MAX_SUM_WDTH_L-1:0]        Ie16dc913f571ae73ce03d755077345a9;
wire [flogtanh_WDTH -1:0]        I452794105cca79653f5509dac3794327;
wire [MAX_SUM_WDTH_L-1:0]        I00b3675542777a857263214ae2fa08cd;
wire [MAX_SUM_WDTH_L-1:0]        I86e53eed5b857c439039238bb486067c;
wire [flogtanh_WDTH -1:0]        I33431ed9c549f5525adfa5d45fbc7653;
wire [MAX_SUM_WDTH_L-1:0]        I695c8725ab88beb04f4eeb9d1ec5cbab;
wire [MAX_SUM_WDTH_L-1:0]        I89433799cfa534afd66e8d6b9f1b62b9;
wire [flogtanh_WDTH -1:0]        I4b8b4fd334b176cb449ad0296ebff4c8;
wire [MAX_SUM_WDTH_L-1:0]        I3317b620629d4ed1162708dd76c7fea0;
wire [MAX_SUM_WDTH_L-1:0]        I80f2e8f6743e28e86e4d85b295e2f768;
wire [flogtanh_WDTH -1:0]        I66e7dacba9dbfb14e9a71b9d57229880;
wire [MAX_SUM_WDTH_L-1:0]        I13a81876edd15dc11e22d573b5a33e83;
wire [MAX_SUM_WDTH_L-1:0]        I1391018fb93372ccc2fcc08700e38b65;
wire [flogtanh_WDTH -1:0]        If3a842c52c8c0b2fd24ef265e8cfe330;
wire [MAX_SUM_WDTH_L-1:0]        I64528d9704c63c85bdf41fb3bd66587d;
wire [MAX_SUM_WDTH_L-1:0]        I8fd26d47ecd4cdd08294cf6133468d17;
wire [flogtanh_WDTH -1:0]        I0f3aea4265966e7bc673d3a08ad1c2e4;
wire [MAX_SUM_WDTH_L-1:0]        I38228bcb39eb9ea57aa0bd811e6976a2;
wire [MAX_SUM_WDTH_L-1:0]        I7097c9518bb3351818b96f31ed49c6d3;
wire [flogtanh_WDTH -1:0]        Ia9de78211d220e68835ff757eb75d919;
wire [MAX_SUM_WDTH_L-1:0]        I6ddd4fd20c147c6dff337057753a4ec2;
wire [MAX_SUM_WDTH_L-1:0]        Id683d693cd50645c3d6d657aa1c8bdb2;
wire [flogtanh_WDTH -1:0]        I2c1c31b8bda73b145cdf74b18bc46a4d;
wire [MAX_SUM_WDTH_L-1:0]        I73f34929e9a61c1a6b95107e277fb254;
wire [MAX_SUM_WDTH_L-1:0]        I88bd8012c93dd9e2ed52ea5e9b8b0004;
wire [flogtanh_WDTH -1:0]        I300a84deada851e18835d6af55c5e2a3;
wire [MAX_SUM_WDTH_L-1:0]        Ib078dd08f08128d55534715ee61ea4b8;
wire [MAX_SUM_WDTH_L-1:0]        Ia8d3667adc34b2b50acf7edb970538d8;
wire [flogtanh_WDTH -1:0]        I1fc6745ba86be641dc9bdac044c19519;
wire [MAX_SUM_WDTH_L-1:0]        I3f723dfd62f8ae0057a07480d74562db;
wire [MAX_SUM_WDTH_L-1:0]        I3f0bba472e912f11dea8e788fbc1cb63;
wire [flogtanh_WDTH -1:0]        I2791cc5f69dd0e7f306760048c759af7;
wire [MAX_SUM_WDTH_L-1:0]        Iff7040b14913e56cdf2b36168dcd751e;
wire [MAX_SUM_WDTH_L-1:0]        I6dc671e73b4e9c70cabfdeaac2e5c40b;
wire [flogtanh_WDTH -1:0]        Ie8157cde860052619820431f87e13c83;
wire [MAX_SUM_WDTH_L-1:0]        I72540f5da4495184c7ae5ecc11a96939;
wire [MAX_SUM_WDTH_L-1:0]        Ia6255a136d5f36ea6cba654bd5823850;
wire [flogtanh_WDTH -1:0]        I9059b74a8f3cf2e4905756cc9c71597f;
wire [MAX_SUM_WDTH_L-1:0]        I6174d9699747eed0b49d44974bfb21b0;
wire [MAX_SUM_WDTH_L-1:0]        I2b9584392ef9a7828ff57bd4c522a302;
wire [flogtanh_WDTH -1:0]        I99584eabd3cbd2546c85f474afa6fabb;
wire [MAX_SUM_WDTH_L-1:0]        Iadc74d3274cb3d595c39a8118b2410aa;
wire [MAX_SUM_WDTH_L-1:0]        I6c1235e88ae444a96ea64fd1bfd04d8f;
wire [flogtanh_WDTH -1:0]        I047abade6abf10a65a5b835ac725fa7c;
wire [MAX_SUM_WDTH_L-1:0]        I27493e743da259f4886f63a08165560e;
wire [MAX_SUM_WDTH_L-1:0]        Id09b8242c22851fb960d55222fe733d4;
wire [flogtanh_WDTH -1:0]        Icf7ab1d1113bc44358c56a56fca7caf9;
wire [MAX_SUM_WDTH_L-1:0]        I834b01b9c0bdcbe8cd616ab7dc5e2b91;
wire [MAX_SUM_WDTH_L-1:0]        Ie355fa27abbc41291eaf08f2cf9a6ff7;
wire [flogtanh_WDTH -1:0]        I4d24650be7a1088c2310d93000d6392a;
wire [MAX_SUM_WDTH_L-1:0]        Id69fd2756995da4325484ac912de043a;
wire [MAX_SUM_WDTH_L-1:0]        I566224393f6bb27bfd8b0b0d6b8e53d6;
wire [flogtanh_WDTH -1:0]        Ic3aea8ebb8eab44a92e7d7d950e1a917;
wire [MAX_SUM_WDTH_L-1:0]        Ia23d77f7fcff89e09068364cf3de713a;
wire [MAX_SUM_WDTH_L-1:0]        I8fcad6e7d5ffc9f79eaaf634f6fe8cda;
wire [flogtanh_WDTH -1:0]        I82af0956870500474eac2505bbf15e35;
wire [MAX_SUM_WDTH_L-1:0]        I781d4698facda706103ef8265810eaf6;
wire [MAX_SUM_WDTH_L-1:0]        I6f0f74dcc830fdcb0af9df75a2b722f7;
wire [flogtanh_WDTH -1:0]        I2d8a8efaa0179340bf5d3ebbd4c11831;
wire [MAX_SUM_WDTH_L-1:0]        Ia92f18f2e26ec8ad3578f230d2201274;
wire [MAX_SUM_WDTH_L-1:0]        Idd95fd099dd2b53c46d02f09575b8032;
wire [flogtanh_WDTH -1:0]        I32ff895ff659ec448270067f76e97a90;
wire [MAX_SUM_WDTH_L-1:0]        I1b1a08cc28279b3ffdd544d38704c1ec;
wire [MAX_SUM_WDTH_L-1:0]        I0f277bc88d46a4e6e9f1f2c410b503fd;
wire [flogtanh_WDTH -1:0]        I15a7fd79aeb5eed24b1c7be3d48296e0;
wire [MAX_SUM_WDTH_L-1:0]        Ie12755a265f6a32154b88d22f2037962;
wire [MAX_SUM_WDTH_L-1:0]        I66b92f1de2cf408c3af53b161a6ffa60;
wire [flogtanh_WDTH -1:0]        I12f311f2311e26320a178d6fec95d9d0;
wire [MAX_SUM_WDTH_L-1:0]        I7c27744991b38f3eb69eb9ba2aeb0907;
wire [MAX_SUM_WDTH_L-1:0]        Id28d9545e8d20ac080fbac5e345692da;
wire [flogtanh_WDTH -1:0]        I2b8ce30d1338ad506e4996d2dd1dc11a;
wire [MAX_SUM_WDTH_L-1:0]        I0bbd6f8a9e1e7489421d3b744005b6e6;
wire [MAX_SUM_WDTH_L-1:0]        I4a5cfd6ebd47cda4fa2e06ba9ad6e5b2;
wire [flogtanh_WDTH -1:0]        Ic2b65e7bd42e94f2ad8b6506a6fce7af;
wire [MAX_SUM_WDTH_L-1:0]        Ib9f20533ee570afdeffb0f5279b51d9d;
wire [MAX_SUM_WDTH_L-1:0]        I62bda8dc70e0b5eb38abe094bbe92fc6;
wire [flogtanh_WDTH -1:0]        I0f54a697ea3e2bbf90354c9a6173fb80;
wire [MAX_SUM_WDTH_L-1:0]        I8edc9f2bff969700d0a7e735b533ee9f;
wire [MAX_SUM_WDTH_L-1:0]        I223b05d94c09b095d1988df121aa5e37;
wire [flogtanh_WDTH -1:0]        I6a6c0f8e4399c21285d66ddc0f1f70c0;
wire [MAX_SUM_WDTH_L-1:0]        Id97e6a4e20414f9a23afe284f3e492e3;
wire [MAX_SUM_WDTH_L-1:0]        I5f73e5faf1aca83ee0a415c9ac4a1b9a;
wire [flogtanh_WDTH -1:0]        Ibfcdfc01f09bcff031e359394947efef;
wire [MAX_SUM_WDTH_L-1:0]        If992b3a65059c6e5866c3a03828efb18;
wire [MAX_SUM_WDTH_L-1:0]        I75f9d3a41019dca3044a1c2cf7069662;
wire [flogtanh_WDTH -1:0]        I8efd478f1ae2ea6090774e1ed3bd7b28;
wire [MAX_SUM_WDTH_L-1:0]        Ie7448467fe54559f10316db6ad186b9e;
wire [MAX_SUM_WDTH_L-1:0]        I820fa56328e3919970dd64adb1d4d8e7;
wire [flogtanh_WDTH -1:0]        I502d3210c60c82ca682d8e2168d54be0;
wire [MAX_SUM_WDTH_L-1:0]        I3df80bf9e919f723f65f34362854119f;
wire [MAX_SUM_WDTH_L-1:0]        I05eadf11cdc6c2f2b021e33f2438fa49;
wire [flogtanh_WDTH -1:0]        I337d74c3c773a358a936806f751c1117;
wire [MAX_SUM_WDTH_L-1:0]        Iefe3ca0afaed4b8f7d63ec54591c6cec;
wire [MAX_SUM_WDTH_L-1:0]        I2c487770d606451440eecf358202db32;
wire [flogtanh_WDTH -1:0]        Ia494fdbd70bff11510eb685f3b5d0aae;
wire [MAX_SUM_WDTH_L-1:0]        I1614bb17d0c7c14b07ac4dde98c1fb2a;
wire [MAX_SUM_WDTH_L-1:0]        I082aa8c413d7ef8f054b1c2857cbe39f;
wire [flogtanh_WDTH -1:0]        I547f7a4c3801c1caa4587c9aef397652;
wire [MAX_SUM_WDTH_L-1:0]        Ib1672ae7e0ce15c6fc9eeabc17b8ee97;
wire [MAX_SUM_WDTH_L-1:0]        I420e2c5a8745133f6263a71b458f1e2f;
wire [flogtanh_WDTH -1:0]        I8009d84fd826dd21eb7091744792f4a7;
wire [MAX_SUM_WDTH_L-1:0]        I5efb28aa360b27578d1bbda19162507c;
wire [MAX_SUM_WDTH_L-1:0]        I4b8d520ee88fd39d83a16432e962f731;
wire [flogtanh_WDTH -1:0]        If724b1c92350989910925d275353e544;
wire [MAX_SUM_WDTH_L-1:0]        Ic661342fb3f026ac5b7ca0d5712f572c;
wire [MAX_SUM_WDTH_L-1:0]        Ia3f7f07ddb09ea33218afe14281ac3c6;
wire [flogtanh_WDTH -1:0]        I26f4a180e992f5de04bc047f539bcb48;
wire [MAX_SUM_WDTH_L-1:0]        I84437247e54c9c225c1441622ec111c4;
wire [MAX_SUM_WDTH_L-1:0]        I25aefb53f59a00abe88b9dcf6be6907a;
wire [flogtanh_WDTH -1:0]        I83ca10d71caf5ac98fef3d45d228be8e;
wire [MAX_SUM_WDTH_L-1:0]        I9e0295a7fa30f62feb64d3b4ed2dd4d2;
wire [MAX_SUM_WDTH_L-1:0]        I22c3140a8db02352d2e2a2a11eeba117;
wire [flogtanh_WDTH -1:0]        Ib8407faa17d1e96cd317c65459c4fa71;
wire [MAX_SUM_WDTH_L-1:0]        I1042cc8af315aa7120ea813ae2c5755a;
wire [MAX_SUM_WDTH_L-1:0]        I954dd66f60316803a8f13a39c460a39a;
wire [flogtanh_WDTH -1:0]        I73829d98e5e2f368c4a2020e3d7814be;
wire [MAX_SUM_WDTH_L-1:0]        I1f64264a2c913aeaf4db38f4190cd2dd;
wire [MAX_SUM_WDTH_L-1:0]        I37b3988d699a1ed42923e3fd1584ecc0;
wire [flogtanh_WDTH -1:0]        I9a120c441f8d9ccb617057e042587ba1;
wire [MAX_SUM_WDTH_L-1:0]        I7fa463286e319877ffc9682e696aae89;
wire [MAX_SUM_WDTH_L-1:0]        If79bc5a35cb55036a367efb88c7d5510;
wire [flogtanh_WDTH -1:0]        I8064df8bc33998ad58d460afae699e48;
wire [MAX_SUM_WDTH_L-1:0]        I59c12008dc705cc23fb3093f2ace7c38;
wire [MAX_SUM_WDTH_L-1:0]        Ideab06dc2448a6950cd1a06a0c90c2c6;
wire [flogtanh_WDTH -1:0]        If016e079d3b453444558706ef9073233;
wire [MAX_SUM_WDTH_L-1:0]        I63f19ffd1e2bf12ea726afc806340062;
wire [MAX_SUM_WDTH_L-1:0]        I1d7d7a68fc53b8be89c4637ac8f29380;
wire [flogtanh_WDTH -1:0]        I51cc187d91ee3c480a759104aed41b1b;
wire [MAX_SUM_WDTH_L-1:0]        Ib5408f87beae3f337dfb1e8a75a42a19;
wire [MAX_SUM_WDTH_L-1:0]        Ib34ad1d14978608d1440f59998a31672;
wire [flogtanh_WDTH -1:0]        I4b8068a6a866c2424439b2956245ac8d;
wire [MAX_SUM_WDTH_L-1:0]        I71c3e022d15f1fb4f7b8ffc67c61ab90;
wire [MAX_SUM_WDTH_L-1:0]        Id081512cd113e4d09df0fb13e443d76b;
wire [flogtanh_WDTH -1:0]        I60513d924016bd300559b7a1bea7f521;
wire [MAX_SUM_WDTH_L-1:0]        Ifd815e691b57a5d6f200b40f3953327c;
wire [MAX_SUM_WDTH_L-1:0]        I57a0f8c3710cf8e216d6dc2420f7621c;
wire [flogtanh_WDTH -1:0]        Iec98284ab12724bb63360f29d00f1ecb;
wire [MAX_SUM_WDTH_L-1:0]        I507e631ff186c6a13a989e3bf09dfda0;
wire [MAX_SUM_WDTH_L-1:0]        Iaa164a078c8cdaad694a053c9c1e0313;
wire [flogtanh_WDTH -1:0]        I3e3eba8135eb797d0a5e8ac1feefce0c;
wire [MAX_SUM_WDTH_L-1:0]        I7b0ca33814446a75f820ed3983b8f806;
wire [MAX_SUM_WDTH_L-1:0]        I7eb76b3d17296fdae702d8f820f1428d;
wire [flogtanh_WDTH -1:0]        I6aa98bc7265b8b7c25181a06e75c24c0;
wire [MAX_SUM_WDTH_L-1:0]        Ic0dd354cd8b9e5eb33fffc13285f00e9;
wire [MAX_SUM_WDTH_L-1:0]        I00ecb5e329390023b318a2ceba0df231;
wire [flogtanh_WDTH -1:0]        I47f9c7018999e1cea25feddbe399e6b7;
wire [MAX_SUM_WDTH_L-1:0]        Ifa81b0a7df922d4d85e99dec97ca6c9a;
wire [MAX_SUM_WDTH_L-1:0]        Iea32ebc385c6cfc9212ff37973a0a05d;
wire [flogtanh_WDTH -1:0]        I7224803ba8f0a16a7b2e969fe727bfa1;
wire [MAX_SUM_WDTH_L-1:0]        I91549d4c802e94f6b0400b459b1b5f50;
wire [MAX_SUM_WDTH_L-1:0]        If845af0d620024f04525244753ba5d18;
wire [flogtanh_WDTH -1:0]        I65bc4e0d837f94c4301cb2c87e24969c;
wire [MAX_SUM_WDTH_L-1:0]        Id002cb5fd3d0c0a5c0f7ab1ad6cef723;
wire [MAX_SUM_WDTH_L-1:0]        I08e907b0619bec3ef2cf4cb3779e0794;
wire [flogtanh_WDTH -1:0]        I444f8e61602b8994f7a01f3ebd4ac6ab;
wire [MAX_SUM_WDTH_L-1:0]        I4c6a3ad23b392e26c465731aa152c61c;
wire [MAX_SUM_WDTH_L-1:0]        I68e5b12792a86dda0576742831d3b728;
wire [flogtanh_WDTH -1:0]        I86c51ec7ff965132e195835d21c24881;
wire [MAX_SUM_WDTH_L-1:0]        Iebf49da6d6689a63afa17717ce18e786;
wire [MAX_SUM_WDTH_L-1:0]        I72db05084d30d7c59ba1cb06d3b09400;
wire [flogtanh_WDTH -1:0]        I07aa1b2db5dedc3230dff10534311a56;
wire [MAX_SUM_WDTH_L-1:0]        Id2f4466e93345d0e36e5d72ab56c495c;
wire [MAX_SUM_WDTH_L-1:0]        Ib1f1aef6c0a9291553b62fd555feb2e7;
wire [flogtanh_WDTH -1:0]        Ia8809cc89c377e8b4109cdc8976daa54;
wire [MAX_SUM_WDTH_L-1:0]        I804df90e3a9f73c97b372fc4ecf3dcac;
wire [MAX_SUM_WDTH_L-1:0]        Ib504b808f724ca6032e7c746517cd4fd;
wire [flogtanh_WDTH -1:0]        I7402dc21bfbc0af749dd8fb03c516a50;
wire [MAX_SUM_WDTH_L-1:0]        I52aa4e2bc75f024d35a92ae35bf1b627;
wire [MAX_SUM_WDTH_L-1:0]        Ia47f7fb27f2d965cfd2989569c257356;
wire [flogtanh_WDTH -1:0]        I8ca06f4250a69dde75889f7a6ba3f456;
wire [MAX_SUM_WDTH_L-1:0]        Iefe341800d7dacd81be0ab984ab16f9f;
wire [MAX_SUM_WDTH_L-1:0]        If2b17f9e9186542117f43d0dd342326e;
wire [flogtanh_WDTH -1:0]        Ibab00faeaa6a7be99fa6a239193b92cb;
wire [MAX_SUM_WDTH_L-1:0]        Ic8a0166e91618bc4c689d8b1cb063fdd;
wire [MAX_SUM_WDTH_L-1:0]        I6c4ba0863ab4c8d1a56324a4d89ccbeb;
wire [flogtanh_WDTH -1:0]        I8e44b109466e00487db9dfb7ae225f89;
wire [MAX_SUM_WDTH_L-1:0]        I5097124bb6e421210e0884fcac4f151a;
wire [MAX_SUM_WDTH_L-1:0]        I4dbd1bb8f1641f15e3a4f1e309962811;
wire [flogtanh_WDTH -1:0]        Ib3e38e46bfa9e1bdc032918269223b32;
wire [MAX_SUM_WDTH_L-1:0]        I7334aa542e79be53450da08709732f13;
wire [MAX_SUM_WDTH_L-1:0]        I26781ef851ed43c6f88ff1215cddca6b;
wire [flogtanh_WDTH -1:0]        I659fb1602b9d248940523c14c628ce86;
wire [MAX_SUM_WDTH_L-1:0]        Ice3479ba2aeeccb88630056b7ed6b114;
wire [MAX_SUM_WDTH_L-1:0]        Ia349e1f7c10a63ddccb3f300c73b4572;
wire [flogtanh_WDTH -1:0]        I1a264a901911abed928628d819c162b2;
wire [MAX_SUM_WDTH_L-1:0]        I02dba95d878330150c37c8b9ff4475fe;
wire [MAX_SUM_WDTH_L-1:0]        I50c4e1d3a3f63b93bc36b5141226fb3c;
wire [flogtanh_WDTH -1:0]        I2a53bd293919bc846ab816144b42592a;
wire [MAX_SUM_WDTH_L-1:0]        Iecdd6e6f19312081a8d1ecfdf064e85f;
wire [MAX_SUM_WDTH_L-1:0]        I12334038c2be8634c47869f397503019;
wire [flogtanh_WDTH -1:0]        I35ce9e616a3213f2b4ce0597a47f998c;
wire [MAX_SUM_WDTH_L-1:0]        Iabe6eb7899a7a53e914f54167c877c95;
wire [MAX_SUM_WDTH_L-1:0]        I64692d5168554dfd7ce1c7a046aecf72;
wire [flogtanh_WDTH -1:0]        Ic3f28aa77fc84cb8e2fe43bac7ede253;
wire [MAX_SUM_WDTH_L-1:0]        Ifb841b166cfe3dc103d1cd92e990ea50;
wire [MAX_SUM_WDTH_L-1:0]        Ia4b438844530fff602ea04e72b07db8d;
wire [flogtanh_WDTH -1:0]        I7f91c0e606b4082c6aec2e1f111079c5;
wire [MAX_SUM_WDTH_L-1:0]        I4f9506d81ccabb58d8a95431289c937b;
wire [MAX_SUM_WDTH_L-1:0]        I9574759e112f27778f3645d5d49126b7;
wire [flogtanh_WDTH -1:0]        I8e0d66c2112193437146e0f503623559;
wire [MAX_SUM_WDTH_L-1:0]        Id02f4b88464b945a30c33049c759587f;
wire [MAX_SUM_WDTH_L-1:0]        I2ffb7c2ad09bac694ef13ec41e5de327;
wire [flogtanh_WDTH -1:0]        Iabe6bf045784762fb6b97be3587fd68d;
wire [MAX_SUM_WDTH_L-1:0]        I66f957fcfe83e2474c7fbfa3f6ca7fb0;
wire [MAX_SUM_WDTH_L-1:0]        Ib190f589f4d663dbc0a3c166a8dcf5fa;
wire [flogtanh_WDTH -1:0]        I11f0fd7033065e1695d846f08d11aed5;
wire [MAX_SUM_WDTH_L-1:0]        Icdbc4ac0db607b9959380b85ca6f6a7c;
wire [MAX_SUM_WDTH_L-1:0]        I459c59ac61179d74170db53bf45ba89e;
wire [flogtanh_WDTH -1:0]        Ife1589d99f0764e3757de2a7d8b43008;
wire [MAX_SUM_WDTH_L-1:0]        I889d2418e278c2787154d3bf2a3b3b38;
wire [MAX_SUM_WDTH_L-1:0]        Ie5e432a991aff25577639f1b4ffd594f;
wire [flogtanh_WDTH -1:0]        I7cb3f1f2e7f997b861d6c63d55c0f4ca;
wire [MAX_SUM_WDTH_L-1:0]        I406358d104cee15dd2b7180a1227f7bc;
wire [MAX_SUM_WDTH_L-1:0]        I72064a6a84ff956d76a5aa590bbc05a9;
wire [flogtanh_WDTH -1:0]        Iae2f185d6338026f3e37696327f214df;
wire [MAX_SUM_WDTH_L-1:0]        I94aea1698b59b7a5bee244015bfec001;
wire [MAX_SUM_WDTH_L-1:0]        Iea74ecbac92e1b8f2ec7ad68d10b8e7d;
wire [flogtanh_WDTH -1:0]        I4da8f5b31f5cf7c70bba0cf661d727d8;
wire [MAX_SUM_WDTH_L-1:0]        Ib871d01d3ccfcd49906cd631b4863880;
wire [MAX_SUM_WDTH_L-1:0]        I4f72d0db9fcc358c6fbec9964fbe0bbb;
wire [flogtanh_WDTH -1:0]        I46dd3a6d37d3df901689403a6215b65d;
wire [MAX_SUM_WDTH_L-1:0]        I3e891af010063eeb5059e18c38ca1a9f;
wire [MAX_SUM_WDTH_L-1:0]        Ifd958901d2ea2284f506e04a058012fa;
wire [flogtanh_WDTH -1:0]        I84f43bb1814bdd83a682f7a859cfd611;
wire [MAX_SUM_WDTH_L-1:0]        I58ea1ef4bc81f85225c8028171e8a161;
wire [MAX_SUM_WDTH_L-1:0]        Ie317bbd70b9092b840c0f2713204fb9d;
wire [flogtanh_WDTH -1:0]        I476ea921894e07d3f1d2ff3e7c3b660a;
wire [MAX_SUM_WDTH_L-1:0]        I9f78607e0bc87e0bc7d86de85ffa838a;
wire [MAX_SUM_WDTH_L-1:0]        I2f9e56d570e72714a06c59aa9e4334c0;
wire [flogtanh_WDTH -1:0]        I5cc52764eb8a9961469e1892559ed7ee;
wire [MAX_SUM_WDTH_L-1:0]        I9f1f04e7bc9539c7aa49815fe1515427;
wire [MAX_SUM_WDTH_L-1:0]        I5b53fd45210b92703cb10d583f471ab9;
wire [flogtanh_WDTH -1:0]        I76f68c50b69a7545c0077f5333bfa3e2;
wire [MAX_SUM_WDTH_L-1:0]        Ie07e94ec114e52df8086f86dc5fbc424;
wire [MAX_SUM_WDTH_L-1:0]        I8edbe77bacf1975e014faeee6b861980;
wire [flogtanh_WDTH -1:0]        Id0bd4407ef72994435b3794096636553;
wire [MAX_SUM_WDTH_L-1:0]        Ia048dc6a01575d1733276742fd45bdf5;
wire [MAX_SUM_WDTH_L-1:0]        I174fcbc2ee01fc55edbc8238e5da7f0c;
wire [flogtanh_WDTH -1:0]        I0879a96ba0ef5eb523ae807c40c66a63;
wire [MAX_SUM_WDTH_L-1:0]        Ice646ce92235cc21cb7fc0799053b50a;
wire [MAX_SUM_WDTH_L-1:0]        Id4dc304aef5f35f6ceb91796c278e716;
wire [flogtanh_WDTH -1:0]        I8304ab4dc851d69a7ad7db75ced3eb9e;
wire [MAX_SUM_WDTH_L-1:0]        I6ea1aaf77ecc0369ff33b58439a99d1b;
wire [MAX_SUM_WDTH_L-1:0]        I0cbdfae6f75a639eb591d9c0022f5838;
wire [flogtanh_WDTH -1:0]        I24d773b608ba1ee21855540ee84028da;
wire [MAX_SUM_WDTH_L-1:0]        I93eed7c401e8f511efa112a82b9b9a4f;
wire [MAX_SUM_WDTH_L-1:0]        I088898ee932a96c14f2f0f568f5455b6;
wire [flogtanh_WDTH -1:0]        I9458b9a213600ce0c8c1d54d31c8c5c2;
wire [MAX_SUM_WDTH_L-1:0]        I9ef8088456f239e42f67e7b0ec062c35;
wire [MAX_SUM_WDTH_L-1:0]        Ide0abde3644a4fafb436aa59768d016e;
wire [flogtanh_WDTH -1:0]        Idb6b8e6f2df9b8d96efa93830df86a71;
wire [MAX_SUM_WDTH_L-1:0]        I5529826cbbfacc566e550b2fb6d34200;
wire [MAX_SUM_WDTH_L-1:0]        I08581dc8d42be712cfb36d744f2786e0;
wire [flogtanh_WDTH -1:0]        I0a8fb8a7a28b364bc8cf49b96fdc66a4;
wire [MAX_SUM_WDTH_L-1:0]        I71d41f3f13a20950a8f5e5dace0b9754;
wire [MAX_SUM_WDTH_L-1:0]        I29fb3830a5fc5922f1ec687a38941e97;
wire [flogtanh_WDTH -1:0]        I938f8896ddbf95751aea2b327f5d40f0;
wire [MAX_SUM_WDTH_L-1:0]        Id031c3a3b6acda879451d8d73153bc49;
wire [MAX_SUM_WDTH_L-1:0]        I715d59fb27e519a9b76bdd8b5139a619;
wire [flogtanh_WDTH -1:0]        Ib5b964583d3ef33b47643ca212bc0ada;
wire [MAX_SUM_WDTH_L-1:0]        Idf0dedc8613d3ebf20cfbbe7d4337be9;
wire [MAX_SUM_WDTH_L-1:0]        Ibe6a876a041198a581c95457a7d1fcf8;
wire [flogtanh_WDTH -1:0]        I4bae2a264af742ffe7be73f9a1129efe;
wire [MAX_SUM_WDTH_L-1:0]        I034f9d302ce082349a9d812c9fe46411;
wire [MAX_SUM_WDTH_L-1:0]        Iec078a95a69b081cfb5e987ba9c5a613;
wire [flogtanh_WDTH -1:0]        I041c1a7ef6128c7a1a8f8593d4401f1b;
wire [MAX_SUM_WDTH_L-1:0]        Id1ad76a0501d9ea66134873e99cb211d;
wire [MAX_SUM_WDTH_L-1:0]        I0e8f3f56bce3be1ee4d5f780a2f2a9fe;
wire [flogtanh_WDTH -1:0]        I22c6d2c87ef183ef45805a7c99a7e473;
wire [MAX_SUM_WDTH_L-1:0]        Iec5b39a66a2fd9920c3bed36edb32f02;
wire [MAX_SUM_WDTH_L-1:0]        Ia73cacadbf80c0701a5b5b430c0d5c98;
wire [flogtanh_WDTH -1:0]        I45fef5261954fc84be265f39eb8f9647;
wire [MAX_SUM_WDTH_L-1:0]        Iedeaa45a179ec994bce6b6cc6da0995c;
wire [MAX_SUM_WDTH_L-1:0]        Ic634d26fc09589a29a160e4efb5613a8;
wire [flogtanh_WDTH -1:0]        I3b292cf842e3a7ca9e6d0c4ab345446f;
wire [MAX_SUM_WDTH_L-1:0]        I915031fb071f83ac6eb7357933151d20;
wire [MAX_SUM_WDTH_L-1:0]        Ie1374cac341cf353b1863dae9f544e8b;
wire [flogtanh_WDTH -1:0]        Ie7bff678d39738eb49b599772586210a;
wire [MAX_SUM_WDTH_L-1:0]        If7df947e519a3cd29b42434a9519fbb5;
wire [MAX_SUM_WDTH_L-1:0]        Ia07447985347e9a7f3739bd98867cdfb;
wire [flogtanh_WDTH -1:0]        Ib9d80aab3818d682b54122974fa3a424;
wire [MAX_SUM_WDTH_L-1:0]        I5bac22cea76db3326f60e45aa8ed14c1;
wire [MAX_SUM_WDTH_L-1:0]        I2121318f589878b4a9260625f97de518;
wire [flogtanh_WDTH -1:0]        Iaa05186a94ba0559ab57ced9202ccefb;
wire [MAX_SUM_WDTH_L-1:0]        I2e9180aad8498bc69a9c74af78238e6d;
wire [MAX_SUM_WDTH_L-1:0]        Ibd8424c228f87f85df3da6204edff2b5;
wire [flogtanh_WDTH -1:0]        I506f39735c3743b3705980c73295c035;
wire [MAX_SUM_WDTH_L-1:0]        Id965c3c3f0ab3fc022737b6b577ad6e0;
wire [MAX_SUM_WDTH_L-1:0]        I8a7fb51566bf215af214cd2fb5209974;
wire [flogtanh_WDTH -1:0]        I8f16ead6735608b15b364b9af9b3a22a;
wire [MAX_SUM_WDTH_L-1:0]        I0ecfcdb358eb5e5ed3eb9c5f3f137dd0;
wire [MAX_SUM_WDTH_L-1:0]        I7c0f872988488ac69815d288885dfd2f;
wire [flogtanh_WDTH -1:0]        Id07af023803badc88c51b891cad1b7e5;
wire [MAX_SUM_WDTH_L-1:0]        I094f9bedec7e86f01b6f7e223d13b82f;
wire [MAX_SUM_WDTH_L-1:0]        I3521b10b97b0e74888ce385cfc772945;
wire [flogtanh_WDTH -1:0]        Iecb522fa10764b2c0c044be6c1ca807d;
wire [MAX_SUM_WDTH_L-1:0]        Ib67397a1a44a6cfd5ea04983f1847686;
wire [MAX_SUM_WDTH_L-1:0]        I58f0b81a46549cab8e74ecbc285df23a;
wire [flogtanh_WDTH -1:0]        I58b9a09be96353ba6c18f310e1987742;
wire [MAX_SUM_WDTH_L-1:0]        I2e49a1e612abcd98120c4528eda7c359;
wire [MAX_SUM_WDTH_L-1:0]        I7095040b38bf9d6b5229c11d2a0d7c57;
wire [flogtanh_WDTH -1:0]        I86ced95bff4327e4ab07338663f82029;
wire [MAX_SUM_WDTH_L-1:0]        Id87382649fe91c747a380e2ec4e4cdcd;
wire [MAX_SUM_WDTH_L-1:0]        I675ab6c4fb93b006f3fcafc985fbc405;
wire [flogtanh_WDTH -1:0]        Ia802328754db2d72d6ec8e12a79b2341;
wire [MAX_SUM_WDTH_L-1:0]        Ia29f77138da85cd201325cc411528c73;
wire [MAX_SUM_WDTH_L-1:0]        I239a992ebb62899120a74b1c9e6cc4b4;
wire [flogtanh_WDTH -1:0]        I5b5a9fa50a6e4c7e07017249e5dee137;
wire [MAX_SUM_WDTH_L-1:0]        I29ffc08244342190be5b2adcb968fbea;
wire [MAX_SUM_WDTH_L-1:0]        I927c870d09285dcb47e6d399f319471e;
wire [flogtanh_WDTH -1:0]        I73ef262450353dfcfabe3051ab0006f9;
wire [MAX_SUM_WDTH_L-1:0]        I58ea03377afb90bb2f408efebc0fe7eb;
wire [MAX_SUM_WDTH_L-1:0]        Ie23ed3ee61f468f59f2baf661cb7f85d;
wire [flogtanh_WDTH -1:0]        I959c5d62629333d1d60766a6d935ae4a;
wire [MAX_SUM_WDTH_L-1:0]        I5f7e827df9d731c1ffd418b1ad028b31;
wire [MAX_SUM_WDTH_L-1:0]        I68e58664be09261e5a80d6f8ecdd1b60;
wire [flogtanh_WDTH -1:0]        I659d579ea5b5d24ef0ccbb8160dfe2ae;
wire [MAX_SUM_WDTH_L-1:0]        I6e5a9a96c90b19eb113510e4dc7fe113;
wire [MAX_SUM_WDTH_L-1:0]        Id2808e0f40992c79ead4da7c734e5b79;
wire [flogtanh_WDTH -1:0]        Icae3ba8a84ee6ee051a3caf210f47b51;
wire [MAX_SUM_WDTH_L-1:0]        I9a1438cdffb8de6db7d253106895fd6c;
wire [MAX_SUM_WDTH_L-1:0]        Icb2b390266bff241a688961136db0f51;
wire [flogtanh_WDTH -1:0]        I92a005abe2d27beb2949fe29c0d8bc65;
wire [MAX_SUM_WDTH_L-1:0]        I972c89a3fa5af605d673f846c71f8f57;
wire [MAX_SUM_WDTH_L-1:0]        I54cfd68212d97a2cc8241ef429429453;
wire [flogtanh_WDTH -1:0]        I28fb1164936618d653aa7bf06c03b38f;
wire [MAX_SUM_WDTH_L-1:0]        I6cdde8c6984cc120c0f0a1a0472d50c5;
wire [MAX_SUM_WDTH_L-1:0]        I8d4e3962525c424786ae822a6981a5e6;
wire [flogtanh_WDTH -1:0]        I8720bdf2c91f113b39aa5b6f82421feb;
wire [MAX_SUM_WDTH_L-1:0]        Id2f5757d8a8432506fbffa192a4e0c49;
wire [MAX_SUM_WDTH_L-1:0]        I1a5f22b4e326d1684c0a8c7a7e754ab4;
wire [flogtanh_WDTH -1:0]        I07320e5fb3beddb93ae325a98c5e3782;
wire [MAX_SUM_WDTH_L-1:0]        Iefdb7ed85a168a0fa2e5e93d1d67701e;
wire [MAX_SUM_WDTH_L-1:0]        I8c2e0c83a8204d6b21e0e3e458d56f05;
wire [flogtanh_WDTH -1:0]        Ib8b29bc86ad9c07d7ae5b358f66cb9ba;
wire [MAX_SUM_WDTH_L-1:0]        If1f93a57723e97173a4289a0052945b8;
wire [MAX_SUM_WDTH_L-1:0]        Ie0622ff815747e4a9f368c74787026ec;
wire [flogtanh_WDTH -1:0]        I8e2ed2040f5bf8ea125e5b953cf89300;
wire [MAX_SUM_WDTH_L-1:0]        Ia5ec300f6b8946d5e6ff0cfb22eba4ed;
wire [MAX_SUM_WDTH_L-1:0]        I5ffed139764d90825b9f2eddacd0eddc;
wire [flogtanh_WDTH -1:0]        I4ad3a5b591cd6b13de04897fbbd068ec;
wire [MAX_SUM_WDTH_L-1:0]        I0c27572b0776655756ce831c506bef53;
wire [MAX_SUM_WDTH_L-1:0]        I5a3297f48e1045273db6522744582b05;
wire [flogtanh_WDTH -1:0]        If5208f94e99b0e7ff353c048b55ad7ba;
wire [MAX_SUM_WDTH_L-1:0]        I088d29bd92758302c48dabb469993251;
wire [MAX_SUM_WDTH_L-1:0]        I9858bb2a3cc458aca5bf7eb077ee55dd;
wire [flogtanh_WDTH -1:0]        I66106fad536bb49418e7d09e3f4221ac;
wire [MAX_SUM_WDTH_L-1:0]        Iec3bf0eb952518b856f1596f964e3ae5;
wire [MAX_SUM_WDTH_L-1:0]        I6e7e27bb176196e4493bf9c45ca19719;
wire [flogtanh_WDTH -1:0]        I6af88c096ca3af849bbedb15b2ac7153;
wire [MAX_SUM_WDTH_L-1:0]        I990ed4f7284e44d83197a4cc987c8ff1;
wire [MAX_SUM_WDTH_L-1:0]        I4cff1804df738cbf4f940c775236df9c;
wire [flogtanh_WDTH -1:0]        I15d6e1e431457b954b5f86cd4fb16a77;
wire [MAX_SUM_WDTH_L-1:0]        I7d0dc027656ba91703f0ac89aae218d3;
wire [MAX_SUM_WDTH_L-1:0]        I0c1e22375d5e023c24519901b92eceb5;
wire [flogtanh_WDTH -1:0]        Ifd67d6dec292171610a805560d7cb9a0;
wire [MAX_SUM_WDTH_L-1:0]        I421d6fb792792366ca3d3bf8f8520f56;
wire [MAX_SUM_WDTH_L-1:0]        Ida5b16851dc06534844a0b037d74feb3;
wire [flogtanh_WDTH -1:0]        I681c4ec303ff366746d35234fe5a1ff4;
wire [MAX_SUM_WDTH_L-1:0]        If538078378e360ac004d4b122f75cb42;
wire [MAX_SUM_WDTH_L-1:0]        Iac3cb5b4481687fcf430c8bf52cfb74d;
wire [flogtanh_WDTH -1:0]        I5df2eac3ace0bcef9e48b0850d975cce;
wire [MAX_SUM_WDTH_L-1:0]        Ia144749f2f8b6f0e06f00dd3a6954616;
wire [MAX_SUM_WDTH_L-1:0]        Ia1499972c4995268acd828c1289f353d;
wire [flogtanh_WDTH -1:0]        Icf6f5254160a82036c4ba0367e8f0404;
wire [MAX_SUM_WDTH_L-1:0]        I8dff03248f37764bfe0c2c6b4fcc795f;
wire [MAX_SUM_WDTH_L-1:0]        Ie559401a3a913400dc5e3e5641297fa6;
wire [flogtanh_WDTH -1:0]        If1de12bbb90e49cc1b28eafc2aa551e5;
wire [MAX_SUM_WDTH_L-1:0]        I5d98e3e3fbce58307f7df7fc7d580ac8;
wire [MAX_SUM_WDTH_L-1:0]        Ie0667fbe76244eaec0b155d69dcc9447;
wire [flogtanh_WDTH -1:0]        Ibf9f7f1f6a759af21ac82d6e6ff7df43;
wire [MAX_SUM_WDTH_L-1:0]        Ia47119d76cf6a40b200cd5ecfd4b1409;
wire [MAX_SUM_WDTH_L-1:0]        I1d0f031e8ae9c0335d501d1565118220;
wire [flogtanh_WDTH -1:0]        Ie44bc9632854c4c2077bcec5f46d29ad;
wire [MAX_SUM_WDTH_L-1:0]        Ia10ec5bac071d9ad1941489d7457e0ef;
wire [MAX_SUM_WDTH_L-1:0]        Ie2c801b2de066c3218d7312615b7bfda;
wire [flogtanh_WDTH -1:0]        I97ae894cd928e17cad4c4631aec2c7a0;
wire [MAX_SUM_WDTH_L-1:0]        I048bdd98d2fdac75bdae08d64fa7ef22;
wire [MAX_SUM_WDTH_L-1:0]        I64c4bb0d40d80ec52aab61ce46954f43;
wire [flogtanh_WDTH -1:0]        I500a903104b4b532b3c07d1640e80b55;
wire [MAX_SUM_WDTH_L-1:0]        Ie8075a19a463a00c303aea3814991070;
wire [MAX_SUM_WDTH_L-1:0]        I512f57a40c7c8cb2f040bdde73e44ca3;
wire [flogtanh_WDTH -1:0]        I1d3ae54c8fa3d87a39e3a51018a20727;
wire [MAX_SUM_WDTH_L-1:0]        Iaa6e4f7efa27d63fff2fae677e914cdb;
wire [MAX_SUM_WDTH_L-1:0]        Id60cbf534604e5dba988050ef5abe625;
wire [flogtanh_WDTH -1:0]        I23d3b6da58b66185ddb3c5eae0f68dae;
wire [MAX_SUM_WDTH_L-1:0]        I3eb15cc35c68ee4a5f5294eb5b993259;
wire [MAX_SUM_WDTH_L-1:0]        I37998a91d20db2248ebdd8e661d42f70;
wire [flogtanh_WDTH -1:0]        I88b1352db9aa35be019bc0f345c7131e;
wire [MAX_SUM_WDTH_L-1:0]        I094201803df7b2720fd55ca7a7d870c4;
wire [MAX_SUM_WDTH_L-1:0]        Ib65ff82aff398f6ff7ba711a36f41ee4;
wire [flogtanh_WDTH -1:0]        I1115071c073981f4db4917844fb12a73;
wire [MAX_SUM_WDTH_L-1:0]        I3831fdb5ff3d1597900808314bfa0fd5;
wire [MAX_SUM_WDTH_L-1:0]        I3d1dd8b9c7c6d3913f7ac369ad7e625c;
wire [flogtanh_WDTH -1:0]        Ia9e4e593fd82657c81aeea8fbcd1194b;
wire [MAX_SUM_WDTH_L-1:0]        I092c808c76ddb6c2dc97a552d1f903cf;
wire [MAX_SUM_WDTH_L-1:0]        I097722547450582dc5776bdaff914741;
wire [flogtanh_WDTH -1:0]        I22300986ed621a97a6dac1f3b4d59b8e;
wire [MAX_SUM_WDTH_L-1:0]        I21dc24999451f1e4d8f14813d7d0e58d;
wire [MAX_SUM_WDTH_L-1:0]        Id4a213e494f9c9be0fd1a307e87c756a;
wire [flogtanh_WDTH -1:0]        Icc08ab7c64b40e53278a93f4ae0f9209;
wire [MAX_SUM_WDTH_L-1:0]        I779162012544d75b0d1559145dd29468;
wire [MAX_SUM_WDTH_L-1:0]        I21594c8b0169efd7c2aa6cbc31f4a901;
wire [flogtanh_WDTH -1:0]        I8cc9f5531f2675b3058df110912551b6;
wire [MAX_SUM_WDTH_L-1:0]        I0c0f66943d6470070aeddf77435e28f7;
wire [MAX_SUM_WDTH_L-1:0]        I15022e1b349eee259d3567837283dbf6;
wire [flogtanh_WDTH -1:0]        Icdba6332ba9ea91ffefd690150fba09f;
wire [MAX_SUM_WDTH_L-1:0]        I30faa261a877ce65b3a057bae448bf7f;
wire [MAX_SUM_WDTH_L-1:0]        I1070940dc2ef6e8ee3d1227ec9ff3162;
wire [flogtanh_WDTH -1:0]        Idaef789d04cd5c6291dae88f616460e6;
wire [MAX_SUM_WDTH_L-1:0]        Ia0f7dfeea453a44869ad21670b100db5;
wire [MAX_SUM_WDTH_L-1:0]        I8922cc37cde6ba132f632743113e42af;
wire [flogtanh_WDTH -1:0]        I016cb9c8307b28a7cabf9a91e8da03d6;
wire [MAX_SUM_WDTH_L-1:0]        I32165a54dc2b00d05357e4512ff40ae3;
wire [MAX_SUM_WDTH_L-1:0]        Ia66c399023e500ed67197dcf236f5d42;
wire [flogtanh_WDTH -1:0]        I54517f62dd6f2e7de7d522dfc506383e;
wire [MAX_SUM_WDTH_L-1:0]        I94df0a38de39d37156cb5d84f3c360fc;
wire [MAX_SUM_WDTH_L-1:0]        I1171dc208d5db1024dc3f09a90c78ca0;
wire [flogtanh_WDTH -1:0]        I6b0c1ef6f0a94adaf62425829edf28dd;
wire [MAX_SUM_WDTH_L-1:0]        I85c46907cc9da850a5123a2140d7d75c;
wire [MAX_SUM_WDTH_L-1:0]        Ic28b148967a5b3d05409976fa9001ac8;
wire [flogtanh_WDTH -1:0]        I067ce754b1084de762c33b295f2f47b2;
wire [MAX_SUM_WDTH_L-1:0]        Ib09c12fe109a9604c5877b84c0d09874;
wire [MAX_SUM_WDTH_L-1:0]        I79fe46308b93fbb24245fe1c75edf4a5;
wire [flogtanh_WDTH -1:0]        Ib2fe88cfe23c363993dfcb7722c4fef0;
wire [MAX_SUM_WDTH_L-1:0]        I4e8f05ec6bda855c0625055f7d7d015e;
wire [MAX_SUM_WDTH_L-1:0]        I3bfcd63e92f1949234ab1d2701dbb499;
wire [flogtanh_WDTH -1:0]        I71f836227a1f7f81500a6c980c06f1f7;
wire [MAX_SUM_WDTH_L-1:0]        If3e09ed5717deb2229298308143c32ce;
wire [MAX_SUM_WDTH_L-1:0]        I5e2331edf6e881e9f3a8c47eebda0ac4;
wire [flogtanh_WDTH -1:0]        I6faf34757a61a0b64e61ba059aca33fa;
wire [MAX_SUM_WDTH_L-1:0]        I6cf5a36287d132e0eb71d9006b816cf9;
wire [MAX_SUM_WDTH_L-1:0]        I4b66c202450986ef0df05e979cc8bc7f;
wire [flogtanh_WDTH -1:0]        Ib1821b79b79aadf1486fe1e2df2f297c;
wire [MAX_SUM_WDTH_L-1:0]        If651c14f270904442ab9c299d25a4c16;
wire [MAX_SUM_WDTH_L-1:0]        I737daf208eccf95feb3192897586cdce;
wire [flogtanh_WDTH -1:0]        I84daf07d3f3790c691b9192f7e2018c1;
wire [MAX_SUM_WDTH_L-1:0]        Iebc916f489d40512cab9ad4494fe3405;
wire [MAX_SUM_WDTH_L-1:0]        I29c8133231cfda17668bbe7b692bdfe2;
wire [flogtanh_WDTH -1:0]        Ib4b3ed1f9d1dee96a3ec846424412e2f;
wire [MAX_SUM_WDTH_L-1:0]        I5a0259d2bf5c8a842f607743dcff5851;
wire [MAX_SUM_WDTH_L-1:0]        Id9d56f09595e80d66c2ac300f7d1d972;
wire [flogtanh_WDTH -1:0]        Ibe73f00bb6f1494ede2e6f11f5e7d3f8;
wire [MAX_SUM_WDTH_L-1:0]        Icac9d2c51408fe77883a998c48953a3a;
wire [MAX_SUM_WDTH_L-1:0]        I97e89a2ee18d2688d7c1a640318a1e0d;
wire [flogtanh_WDTH -1:0]        I1542461b996a466d7d3d50bb48ebd690;
wire [MAX_SUM_WDTH_L-1:0]        Icaca84de45cecbfbbc4613ee6b1ebd78;
wire [MAX_SUM_WDTH_L-1:0]        Ife123bf57fe693dabe6aeaa236c4e058;
wire [flogtanh_WDTH -1:0]        If97a5a2c523f51c5881496c5dc8ad11e;
wire [MAX_SUM_WDTH_L-1:0]        I2dc2f2119d90018c1376658e22e66c56;
wire [MAX_SUM_WDTH_L-1:0]        I0c0d844fe3b7d35c1ed6bd7cc4e0dc24;
wire [flogtanh_WDTH -1:0]        Ie19ea558cf2a95ca0c8ae769a809d908;
wire [MAX_SUM_WDTH_L-1:0]        If570315645da3ffaedc01b9bb830e1e5;
wire [MAX_SUM_WDTH_L-1:0]        I2d9632ae6a0f3ba44c3da8f56ba3fedf;
wire [flogtanh_WDTH -1:0]        I6532e6299b8c1fdf7f61b3a44b61c35c;
wire [MAX_SUM_WDTH_L-1:0]        Id5083f0249f7b1bd62260a38e2ad71c9;
wire [MAX_SUM_WDTH_L-1:0]        I38cc7b117c0bcd5e3060cd370d710d7e;
wire [flogtanh_WDTH -1:0]        Ic7102fb8b5df222fff6151e8794bec3c;
wire [MAX_SUM_WDTH_L-1:0]        I7b4308ad008be7a70f2d1d5d7a259479;
wire [MAX_SUM_WDTH_L-1:0]        I793ddbf6a5d026a57ab72984ca19deac;
wire [flogtanh_WDTH -1:0]        I1f97ea0e7bf46382824cbffc3e94e9df;
wire [MAX_SUM_WDTH_L-1:0]        I6b0d8c39fbd70231e5bf5c9b9690476b;
wire [MAX_SUM_WDTH_L-1:0]        I79458089b042e181e37cc44c06d08681;
wire [flogtanh_WDTH -1:0]        I801dfe17655932ad8fe9702cbaad270f;
wire [MAX_SUM_WDTH_L-1:0]        Ie7241b933e5ad5520235b6af19caa8d5;
wire [MAX_SUM_WDTH_L-1:0]        I42460fae0acff25fa2b829e39ddcc4fd;
wire [flogtanh_WDTH -1:0]        Idbd834f0c907b233a8eff58eaca28863;
wire [MAX_SUM_WDTH_L-1:0]        I2a3101f6f107fd42234971ee8ec79ad2;
wire [MAX_SUM_WDTH_L-1:0]        Id3670a6f05d40ab69624544de92b9c64;
wire [flogtanh_WDTH -1:0]        Ic69e0c34630bde15f4172714bc3d92be;
wire [MAX_SUM_WDTH_L-1:0]        Ibc273f3403da77770e246102b6aad94c;
wire [MAX_SUM_WDTH_L-1:0]        I81800fb49855a4fd2737faa07ff15d29;
wire [flogtanh_WDTH -1:0]        I465a735c8e94ddbfdbaeb2a7652e481e;
wire [MAX_SUM_WDTH_L-1:0]        I5a2febf5da7cbbb8bb0aee0830d8122e;
wire [MAX_SUM_WDTH_L-1:0]        Ibfe325e48511372569e0d98d9c4e70e3;
wire [flogtanh_WDTH -1:0]        Id1c6a3f52dd7972f47cbd8103ace643f;
wire [MAX_SUM_WDTH_L-1:0]        I166fdc6588cbe080275b58ccae50fd80;
wire [MAX_SUM_WDTH_L-1:0]        I326660e98f61bb2ced4c23c7bcc9324a;
wire [flogtanh_WDTH -1:0]        I26b9e2d073b20376980662c249bf9d43;
wire [MAX_SUM_WDTH_L-1:0]        Ifde315b0389f701a061b3f765cf35ce7;
wire [MAX_SUM_WDTH_L-1:0]        Ic6fa98631d742b27f252fe7c95caef55;
wire [flogtanh_WDTH -1:0]        Id4cc1b15055941d401ded6ff8b777461;
wire [MAX_SUM_WDTH_L-1:0]        I0df682bffaf274789733b11506a1630f;
wire [MAX_SUM_WDTH_L-1:0]        Iab6d0f72579687407e029c630b107f7d;
wire [flogtanh_WDTH -1:0]        I064bd1f4b7fa40b2cae3ea361edf9167;
wire [MAX_SUM_WDTH_L-1:0]        Ia39290e9e73e101284fb99f7aa472db4;
wire [MAX_SUM_WDTH_L-1:0]        I19eae741ef89baa1a64c403fb29f14f4;
wire [flogtanh_WDTH -1:0]        I4b5aadc25b0ed6811a665b33d6c4ae2a;
wire [MAX_SUM_WDTH_L-1:0]        Ib4f9fe5e96247d914bbdcc12be4044a0;
wire [MAX_SUM_WDTH_L-1:0]        I749b9c345f23aae03c595a2c76126ecb;
wire [flogtanh_WDTH -1:0]        Ic883bcc70572a237ba0e3d465337bc59;
wire [MAX_SUM_WDTH_L-1:0]        I3b06a47b2157c79d4a63dc94865a43c8;
wire [MAX_SUM_WDTH_L-1:0]        Idc77c7d5123717fc2596a51d904c6d82;
wire [flogtanh_WDTH -1:0]        I7181ab1d663b0cbe30861e29fc3f8532;
wire [MAX_SUM_WDTH_L-1:0]        I9f91a577741c480378c018f313c68030;
wire [MAX_SUM_WDTH_L-1:0]        I779da979707d9712c1626d6025f97599;
wire [flogtanh_WDTH -1:0]        Id3fbb6d083344684de89d99c040b2100;
wire [MAX_SUM_WDTH_L-1:0]        I9997a7033ca3806006f2706960325d6d;
wire [MAX_SUM_WDTH_L-1:0]        I97aede8502e443f98938487a5a5c072c;
wire [flogtanh_WDTH -1:0]        Iee8d139aa5a8ae046f5019abecdbc3c4;
wire [MAX_SUM_WDTH_L-1:0]        I0dea21c66fdec2b891938d4cfb4452cd;
wire [MAX_SUM_WDTH_L-1:0]        Ie7820d1a242bc28c19ec32d2c91e47b7;
wire [flogtanh_WDTH -1:0]        Idc0bfe36a3a9b3006a04d5dfc31b8107;
wire [MAX_SUM_WDTH_L-1:0]        Ia6e3665657bc28e92fa4ffb8ddcbc537;
wire [MAX_SUM_WDTH_L-1:0]        I82a14e1ee4723e7d9a13c1f2b8b13691;
wire [flogtanh_WDTH -1:0]        Ia2462ec52aaccc97597d1dfc2e33b7e2;
wire [MAX_SUM_WDTH_L-1:0]        I4097acfa6a9dbc9297745f4891286bd0;
wire [MAX_SUM_WDTH_L-1:0]        I77a94cd9186ca546ca9664942ea3537f;
wire [flogtanh_WDTH -1:0]        I8048bbe27b49b9d248fee919be6dc977;
wire [MAX_SUM_WDTH_L-1:0]        Icef9faf2ee30e443183708bda55cf706;
wire [MAX_SUM_WDTH_L-1:0]        I3c0ddec25c53c166d30eb78d4518840e;
wire [flogtanh_WDTH -1:0]        I838d1cc5e9ca5058c25223ec53d9c34f;
wire [MAX_SUM_WDTH_L-1:0]        I68c9c1da797be9d6d1093884fef3ec3e;
wire [MAX_SUM_WDTH_L-1:0]        I98bbe3b75958f10195dee6460cf2aca6;
wire [flogtanh_WDTH -1:0]        Id9e5147e089e6e52ef2a687d76534f16;
wire [MAX_SUM_WDTH_L-1:0]        Iff7f4a450dee1fe869764249a7a4e612;
wire [MAX_SUM_WDTH_L-1:0]        If6d436031f68ef587750c5c1dfcfffc2;
wire [flogtanh_WDTH -1:0]        Ia043941abbcf10c16f086fe8d61dd456;
wire [MAX_SUM_WDTH_L-1:0]        I323b8c5e397420e5eb3c0872162dc013;
wire [MAX_SUM_WDTH_L-1:0]        I461398638cb8280f1779915298540b00;
wire [flogtanh_WDTH -1:0]        I625ab32380498dfbf9d3290c2053bf3d;
wire [MAX_SUM_WDTH_L-1:0]        Ib62e0c5c630f77706a8bc2ef1409214c;
wire [MAX_SUM_WDTH_L-1:0]        I20c65000bbc10299168af7390776a03c;
wire [flogtanh_WDTH -1:0]        I903f7844e55d1cd6969352490c275c8e;
wire [MAX_SUM_WDTH_L-1:0]        Id51115ce716fdb681e7d5d4cad1fa1c5;
wire [MAX_SUM_WDTH_L-1:0]        Ia840e19ca36795a50ab1a6e6a1729edb;
wire [flogtanh_WDTH -1:0]        Ie5951bc919195ba594fe87375ad41269;
wire [MAX_SUM_WDTH_L-1:0]        Ifbb85fd268ca90f905cbe5587d34cbbb;
wire [MAX_SUM_WDTH_L-1:0]        I7d98d1e5f07fccff5f20eaca6363c700;
wire [flogtanh_WDTH -1:0]        Ieeed8d4eebc0adea7ee0af6a5dbe045c;
wire [MAX_SUM_WDTH_L-1:0]        I7e91bd3d8b70220941a7eb290852b898;
wire [MAX_SUM_WDTH_L-1:0]        I97a75b8625ae2a143cf364790ae77753;
wire [flogtanh_WDTH -1:0]        I266cd5f0a56cd5171da8d59df0042d5d;
wire [MAX_SUM_WDTH_L-1:0]        I366001777963d791fb7811c0fed5f268;
wire [MAX_SUM_WDTH_L-1:0]        Idbea892c8109117f90b453efe8ae25af;
wire [flogtanh_WDTH -1:0]        Ie5a57c603ad520441bc5819c81fb877f;
wire [MAX_SUM_WDTH_L-1:0]        I5db5b227fee3a0a53935d1fd86b1ec77;
wire [MAX_SUM_WDTH_L-1:0]        Icfc1c6d96a3598af73e99a350c387d72;
wire [flogtanh_WDTH -1:0]        I17ac503f4f952f9e2fcdea3f955cc1a9;
wire [MAX_SUM_WDTH_L-1:0]        Id9a0ece818dcc0a00e66ebc35c664c73;
wire [MAX_SUM_WDTH_L-1:0]        I523e9b6f828ec7f166750112f8a3f676;
wire [flogtanh_WDTH -1:0]        Id8b704aada09411d5f5153d088c1c613;
wire [MAX_SUM_WDTH_L-1:0]        I24326227bfacd8f0de4b746ba973242b;
wire [MAX_SUM_WDTH_L-1:0]        I79259217f63b2f6263552c434d0e5c93;
wire [flogtanh_WDTH -1:0]        If64a200b2dac7049b77e5b6bb03b9cc3;
wire [MAX_SUM_WDTH_L-1:0]        Ic96744b0858aea49e052758e4efd4d8a;
wire [MAX_SUM_WDTH_L-1:0]        Ice6db5ba70d3c7499df6723a2df56bfe;
wire [flogtanh_WDTH -1:0]        Iee1b48cae01fe51344b8d662ace9c6f1;
wire [MAX_SUM_WDTH_L-1:0]        I98de4ec4bf1dc2402f1417c2d42a1e2f;
wire [MAX_SUM_WDTH_L-1:0]        I28aa517220bf597cf898660f698ef19d;
wire [flogtanh_WDTH -1:0]        Ic879cd355d61eb021250d62841115a52;
wire [MAX_SUM_WDTH_L-1:0]        I1174526f0aeaaaaa3f10802ea73526f2;
wire [MAX_SUM_WDTH_L-1:0]        I07048dc5cbe24ff72d24902d572face0;
wire [flogtanh_WDTH -1:0]        I46e2d889b9ba7eccad5529200852ca17;
wire [MAX_SUM_WDTH_L-1:0]        Ia49bff02824813d4823f50058348f4e1;
wire [MAX_SUM_WDTH_L-1:0]        Iab3876e5107e3a56b1fafe41e16d9482;
wire [flogtanh_WDTH -1:0]        Ia4e080f13520998be95b64eb883f8e32;
wire [MAX_SUM_WDTH_L-1:0]        I30b6fe386734293d3541f1705a7e2f18;
wire [MAX_SUM_WDTH_L-1:0]        I511a55c2f4d6d3727dff5825597f55a9;
wire [flogtanh_WDTH -1:0]        I2ad2ede07f1ffac643211e88bf8ddbd6;
wire [MAX_SUM_WDTH_L-1:0]        If7541af81460bd2457931a0f435716d8;
wire [MAX_SUM_WDTH_L-1:0]        I2493237a24acdcab8b5bda10e804a5cf;
wire [flogtanh_WDTH -1:0]        I5bc390dc300be5f8bc85f928cca1cd0b;
wire [MAX_SUM_WDTH_L-1:0]        I47cd82d1a6107cbc86188bf1ff4a55a6;
wire [MAX_SUM_WDTH_L-1:0]        I03829256e357ac17c7ca7cae2f980f41;
wire [flogtanh_WDTH -1:0]        I3e7efaed64fd3c276e882ab38109d538;
wire [MAX_SUM_WDTH_L-1:0]        I41f07d0c85ebaf33ef8dd9b96a438df2;
wire [MAX_SUM_WDTH_L-1:0]        Iae32c44b88fe7ddb5d4f19cf8fff3ba6;
wire [flogtanh_WDTH -1:0]        Ib4738fe629dbe40eefed821b40ab93c8;
wire [MAX_SUM_WDTH_L-1:0]        I95a440b3890f6d285bde57a8d879c9aa;
wire [MAX_SUM_WDTH_L-1:0]        I3bdc5ba374f85dc61346e4868c41a6bf;
wire [flogtanh_WDTH -1:0]        I30268ed341753c3ab53b65ad43e94923;
wire [MAX_SUM_WDTH_L-1:0]        I2d3ee951489a62634a7b7332d5fd2450;
wire [MAX_SUM_WDTH_L-1:0]        I557ef77ce931535467a07a8d70145f55;
wire [flogtanh_WDTH -1:0]        I2f10be9cbe2a935475077c0218031a5a;
wire [MAX_SUM_WDTH_L-1:0]        I9f4acc72fd3769c7c300fc36aac958b3;
wire [MAX_SUM_WDTH_L-1:0]        Ib4695d4389db72c5ac7e31809072c290;
wire [flogtanh_WDTH -1:0]        I41d598b80334ab12e5f53b2a6c721517;
wire [MAX_SUM_WDTH_L-1:0]        I4de1d4373a309ecd3278d1891ddce050;
wire [MAX_SUM_WDTH_L-1:0]        Ie81315a3a14a5ef879d8e3f405936365;
wire [flogtanh_WDTH -1:0]        I94b3d895ee69e3ab482ff1aa0798c92a;
wire [MAX_SUM_WDTH_L-1:0]        Iea0a307bacf40b16646458e5e8ea6d9a;
wire [MAX_SUM_WDTH_L-1:0]        Ia7520053a7c4a94437c6a780b03a28a5;
wire [flogtanh_WDTH -1:0]        I24a25d4725db6bcb4732fa21bc861736;
wire [MAX_SUM_WDTH_L-1:0]        Id171f9ecb8da0298882ae2416c2132d3;
wire [MAX_SUM_WDTH_L-1:0]        Ic308a5413f38b96d244cac3b0bc9462c;
wire [flogtanh_WDTH -1:0]        I1877b73e028c908de9dc734b93cbf8bb;
wire [MAX_SUM_WDTH_L-1:0]        Ic10ae3db593c8fb6a2d2a414b131dace;
wire [MAX_SUM_WDTH_L-1:0]        I034fb3850485fae2d1358041a1c41888;
wire [flogtanh_WDTH -1:0]        Ic99b64430e5dfdabe3634fbddeb41b3c;
wire [MAX_SUM_WDTH_L-1:0]        I9dd17bc57b2d75f3e50f2b2243ea6e0b;
wire [MAX_SUM_WDTH_L-1:0]        I0e7079db66c15210046b997f319ece89;
wire [flogtanh_WDTH -1:0]        I3c0ddec6d702a344930fd04f923bb2f1;
wire [MAX_SUM_WDTH_L-1:0]        I69c326b0728bef980588c914c3118d6f;
wire [MAX_SUM_WDTH_L-1:0]        I9a5388f8aa6e9924a309aa8db4c1983b;
wire [flogtanh_WDTH -1:0]        I41829e511abe1ddf9b67f899143db19a;
wire [MAX_SUM_WDTH_L-1:0]        I52e368d1bc43a02ad9418f54b3fe08b8;
wire [MAX_SUM_WDTH_L-1:0]        Ief76663994991118b1899ea4ddf4527d;
wire [flogtanh_WDTH -1:0]        I41961139f5b650e4f4ba5c2eadda6702;
wire [MAX_SUM_WDTH_L-1:0]        I548594daa8f38ff594534dfa4d6238d9;
wire [MAX_SUM_WDTH_L-1:0]        I6fb63ea54e492bdbc6d1145affc683e9;
wire [flogtanh_WDTH -1:0]        I8ef0ac3bf43f16d2edf5a5045b0eb498;
wire [MAX_SUM_WDTH_L-1:0]        I1080d88996caef7f760f64532883ee93;
wire [MAX_SUM_WDTH_L-1:0]        If83ce1cbe3a73472419520c225b288a6;
wire [flogtanh_WDTH -1:0]        I4084e3c9ba635fc4a8d281015bdeb33a;
wire [MAX_SUM_WDTH_L-1:0]        I49f6d04d31956a1134257027fabdb381;
wire [MAX_SUM_WDTH_L-1:0]        Id1df78ab32daf524b77c0431c782f2bf;
wire [flogtanh_WDTH -1:0]        I199a14038a0ff6ac25dab60162f8c6c9;
wire [MAX_SUM_WDTH_L-1:0]        I2aacba8f2c989ba723b7f65c7c009c64;
wire [MAX_SUM_WDTH_L-1:0]        Iff142b88493149045fc0de355b767c16;
wire [flogtanh_WDTH -1:0]        Ic6859263f79d29d5f4896d85367be2bf;
wire [MAX_SUM_WDTH_L-1:0]        If0cf7facd593ca5190b2e20429c1868a;
wire [MAX_SUM_WDTH_L-1:0]        I28c3818247c7c6de11790f6692882b5a;
wire [flogtanh_WDTH -1:0]        If0af3259e321390fffe518318f0f2545;
wire [MAX_SUM_WDTH_L-1:0]        I40d7acfc8d14404d3669e04dbfd61659;
wire [MAX_SUM_WDTH_L-1:0]        Ib451127b69a0a800332a712af77c6d29;
wire [flogtanh_WDTH -1:0]        Icafbf36da24f4db99e0ce4eeca6ca338;
wire [MAX_SUM_WDTH_L-1:0]        I43e5964e737fd1bf55c876d36d1a573d;
wire [MAX_SUM_WDTH_L-1:0]        I3d601db540da359ae4d22f960d3d5af8;
wire [flogtanh_WDTH -1:0]        Ia614303d31afc0ef4f15ec5b43231cd8;
wire [MAX_SUM_WDTH_L-1:0]        I85cc34b35ec9a6e377263bc8307ae9af;
wire [MAX_SUM_WDTH_L-1:0]        I2c1f2476efe593829ade470fe8ec2526;
wire [flogtanh_WDTH -1:0]        I28ff2f86da2016b00bd0c21cbd1b4530;
wire [MAX_SUM_WDTH_L-1:0]        I0bf108b578bd4decc8b7b8d9db13d4a1;
wire [MAX_SUM_WDTH_L-1:0]        I7e685b06df8a8c2ac351fa9f9b76a81d;
wire [flogtanh_WDTH -1:0]        I2b8c969c11b4117c96470f4f6ed6963a;
wire [MAX_SUM_WDTH_L-1:0]        Idcd92c1ab555e9586c17b939903bc6a1;
wire [MAX_SUM_WDTH_L-1:0]        I1338d211b5d2d409bfe0df76d2ca2701;
wire [flogtanh_WDTH -1:0]        Iea563639beb7fcb0291b5dc1410951d1;
wire [MAX_SUM_WDTH_L-1:0]        I45f165607aba91f1026657ea9c265bb7;
wire [MAX_SUM_WDTH_L-1:0]        Ia40dad546d9c852e2fa8942c62a1c1f8;
wire [flogtanh_WDTH -1:0]        Ic1b35046657e23f42199e39343a652a8;
wire [MAX_SUM_WDTH_L-1:0]        If6a9b9c0cff23cab0ac2af86f2eab66a;
wire [MAX_SUM_WDTH_L-1:0]        I0b0dd019d8bd24684403a29aed668b6d;
wire [flogtanh_WDTH -1:0]        Ie7b26120ee77b43574c1ca171d7ec15f;
wire [MAX_SUM_WDTH_L-1:0]        I5f36159573f16b76a28cca6923881ece;
wire [MAX_SUM_WDTH_L-1:0]        I66a304016a9adfd85a2abb6f8fd39afc;
wire [flogtanh_WDTH -1:0]        I2ed61ced1577d905da91d97592006ed5;
wire [MAX_SUM_WDTH_L-1:0]        Icd396e938ee702fab0f788a7a91b90cf;
wire [MAX_SUM_WDTH_L-1:0]        I177be24718c59688752097fe2a4085c4;
wire [flogtanh_WDTH -1:0]        I332dc26a52194745d19c4d8468e42864;
wire [MAX_SUM_WDTH_L-1:0]        I6cee7c45f29f8e1affd935a441d8a0a7;
wire [MAX_SUM_WDTH_L-1:0]        I7e66a42eb7cdb820cd1297c39f0625e8;
wire [flogtanh_WDTH -1:0]        Ibb4fefe05e94e055e86a743c40fb1c5e;
wire [MAX_SUM_WDTH_L-1:0]        I7d389f1dba81f9205521753c52490695;
wire [MAX_SUM_WDTH_L-1:0]        If2021f0735c6c5649ebac0d230fda87c;
wire [flogtanh_WDTH -1:0]        Ia56a76a20d4f11b0e80cbe31820a6977;
wire [MAX_SUM_WDTH_L-1:0]        I759d027d500e4bf950a89c0a49e135c3;
wire [MAX_SUM_WDTH_L-1:0]        Ie1bf5d97b8f679095d2442bbf9f95608;
wire [flogtanh_WDTH -1:0]        I054ebc7f9e3da325ba0c6e329f2ee770;
wire [MAX_SUM_WDTH_L-1:0]        I378871e4d07eabcf01ff30c299f8f054;
wire [MAX_SUM_WDTH_L-1:0]        I632469889d6bb1c268b45fb805467ebd;
wire [flogtanh_WDTH -1:0]        I3361df26cc86ca8be1653d9376d0c8e0;
wire [MAX_SUM_WDTH_L-1:0]        Id346411c557c6ac494ab4913a44c6cf0;
wire [MAX_SUM_WDTH_L-1:0]        Ie230ba3c73808e102eee9e5868595e7c;
wire [flogtanh_WDTH -1:0]        I586fbde80f0130c4a6ead49de11efdd9;
wire [MAX_SUM_WDTH_L-1:0]        I2ed644da3d2a47eef5788a3139de04ac;
wire [MAX_SUM_WDTH_L-1:0]        Ie1e9326e4eee006ec07abb6bb7d269a5;
wire [flogtanh_WDTH -1:0]        Ifa087137c8a6028b13bfa95aba19fc34;
wire [MAX_SUM_WDTH_L-1:0]        I6e90f86b20562e80e2935d1886123672;
wire [MAX_SUM_WDTH_L-1:0]        Ica4ec1647bdb5a3aad6db6b447bd7995;
wire [flogtanh_WDTH -1:0]        I51a3a6c79c488c092394375891775be3;
wire [MAX_SUM_WDTH_L-1:0]        I5c8c09dcb6623c9dee9772f1409ffc98;
wire [MAX_SUM_WDTH_L-1:0]        Ia17295aec0a40c2b46a595dacfede2d5;
wire [flogtanh_WDTH -1:0]        I01a7ebdc760227ee40b85828e28238a9;
wire [MAX_SUM_WDTH_L-1:0]        I6bbd4143192116282eab3d7fbcb544e6;
wire [MAX_SUM_WDTH_L-1:0]        I4c6d3d6fc2d10066a744fdd9405a7902;
wire [flogtanh_WDTH -1:0]        Ib3f9e4c05e363069775e5de9d240b3dc;
wire [MAX_SUM_WDTH_L-1:0]        I5177a497f9d6aae2f1917987542472f0;
wire [MAX_SUM_WDTH_L-1:0]        Ia9c043c5e8873fd13e39cf6bd8136c51;
wire [flogtanh_WDTH -1:0]        I18664482dcc1371fa4b915af96070539;
wire [MAX_SUM_WDTH_L-1:0]        I7cdb256503fb49f4bc9123c0815ea3dd;
wire [MAX_SUM_WDTH_L-1:0]        I2e802c75c6ce34b05943b678ecbfacb1;
wire [flogtanh_WDTH -1:0]        I6a41c6cf78cb25ad1c47550756449002;
wire [MAX_SUM_WDTH_L-1:0]        Ia116be2c3a094f1f5e1d04db21123309;
wire [MAX_SUM_WDTH_L-1:0]        Ieb3f28762410fb40a0c8a8556b4b3ca0;
wire [flogtanh_WDTH -1:0]        Iaf660a97d66e0d7f8e26f65229b7683f;
wire [MAX_SUM_WDTH_L-1:0]        I75175fd0c716e6fbc022cbbd73a9fefd;
wire [MAX_SUM_WDTH_L-1:0]        Ie3e0c0e40c7a67ce7f957e74bd2a895d;
wire [flogtanh_WDTH -1:0]        I7ded197ff64af1bce0e0d85705900a42;
wire [MAX_SUM_WDTH_L-1:0]        I31809c8a10f68b5058f8db1db8d2f714;
wire [MAX_SUM_WDTH_L-1:0]        I491f2373b2df19a4c22e1787ef034179;
wire [flogtanh_WDTH -1:0]        I7c06179d5424165f8a805754834fd98c;
wire [MAX_SUM_WDTH_L-1:0]        I9f4163bac1b52f4282b51e6767085f7f;
wire [MAX_SUM_WDTH_L-1:0]        Ief96603d41b4f670d2bbfa3d3875c903;
wire [flogtanh_WDTH -1:0]        Id364f2a517a0f3109564a025ffd8eec3;
wire [MAX_SUM_WDTH_L-1:0]        Iccc62d273c738111d4ec9adea8c3aec8;
wire [MAX_SUM_WDTH_L-1:0]        I7a029c27d92754041eb6d605837238dd;
wire [flogtanh_WDTH -1:0]        Ie3ea12584ed3e255073776620d778f06;
wire [MAX_SUM_WDTH_L-1:0]        I0c15c6d14710a00728d755472f83d8aa;
wire [MAX_SUM_WDTH_L-1:0]        I00dad36628d2fa923120fdaa79bf0045;
wire [flogtanh_WDTH -1:0]        I38d885c58b4f7333c679b0b5783418df;
wire [MAX_SUM_WDTH_L-1:0]        I5a1afe8d872b05da9e7eb44dd4bafb9f;
wire [MAX_SUM_WDTH_L-1:0]        I3707f68de059df0af5c652fc0478e543;
wire [flogtanh_WDTH -1:0]        I69251440f80eb2e177307aec4cb0111f;
wire [MAX_SUM_WDTH_L-1:0]        If40a1a450ba33087149fb6cdcf1f202e;
wire [MAX_SUM_WDTH_L-1:0]        I94af4b6b9dc11935db54ba872889392d;
wire [flogtanh_WDTH -1:0]        I0a9bcd4a3b79b003b5df8afa0d6b6782;
wire [MAX_SUM_WDTH_L-1:0]        I7079b578409c284713f6b1045c34b659;
wire [MAX_SUM_WDTH_L-1:0]        I38e2dbba093928b874d447362d89b291;
wire [flogtanh_WDTH -1:0]        I36569656996bf98bce33b2d7a4b79def;
wire [MAX_SUM_WDTH_L-1:0]        I336b37e04a2d76a541fcb62871e0c9d4;
wire [MAX_SUM_WDTH_L-1:0]        Ia48f0029e9e76386f3dd70aacd9adbfa;
wire [flogtanh_WDTH -1:0]        I7e408a50d0511909aeb57d5a00535e80;
wire [MAX_SUM_WDTH_L-1:0]        I82325e0f7a4aa9849d619e8b8617c9b8;
wire [MAX_SUM_WDTH_L-1:0]        Ic2b20168744fafbe15037ed7fa83da72;
wire [flogtanh_WDTH -1:0]        Iacc6f48dd92dc515be06a681cc5b56e9;
wire [MAX_SUM_WDTH_L-1:0]        I8bf35575b614154bed06e946d5daf9eb;
wire [MAX_SUM_WDTH_L-1:0]        I62fdc8936121a2707d94cf3bd6e660ac;
wire [flogtanh_WDTH -1:0]        Icafa051878ad3421c31ed2550ea09945;
wire [MAX_SUM_WDTH_L-1:0]        If13d0317f786afef5e7dbbb9d4cd241a;
wire [MAX_SUM_WDTH_L-1:0]        Ia0932b3fd6a5ae6da2bacd2b86ba3a43;
wire [flogtanh_WDTH -1:0]        If4e4f2776b1467e4f03bf15ff5f43c04;
wire [MAX_SUM_WDTH_L-1:0]        I6caaf723f09fdfc7684e94af6fd94d30;
wire [MAX_SUM_WDTH_L-1:0]        I9fce6091885f1bb97d29fb1f543b1a38;
wire [flogtanh_WDTH -1:0]        I9387cd07e38260005bb3e41807d2d794;
wire [MAX_SUM_WDTH_L-1:0]        I3925ce727ac5b2dfff6a5982d034eb80;
wire [MAX_SUM_WDTH_L-1:0]        Ib402cdbfaa9900820b85bd625415c547;
wire [flogtanh_WDTH -1:0]        I8bede290f421e6a05e49244f0d1d3d9b;
wire [MAX_SUM_WDTH_L-1:0]        I3b949d926e8052d319c9262a80951516;
wire [MAX_SUM_WDTH_L-1:0]        I518a2736384c14c02f27bfa3d8ea7aff;
wire [flogtanh_WDTH -1:0]        I6d8c2489fdeb42411f2e12bfa30752d2;
wire [MAX_SUM_WDTH_L-1:0]        I7e8e247667ba53ee311f29a82574c0b7;
wire [MAX_SUM_WDTH_L-1:0]        I847cf7ff866f8a666872c12d6b67b1b1;
wire [flogtanh_WDTH -1:0]        I082715d1b8943faf11d464087542a83e;
wire [MAX_SUM_WDTH_L-1:0]        If6264b63f2c37286744ad61d579d2cc7;
wire [MAX_SUM_WDTH_L-1:0]        I9e45e3d7117ce48cdbfc5db8c0ccfcf4;
wire [flogtanh_WDTH -1:0]        I4de91d9613edc5c4d096b717d9df5de4;
wire [MAX_SUM_WDTH_L-1:0]        I71f47913679ccca9ab806c95c1152182;
wire [MAX_SUM_WDTH_L-1:0]        I380ff8528cdba4026fac3c4eda8b2c52;
wire [flogtanh_WDTH -1:0]        Ifb2a91a74b87c75592cb046b9bfd9c8b;
wire [MAX_SUM_WDTH_L-1:0]        I7b8e7702e50151938e6bb4bcfe59bcad;
wire [MAX_SUM_WDTH_L-1:0]        Iee8f9b0654f6f6797f11cae0947e454e;
wire [flogtanh_WDTH -1:0]        Ie21cffaecd7fe37601dcaef49a0d6cc3;
wire [MAX_SUM_WDTH_L-1:0]        Ic7799445f86a0bb5bed7a74ebe2531fd;
wire [MAX_SUM_WDTH_L-1:0]        Ie3e54a4700d8d0f6478187e06cb6f85d;
wire [flogtanh_WDTH -1:0]        Ia648c9d395ad2727209229807b4224fb;
wire [MAX_SUM_WDTH_L-1:0]        Ic09ec6636c2f6157512550bfe533ac03;
wire [MAX_SUM_WDTH_L-1:0]        I8c0069e8756bcff203ce21ae3170aa42;
wire [flogtanh_WDTH -1:0]        Ib415da845b88e5a8261beaf88b7ec804;
wire [MAX_SUM_WDTH_L-1:0]        I93edc232c5754d21318c71402ba15dad;
wire [MAX_SUM_WDTH_L-1:0]        I856eada207c5006beb8f83f01d5d74c9;
wire [flogtanh_WDTH -1:0]        I6dffcf934a74385aa716db9d7fa29ed1;
wire [MAX_SUM_WDTH_L-1:0]        I8af3fc54adca45e7dbf26e3bd793cd7b;
wire [MAX_SUM_WDTH_L-1:0]        I79a46279070c53678a5af54f661c5821;
wire [flogtanh_WDTH -1:0]        I13383df545ed8620a17a4fc2493cd770;
wire [MAX_SUM_WDTH_L-1:0]        If111e57b5685180f787cc00a5ca98c39;
wire [MAX_SUM_WDTH_L-1:0]        Ica807adc510a2e32580ca77c18ea0b45;
wire [flogtanh_WDTH -1:0]        I87ea43bfae8fad4e4c26741fd2de5b41;
wire [MAX_SUM_WDTH_L-1:0]        I13886c8ae8cffd0b01f2f3ce76fbe755;
wire [MAX_SUM_WDTH_L-1:0]        Ia8094903aed8dd0ce8e9ff459a5287b0;
wire [flogtanh_WDTH -1:0]        I6d2022ba184980b8e5bc5edb4f4b0ff3;
wire [MAX_SUM_WDTH_L-1:0]        Id2e58c1480df3e5cadf231bbd03aaf8e;
wire [MAX_SUM_WDTH_L-1:0]        Ie018f3003c5f124bddd13c359257bf35;
wire [flogtanh_WDTH -1:0]        I68f98b68c9a3836d0c7dc152a2d441da;
wire [MAX_SUM_WDTH_L-1:0]        I5fbf6c0b386eb14a493c94824ba51dea;
wire [MAX_SUM_WDTH_L-1:0]        Ice18bceb10fec484ffc96155e14c4974;
wire [flogtanh_WDTH -1:0]        I2dc3cec85c37aa943f01df545f952e05;
wire [MAX_SUM_WDTH_L-1:0]        I8a77a7011da9a8d0a14e561b73d7df86;
wire [MAX_SUM_WDTH_L-1:0]        Ib484aa64b795f7e36198b800f302164f;
wire [flogtanh_WDTH -1:0]        Ieed49c262f87c86b30d94e9842525ab0;
wire [MAX_SUM_WDTH_L-1:0]        Ifa70dba64cfba1806028839643ea900b;
wire [MAX_SUM_WDTH_L-1:0]        Icdb143a4ce96029c2441758bf2edd7b0;
wire [flogtanh_WDTH -1:0]        Ib9ab475010c98fc4e06df5c98944387a;
wire [MAX_SUM_WDTH_L-1:0]        If81b9c6cecfb4f03c642cf8ad899833a;
wire [MAX_SUM_WDTH_L-1:0]        I3a76f70ca3bfbcacc6f3342aa71f1912;
wire [flogtanh_WDTH -1:0]        If7c8bdd5bae4a1bffd4bd2c8015bb738;
wire [MAX_SUM_WDTH_L-1:0]        Ia515c4910fdd7af0fbf81e2094be54e0;
wire [MAX_SUM_WDTH_L-1:0]        I9470c7ab9634c01bb832c9e4ff5496bf;
wire [flogtanh_WDTH -1:0]        I6463249144cd032e1c5af9e2987254b3;
wire [MAX_SUM_WDTH_L-1:0]        Ic110a8375139cd038f6fad5631ff6df6;
wire [MAX_SUM_WDTH_L-1:0]        I218ee96418a4f5d734d3d71685bc09c7;
wire [flogtanh_WDTH -1:0]        I5f9e468fc1bc199574d719d866d52dfc;
wire [MAX_SUM_WDTH_L-1:0]        I5b1da643c42d2bf15855112416b6ee01;
wire [MAX_SUM_WDTH_L-1:0]        I924514226fdb5bac110a2650bcb2e85f;
wire [flogtanh_WDTH -1:0]        Ie69f792c606c3162052840dec732ef99;
wire [MAX_SUM_WDTH_L-1:0]        Iefe55f571684afc7c5257ae145de8594;
wire [MAX_SUM_WDTH_L-1:0]        Idc57f37015a48393608e2b026bc7065c;
wire [flogtanh_WDTH -1:0]        If874254c3c6813ff0d5184b574cb613d;
wire [MAX_SUM_WDTH_L-1:0]        I7195c3cd02b5b61f50217c41cd409cf6;
wire [MAX_SUM_WDTH_L-1:0]        I41af7e4c97fc04154fe6de66b82499f5;
wire [flogtanh_WDTH -1:0]        I90969c917df8480d379afef834c1a253;
wire [MAX_SUM_WDTH_L-1:0]        I39f71f309736112e18565c8a18bc594a;
wire [MAX_SUM_WDTH_L-1:0]        I972bee4216f8e532e8fa4bd25fbb9c57;
wire [flogtanh_WDTH -1:0]        I07280ae3417855f994980fbb95696fc6;
wire [MAX_SUM_WDTH_L-1:0]        I4fb6ab2aea28cb0776f52fc291782a27;
wire [MAX_SUM_WDTH_L-1:0]        Ib303ea0240e7ab5f000dd10e975b2274;
wire [flogtanh_WDTH -1:0]        I852c62fffff0fd7bf06939d75fada3eb;
wire [MAX_SUM_WDTH_L-1:0]        I85d1c9d05f286204503b33dc9417c3f4;
wire [MAX_SUM_WDTH_L-1:0]        I5971253546899e9a82f387d5eabcc7b3;
wire [flogtanh_WDTH -1:0]        I9e0a2da5a82f1b509bd502554f4760aa;
wire [MAX_SUM_WDTH_L-1:0]        I8827c931edb38391e37eca5443c0f26a;
wire [MAX_SUM_WDTH_L-1:0]        I1fc36e6f738fab96df356979e1e3a612;
wire [flogtanh_WDTH -1:0]        I6293c2b405087f14b42b423336f6990c;
wire [MAX_SUM_WDTH_L-1:0]        I495c79f2d8ec79a2f03613e0b64bde0e;
wire [MAX_SUM_WDTH_L-1:0]        Ie2d8c84d8c9a4c8f637068a2ae39fdde;
wire [flogtanh_WDTH -1:0]        I70e8d96970e69bc828a6aea5ade3bdd1;
wire [MAX_SUM_WDTH_L-1:0]        I954c51f604d6b8e7557797dd06aec9b7;
wire [MAX_SUM_WDTH_L-1:0]        I114c595caa67a3f777f087a634130a6d;
wire [flogtanh_WDTH -1:0]        I0380003f741eedb994793c2cb7e6c5c3;
wire [MAX_SUM_WDTH_L-1:0]        Icd91fad15b5b5844144ac5c34218955f;
wire [MAX_SUM_WDTH_L-1:0]        Idad14b6383b9af54eb35e72ff3d10035;
wire [flogtanh_WDTH -1:0]        Ia884fcfa49cfe0b404bf49b99d7381aa;
wire [MAX_SUM_WDTH_L-1:0]        I4caf7dc4da499ea51928aa11326e0eae;
wire [MAX_SUM_WDTH_L-1:0]        I46e9c76b19ed1ff21f102efe6ee5c732;
wire [flogtanh_WDTH -1:0]        Ie4ecd4c122ea5b478f3d7d2d632b8bf4;
wire [MAX_SUM_WDTH_L-1:0]        I5461e1657c752f83cca50253e1db6772;
wire [MAX_SUM_WDTH_L-1:0]        Ic75b8bbb1b80001ec188a0cd25623420;
wire [flogtanh_WDTH -1:0]        I82e534ecaabf5af6a9b6a567b862800a;
wire [MAX_SUM_WDTH_L-1:0]        Ib184e1d3a451b69a5206cf83e0b787f6;
wire [MAX_SUM_WDTH_L-1:0]        Idc7df6877bdb7e7d392307d78183d31c;
wire [flogtanh_WDTH -1:0]        I1c9684b45467216a18a3a0d93b555b60;
wire [MAX_SUM_WDTH_L-1:0]        If6d01c60d560e37c2676de16f9c10d20;
wire [MAX_SUM_WDTH_L-1:0]        Ib8b95ece5da3877b261a06e6d0571921;
wire [flogtanh_WDTH -1:0]        Ice212c509101d6d41b52ea0cb85dacc0;
wire [MAX_SUM_WDTH_L-1:0]        Ic191abac086c847828546b8feea4fb23;
wire [MAX_SUM_WDTH_L-1:0]        Ic99654bf4833c9132912eeb4c0dc92fa;
wire [flogtanh_WDTH -1:0]        I37ee7a2fab22cf8e6452fb408b849595;
wire [MAX_SUM_WDTH_L-1:0]        I08c8ec03b53121517a27ff7fa143e5cb;
wire [MAX_SUM_WDTH_L-1:0]        I2461055ef9b1aa2ffca0f5cac3300e71;
wire [flogtanh_WDTH -1:0]        I0ec18ade132eede6849e0607af608726;
wire [MAX_SUM_WDTH_L-1:0]        I52362ce3dd44269cdce0797f54886036;
wire [MAX_SUM_WDTH_L-1:0]        I2bc3ffbe5b42b0833206437d3863278e;
wire [flogtanh_WDTH -1:0]        I4651eab27cb766a1792f9564bcb2764a;
wire [MAX_SUM_WDTH_L-1:0]        Ib36da02cb5325af53c1cebe6e20b9468;
wire [MAX_SUM_WDTH_L-1:0]        Id5e02d4c48fa6c3b0d45a9e66f09448f;
wire [flogtanh_WDTH -1:0]        Ibbdbc4e4fc2ee018a0e7a4da29e85b56;
wire [MAX_SUM_WDTH_L-1:0]        I8be5606ad0efbff7ccb552566592ef15;
wire [MAX_SUM_WDTH_L-1:0]        I40e99289d5762e77a3766eb8251eef00;
wire [flogtanh_WDTH -1:0]        Ic67b9e090d6815b2a745bdc4983f9c69;
wire [MAX_SUM_WDTH_L-1:0]        Ie70af982f7791be92f896afe027c8832;
wire [MAX_SUM_WDTH_L-1:0]        I20beb3fdbe91936f74a200cd8ec9817b;
wire [flogtanh_WDTH -1:0]        I8327267045af5da02c066a5eab25f13a;
wire [MAX_SUM_WDTH_L-1:0]        I93ed828faec287b2295a3f860d818fbe;
wire [MAX_SUM_WDTH_L-1:0]        Id435b68afb53bef4afc7b70a9512e955;
wire [flogtanh_WDTH -1:0]        Id91ef7e27c689cdf5ce50d705017e40e;
wire [MAX_SUM_WDTH_L-1:0]        Ifea8cb28a2e829628ceae6126c81eb1f;
wire [MAX_SUM_WDTH_L-1:0]        I0cf5cb4cd472502b84dbf6fe1af0be78;
wire [flogtanh_WDTH -1:0]        I60498760f3c03cf92ceeb99c5096fe54;
wire [MAX_SUM_WDTH_L-1:0]        Idd12f95ce2cb0eb33dbbb09a235c3ca0;
wire [MAX_SUM_WDTH_L-1:0]        Iacf6340a29a5592b61ea875304a2de48;
wire [flogtanh_WDTH -1:0]        I63169dbc533400e0db5e37a8ebeca1aa;
wire [MAX_SUM_WDTH_L-1:0]        I2cfcf8d0beaa4aceb9182c835352b210;
wire [MAX_SUM_WDTH_L-1:0]        I5dfc71255cba279420b7545df4d35c40;
wire [flogtanh_WDTH -1:0]        I150f11a565ad39c59d8f9e4c94d397e2;
wire [MAX_SUM_WDTH_L-1:0]        I7bcc86543042aa717d956b83566442d2;
wire [MAX_SUM_WDTH_L-1:0]        Ibadcb205c7e9a0f3345cac7eb41b5985;
wire [flogtanh_WDTH -1:0]        Icadb816a238ba165425e5a30bd0bb8e6;
wire [MAX_SUM_WDTH_L-1:0]        I4ae99bdc1aca92e0c7ebec69455db910;
wire [MAX_SUM_WDTH_L-1:0]        I762b2abb876381eff6de97cef0798405;
wire [flogtanh_WDTH -1:0]        I3b55785b9625ac53f6c00ba5a10a481b;
wire [MAX_SUM_WDTH_L-1:0]        I612ab97c8ff0b0000f5321336aa31481;
wire [MAX_SUM_WDTH_L-1:0]        Ib3e7633767b6e09e4ee54f6feaddd31e;
wire [flogtanh_WDTH -1:0]        If7317c81c9b6503386cab33fa812e80e;
wire [MAX_SUM_WDTH_L-1:0]        I837c986c9a0267bcb434c774c307542e;
wire [MAX_SUM_WDTH_L-1:0]        I3f193e9c265c1dfaeada63d59db5b79f;
wire [flogtanh_WDTH -1:0]        I095672e79ca3a6dd8589b7821f06cdb9;
wire [MAX_SUM_WDTH_L-1:0]        I7383d68c9e1c7c663a32233a8385435a;
wire [MAX_SUM_WDTH_L-1:0]        Ie72268e979cf069b88f6eadde789e5ab;
wire [flogtanh_WDTH -1:0]        Ibf2f43980e835dd7ae7535957e3ec131;
wire [MAX_SUM_WDTH_L-1:0]        I8726f6e59d2146674ad4fae01d7f4135;
wire [MAX_SUM_WDTH_L-1:0]        I5732fdb805258fc13c8ba4aaf56574ca;
wire [flogtanh_WDTH -1:0]        Iaa980a50205025e3e1b09c6ce8ee53dd;
wire [MAX_SUM_WDTH_L-1:0]        I3a754b15a3a7d47b3a9741f4982a0a32;
wire [MAX_SUM_WDTH_L-1:0]        I3afe987d8f2c93cc19534a3221d1939c;
wire [flogtanh_WDTH -1:0]        I829aa657f0dd13c3fb86baeda8a3b4c8;
wire [MAX_SUM_WDTH_L-1:0]        I9bd8a06d5fdfe50c340c649a678ba2e2;
wire [MAX_SUM_WDTH_L-1:0]        Ic66af6c3c0268cfb0e9f0776c4f4e961;
wire [flogtanh_WDTH -1:0]        I1ae4334c32094064c19df0dac77bd03d;
wire [MAX_SUM_WDTH_L-1:0]        I215cb4bca0e3579af6474dbd9462304c;
wire [MAX_SUM_WDTH_L-1:0]        Ia605d14205926b3edc6d1c2f69f70ac0;
wire [flogtanh_WDTH -1:0]        I78788f7e0845e4353145012efa04a48c;
wire [MAX_SUM_WDTH_L-1:0]        I6d73cf92b5ad3ded496cf1363c87d3ad;
wire [MAX_SUM_WDTH_L-1:0]        I0071f2168787bd42ab7f2370aed9d0f5;
wire [flogtanh_WDTH -1:0]        I359f3e3bb2a69349f8564466fa81a054;
wire [MAX_SUM_WDTH_L-1:0]        I47851422267c2963b3c93e029e81fe1e;
wire [MAX_SUM_WDTH_L-1:0]        I4936f823841b0ffe32f801f5134c0211;
wire [flogtanh_WDTH -1:0]        I7b630e8ac26638fb858dd3b5d2d56385;
wire [MAX_SUM_WDTH_L-1:0]        Ie9cd13f4f83e446d41fa362d0ca005c2;
wire [MAX_SUM_WDTH_L-1:0]        I5975ef8f6cf53cf2132cdd9d707e7912;
wire [flogtanh_WDTH -1:0]        I859bef71501c2f2a994a0cdf8a94b2a7;
wire [MAX_SUM_WDTH_L-1:0]        I9990a45631a11aa0b051d237de4cb71f;
wire [MAX_SUM_WDTH_L-1:0]        I954ff0f9ee871a31774a3d786128fa13;
wire [flogtanh_WDTH -1:0]        Ib51b9e41161f4273f6469e8965acd7dd;
wire [MAX_SUM_WDTH_L-1:0]        I4be57c0a1c49baa53daba558c939eee0;
wire [MAX_SUM_WDTH_L-1:0]        I31f6bbfbbbd4c20d0c5c71663da1d4c1;
wire [flogtanh_WDTH -1:0]        I78bb23c008613c0f07f6f85172482296;
wire [MAX_SUM_WDTH_L-1:0]        I16d8c346fd377bc293763e9cb683566e;
wire [MAX_SUM_WDTH_L-1:0]        I1898bc3cc6a8b6f71d65c758d1f08366;
wire [flogtanh_WDTH -1:0]        I8b883a5bc22b2cde03f4074357be7c88;
wire [MAX_SUM_WDTH_L-1:0]        I9df0b548fc5a23180b48207dc7fc603e;
wire [MAX_SUM_WDTH_L-1:0]        If86532f849bd392dbf599eeb2fae0545;
wire [flogtanh_WDTH -1:0]        Ic2727e097ffbce70f07fc9f3d9395b54;
wire [MAX_SUM_WDTH_L-1:0]        I0b3b2dd5a443fab695d0ff59634b6cb6;
wire [MAX_SUM_WDTH_L-1:0]        Ia344734d285ac29b53cf401c08a0f987;
wire [flogtanh_WDTH -1:0]        I096397439036b0056c979054528ce1fd;
wire [MAX_SUM_WDTH_L-1:0]        I6f66b0df384980fcbf6a92e5a197575e;
wire [MAX_SUM_WDTH_L-1:0]        I502a8e382aa0881dc86f3c13e0566ca3;
wire [flogtanh_WDTH -1:0]        Ifcc83d9007aafdf32acf04f062e008c8;
wire [MAX_SUM_WDTH_L-1:0]        I2aff93633ddb7f63312e991dab99cfca;
wire [MAX_SUM_WDTH_L-1:0]        Ic462cebbfc39190b22d20013259e39eb;
wire [flogtanh_WDTH -1:0]        I53c01c60f4061d970e4491564ddf88ae;
wire [MAX_SUM_WDTH_L-1:0]        Ic17e0c2adccfc8b88818591fb7c3958a;
wire [MAX_SUM_WDTH_L-1:0]        I385d03def4cfb49f54867687ebd710ed;
wire [flogtanh_WDTH -1:0]        I0b4d34aa164c014f9315debd37fa534b;
wire [MAX_SUM_WDTH_L-1:0]        I835b69f77b77fcb0bb1cc9a05a9964c4;
wire [MAX_SUM_WDTH_L-1:0]        If8aa3ec1b5a4a3c122da82467be917da;
wire [flogtanh_WDTH -1:0]        Iac97aad4ca2c93e387ff0c1340143029;
wire [MAX_SUM_WDTH_L-1:0]        Iac61d3d6b4ebec5460d07a209317dbf6;
wire [MAX_SUM_WDTH_L-1:0]        I8daf79a0a2ee1bac7f055af441539fa4;
wire [flogtanh_WDTH -1:0]        I8b4c2d8a5f2b796029575ecf3b89e2b9;
wire [MAX_SUM_WDTH_L-1:0]        I762215c24e6cfbb27328534b48f6c013;
wire [MAX_SUM_WDTH_L-1:0]        I6261e0d339762cb2364421e6b87086cb;
wire [flogtanh_WDTH -1:0]        I06dd747316fa36a8dbdbb4ddf011230b;
wire [MAX_SUM_WDTH_L-1:0]        I278647e72fba32b7725004a889c40fb0;
wire [MAX_SUM_WDTH_L-1:0]        I0e2f746715b901feb69f6b3c94f3a828;
wire [flogtanh_WDTH -1:0]        I1594e7dfaedd9e7f5818dc4d639bb663;
wire [MAX_SUM_WDTH_L-1:0]        Ib6b14ee93e905e08b910d6011d780bf9;
wire [MAX_SUM_WDTH_L-1:0]        I7b8da162c08f8aa2ae90522ee1526cf6;
wire [flogtanh_WDTH -1:0]        Ic8111eb95e6b6ab35bcd8e2cafcd0c1e;
wire [MAX_SUM_WDTH_L-1:0]        I6f89d12b0e9b153b01cd8fd0e548a5ab;
wire [MAX_SUM_WDTH_L-1:0]        I5e8ecdbb018402b2fbc0049ee44bae8c;
wire [flogtanh_WDTH -1:0]        I650b4641d233096a77ae15c8254a29b1;
wire [MAX_SUM_WDTH_L-1:0]        I63ba8ed824c286ff8f68ffb6cb10a12c;
wire [MAX_SUM_WDTH_L-1:0]        I06d859184884c07a14c83d2f06587ad5;
wire [flogtanh_WDTH -1:0]        Ia905d37c471bdf7258a547be95b85e4f;
wire [MAX_SUM_WDTH_L-1:0]        Ib54c1747fb4316314527140212c7cc60;
wire [MAX_SUM_WDTH_L-1:0]        I79e3e49f57d47231c0fe6aaafdbc57f1;
wire [flogtanh_WDTH -1:0]        Icfc2b5de1aa36d81de3f163880d48a68;
wire [MAX_SUM_WDTH_L-1:0]        Idfaaf824ddb5452930ca1997f057e321;
wire [MAX_SUM_WDTH_L-1:0]        I12c07042202f66db926861c9ce7c2b25;
wire [flogtanh_WDTH -1:0]        I3c6893d360627cd954db1c20f3c9d319;
wire [MAX_SUM_WDTH_L-1:0]        I372410e0c71fce0d0a592bf9f16f822d;
wire [MAX_SUM_WDTH_L-1:0]        I9d0fdb45b9e86bd409740e538a690320;
wire [flogtanh_WDTH -1:0]        Ibc971e0b7ade69365d2c23f30ba0c1ea;
wire [MAX_SUM_WDTH_L-1:0]        Ie9392382734808bcff4da7e0c7f8e4d3;
wire [MAX_SUM_WDTH_L-1:0]        Id5fd6f25dc3df22a322434ae3c90dea6;
wire [flogtanh_WDTH -1:0]        I562d9a1676d27c7966d2920bb6be3b38;
wire [MAX_SUM_WDTH_L-1:0]        If703357df55e47b3ab1fbb1126ad5160;
wire [MAX_SUM_WDTH_L-1:0]        Id812a8ea2a3b4a912d151be582833fcf;
wire [flogtanh_WDTH -1:0]        I8aa258f382bea1eb300b006c3083bec1;
wire [MAX_SUM_WDTH_L-1:0]        I69e05d54d008abdfb8d0b2d1ddc0fd49;
wire [MAX_SUM_WDTH_L-1:0]        Ifd3638d44e1ba2285891fac152dee327;
wire [flogtanh_WDTH -1:0]        Iec0e7232ec94c15d7d50866ad5eb85fb;
wire [MAX_SUM_WDTH_L-1:0]        Ic79dc94346350619e49087d1d399bc39;
wire [MAX_SUM_WDTH_L-1:0]        Idd1b6014de2f053554ed09c29bf3e640;
wire [flogtanh_WDTH -1:0]        I0d252b23e06d25aee4afd84b4c5b4ba9;
wire [MAX_SUM_WDTH_L-1:0]        Ib805b36c4865846137bb8c620ee711bb;
wire [MAX_SUM_WDTH_L-1:0]        I0d96336eb4d5071d7e1d350e86513b25;
wire [flogtanh_WDTH -1:0]        I430703cef7ec173f9099c8391132e5c4;
wire [MAX_SUM_WDTH_L-1:0]        I8af4ba916324c47b2773e25e81eec395;
wire [MAX_SUM_WDTH_L-1:0]        I31e5b2cdc3dc571eafa37510076bcc64;
wire [flogtanh_WDTH -1:0]        I5788d966ba8393f5d76dcfcb9294b52e;
wire [MAX_SUM_WDTH_L-1:0]        I43bf51dd2065c4699e2efb0d23ca67fc;
wire [MAX_SUM_WDTH_L-1:0]        Ia8849f78971a45ed0daa2489e7d27dd7;
wire [flogtanh_WDTH -1:0]        Ied561890134d28b451f26da773ea5525;
wire [MAX_SUM_WDTH_L-1:0]        Ie42fb8850ec075e738c9265ef746d0a2;
wire [MAX_SUM_WDTH_L-1:0]        Ie4749f8e9ad2b370f9f9814b5a463c43;
wire [flogtanh_WDTH -1:0]        I52e018ad790a1e406777510a0f4b6c29;
wire [MAX_SUM_WDTH_L-1:0]        I734fecd29be258bbcf174ce05a4ad7c7;
wire [MAX_SUM_WDTH_L-1:0]        I3096d11098113da669ee0a94686e600d;
wire [flogtanh_WDTH -1:0]        I25eb66d8589cbb35b32cd25539a24f7f;
wire [MAX_SUM_WDTH_L-1:0]        I90c0a469b49cec5817be9ee089d7f035;
wire [MAX_SUM_WDTH_L-1:0]        I09a1d04c307fcb8a0e30925d86df3fe9;
wire [flogtanh_WDTH -1:0]        Icd4716d0d66d95a532544461c4872d11;
wire [MAX_SUM_WDTH_L-1:0]        I20467038010337e3e125bf2a7e1302d4;
wire [MAX_SUM_WDTH_L-1:0]        Idb0a98cea3ee6cd4308bfc2414a003e1;
wire [flogtanh_WDTH -1:0]        I266ba4229056534d310d982253b5f9b9;
wire [MAX_SUM_WDTH_L-1:0]        Idc01d14ecbd22e73d7ee052989eacff6;
wire [MAX_SUM_WDTH_L-1:0]        Id4788855f9a503e8b506d012aaeea445;
wire [flogtanh_WDTH -1:0]        I86498c8c820d276ac12764b5df267252;
wire [MAX_SUM_WDTH_L-1:0]        If3410ef0f48854e7b788d74904d03dad;
wire [MAX_SUM_WDTH_L-1:0]        I5b937934e7aae1f916c2848889f12685;
wire [flogtanh_WDTH -1:0]        I7bb9ad1a2cd32966746b05b7604a09b6;
wire [MAX_SUM_WDTH_L-1:0]        Icba9bcbb58a3fef701c5572510dbba65;
wire [MAX_SUM_WDTH_L-1:0]        I9275bb36e58e0f17964e13ee7f027ab7;
wire [flogtanh_WDTH -1:0]        Id0998cc2848a6a72ed2701a8e720946e;
wire [MAX_SUM_WDTH_L-1:0]        Ice5cb3b187d142f36c9fe4673952b229;
wire [MAX_SUM_WDTH_L-1:0]        I02330ade2eed926076cc071e45eed82c;
wire [flogtanh_WDTH -1:0]        If1ed051cd94d42e7836f82c10538b302;
wire [MAX_SUM_WDTH_L-1:0]        Id382353b13f6d198e0e9b90c5c3c16b3;
wire [MAX_SUM_WDTH_L-1:0]        I296bc392d4223cbdd6f77be6523df819;
wire [flogtanh_WDTH -1:0]        I780afd116929565d1ff9b3833ba242d5;
wire [MAX_SUM_WDTH_L-1:0]        I83efee0bf505cf1258bb68e419ffccf7;
wire [MAX_SUM_WDTH_L-1:0]        I31b0f2fe98cfddbc05dbd14be8be394b;
wire [flogtanh_WDTH -1:0]        I89ee99e699676bcec20031b6cad0e2ac;
wire [MAX_SUM_WDTH_L-1:0]        Id54f91bbae7215f942f539ca0834bd1f;
wire [MAX_SUM_WDTH_L-1:0]        Ia71663e8f563041c27cd21a0c9c27a28;
wire [flogtanh_WDTH -1:0]        I862b467403c045e4694fb57d59e10064;
wire [MAX_SUM_WDTH_L-1:0]        I810c80a4b57d13add447ee8964844ce1;
wire [MAX_SUM_WDTH_L-1:0]        Ib46b13498ec14ceaa56719f26f18febb;
wire [flogtanh_WDTH -1:0]        Ic3b554c66f652f027159dbc0fccc5ba3;
wire [MAX_SUM_WDTH_L-1:0]        Icf6d317a1bca3a6f3dfafdc9bdc0b805;
wire [MAX_SUM_WDTH_L-1:0]        I9bc2d5692474b8368c570d92835191b3;
wire [flogtanh_WDTH -1:0]        I04635713f6d70142b7ab3ecb5ffe6ac9;
wire [MAX_SUM_WDTH_L-1:0]        I47ca60b0a9bec684ec4e52f28f76c6d7;
wire [MAX_SUM_WDTH_L-1:0]        If8b0b96a659183e3651c691a2848b86b;
wire [flogtanh_WDTH -1:0]        I1917eae0dbcc0a941718c3248c7d4b11;
wire [MAX_SUM_WDTH_L-1:0]        I6ae68bcd4f3d39661626e4b671acf4ea;
wire [MAX_SUM_WDTH_L-1:0]        I87d958c00fc6209d901147831b0c951c;
wire [flogtanh_WDTH -1:0]        Ifa60c3079164485f31442d9cf12bd2ad;
wire [MAX_SUM_WDTH_L-1:0]        Iaa25b6dc9ec478e1fe096bfb9013752c;
wire [MAX_SUM_WDTH_L-1:0]        Ie4e4eaf3e5d2f581210af8054df71c6c;
wire [flogtanh_WDTH -1:0]        I5616405acf49c3e8608ae4d2b544b0d6;
wire [MAX_SUM_WDTH_L-1:0]        If7f010576686a2eb7aa5b2307c02ad6b;
wire [MAX_SUM_WDTH_L-1:0]        I0b557cf102da41afd26936cbdb64b6e8;
wire [flogtanh_WDTH -1:0]        Ie6f9ae463fa1add4de23463435a23d25;
wire [MAX_SUM_WDTH_L-1:0]        Ie8a683efbffce7c5676fa831573299d7;
wire [MAX_SUM_WDTH_L-1:0]        I49eb064043f91112c854e31e4eb9b885;
wire [flogtanh_WDTH -1:0]        Ib16a67d67a4650e53547312e3af60363;
wire [MAX_SUM_WDTH_L-1:0]        I50a4545b75d92b3c3209d473f8d0647c;
wire [MAX_SUM_WDTH_L-1:0]        I1039bc43e88eee527d2ed6adb8c7d1ba;
wire [flogtanh_WDTH -1:0]        I8fa4ad645ca2ef21dea8669d2e2afbe2;
wire [MAX_SUM_WDTH_L-1:0]        Ib0e11d415f14d70a626c6f0dfeed2e37;
wire [MAX_SUM_WDTH_L-1:0]        I9aab16e89f1b64117caece8ca8af5940;
wire [flogtanh_WDTH -1:0]        I41ea2e3d798ff8e0a95f04e4773c59b4;
wire [MAX_SUM_WDTH_L-1:0]        I3a6167a349b5dce1dfa66859bfd5eee7;
wire [MAX_SUM_WDTH_L-1:0]        I343df614f97cf732e57cf2ad3f95dc9e;
wire [flogtanh_WDTH -1:0]        Id7f4c6208197cdbf48fecdb2a18b81fc;
wire [MAX_SUM_WDTH_L-1:0]        I566fd98c8c6ebf6e2d8ebace4b8b358b;
wire [MAX_SUM_WDTH_L-1:0]        Ie02de90d8eb06b16314946d21299500c;
wire [flogtanh_WDTH -1:0]        I0adb66417482782dd71da1678c1f7412;
wire [MAX_SUM_WDTH_L-1:0]        Ib777f0ff44b2847294370d74f741b70b;
wire [MAX_SUM_WDTH_L-1:0]        I3353a7916b569f2c0ca122180608dccc;
wire [flogtanh_WDTH -1:0]        I2abe89a1366a1ad862266ad88101baa2;
wire [MAX_SUM_WDTH_L-1:0]        I6cd7374654c74b4be21b6a3639ddac0f;
wire [MAX_SUM_WDTH_L-1:0]        Ibfe760474fcac99f1e5ffa2e008fef99;
wire [flogtanh_WDTH -1:0]        I8d10f0c6dc026005f7882ca013283099;
wire [MAX_SUM_WDTH_L-1:0]        I930319dcb4988822341ac101fef3dc52;
wire [MAX_SUM_WDTH_L-1:0]        I3caf1211dcbcdc746a3e4c7fbbdae4a8;
wire [flogtanh_WDTH -1:0]        I4ef16908ce9b89771f94068eec1a983e;
wire [MAX_SUM_WDTH_L-1:0]        If556f828f8cb4c1f1721e9d12977ec5a;
wire [MAX_SUM_WDTH_L-1:0]        I2dcc0d17b9fcac35693bf32b5c5540fd;
wire [flogtanh_WDTH -1:0]        I4f6bcd6e0bcd77730248b69d2b93c904;
wire [MAX_SUM_WDTH_L-1:0]        If7df1cceb63540263742300063a2febb;
wire [MAX_SUM_WDTH_L-1:0]        Ie6764a631310e312ba5c2c1e601d828f;
wire [flogtanh_WDTH -1:0]        Iea1ae39e18f083fb8f855fd9ad3d4f8e;
wire [MAX_SUM_WDTH_L-1:0]        Idb605ffe97f2a0cbc2b260464afd1479;
wire [MAX_SUM_WDTH_L-1:0]        I220f8e45e5fe6e69f02cded87f12e1e5;
wire [flogtanh_WDTH -1:0]        I795ae30dec63ef2952917eb3355148a2;
wire [MAX_SUM_WDTH_L-1:0]        I8690851e49869591791e5202e2ef2432;
wire [MAX_SUM_WDTH_L-1:0]        I896cd566a3d078b0f697a788efd223f2;
wire [flogtanh_WDTH -1:0]        I188813c5474bf304b59dbe07c78bef6f;
wire [MAX_SUM_WDTH_L-1:0]        I60d3d03ea9219db9501568fb71d87df0;
wire [MAX_SUM_WDTH_L-1:0]        I7caa41076a293edf18c7c4309fdcfc91;
wire [flogtanh_WDTH -1:0]        I1760a42d85513ea751e94a8b829b5f1a;
wire [MAX_SUM_WDTH_L-1:0]        Ib7f80c4193c311c6c553f15f0d9e0e09;
wire [MAX_SUM_WDTH_L-1:0]        I928a0e4951208aab170656596f456209;
wire [flogtanh_WDTH -1:0]        I8c652055cfcd230426887e171eaf2511;
wire [MAX_SUM_WDTH_L-1:0]        I3dfabb54fefcb9b9896e52446a1edc25;
wire [MAX_SUM_WDTH_L-1:0]        Ia3d129fd297905bee180293c0c39d9ef;
wire [flogtanh_WDTH -1:0]        I9a88a91b0fcc6dd1a7b4ed24e676d9e1;
wire [MAX_SUM_WDTH_L-1:0]        If35ab032940f067a7905284b5f34a795;
wire [MAX_SUM_WDTH_L-1:0]        Id555c88cf7f0904db74d45cc75c8f5d6;
wire [flogtanh_WDTH -1:0]        I89f6566e2295d58668e63b9529d94df8;
wire [MAX_SUM_WDTH_L-1:0]        I11cbc38d0e7e8bb159707d0b6a312049;
wire [MAX_SUM_WDTH_L-1:0]        I1ddfd31bbf062aa5c3c71d61e492e3a2;
wire [flogtanh_WDTH -1:0]        I08295c218fd06a8900974edc9c2924f2;
wire [MAX_SUM_WDTH_L-1:0]        Ib39a30cd08168accc0c3ca3bda467878;
wire [MAX_SUM_WDTH_L-1:0]        Iae9e023628eb6686708b2656f15616cc;
wire [flogtanh_WDTH -1:0]        I0a39fdea8b5bfac1862f199152e26ffe;
wire [MAX_SUM_WDTH_L-1:0]        I44afd98669c6e6bf5054d677de2b919c;
wire [MAX_SUM_WDTH_L-1:0]        If4b100d26126e460c41b8c1bc8fbbb96;
wire [flogtanh_WDTH -1:0]        Ib36a71ff310882325be0a2745e48f708;
wire [MAX_SUM_WDTH_L-1:0]        Ic75ef170613d6b56ad3928b88f1abef5;
wire [MAX_SUM_WDTH_L-1:0]        I85a7fede715578be0634d71e9c7951cd;
wire [flogtanh_WDTH -1:0]        I75e4d037cc2ed0b0f75fc1fe9cb21da3;
wire [MAX_SUM_WDTH_L-1:0]        If541dad0db59ce6598cc87b2ecf6d76a;
wire [MAX_SUM_WDTH_L-1:0]        I2d7715a3af03d9664729fa6df85034a2;
wire [flogtanh_WDTH -1:0]        Iee9e9849924642a9579a10655624fa17;
wire [MAX_SUM_WDTH_L-1:0]        I3e9f3d8ae099408fe2ff46ae3aff430e;
wire [MAX_SUM_WDTH_L-1:0]        I571ddcb0a10938e4c0816c965214b4a8;
wire [flogtanh_WDTH -1:0]        I0a267feb8313c9fa5c663a3fe68284dd;
wire [MAX_SUM_WDTH_L-1:0]        I6688f7cccc769490e870707ba9c14991;
wire [MAX_SUM_WDTH_L-1:0]        I8bf8b0cf27a2654a0e7fdf3255945b67;
wire [flogtanh_WDTH -1:0]        I0e0ff3511e65a1dda10ec944c89d09d7;
wire [MAX_SUM_WDTH_L-1:0]        I89d5eb773f6c952c1ed5e5c57fed6fe1;
wire [MAX_SUM_WDTH_L-1:0]        I63f82f075d53205b5b556c0054f1a0b8;
wire [flogtanh_WDTH -1:0]        I4504a0a17633d26163a0afae21ad0f43;
wire [MAX_SUM_WDTH_L-1:0]        Ia55fb2a1a8fcd959e3dd99403cd39a97;
wire [MAX_SUM_WDTH_L-1:0]        I3c6fb0df5846a19228a4e6cf9f9106ac;
wire [flogtanh_WDTH -1:0]        Ibd7b7f4ba86b6c61a0dd38f71c67ae05;
wire [MAX_SUM_WDTH_L-1:0]        I51a2b9abfab582408aeea3130d1e8334;
wire [MAX_SUM_WDTH_L-1:0]        I7168b0efdd2fae57292379c9d15c62eb;
wire [flogtanh_WDTH -1:0]        Icddd184270ffda26b803956883400ad0;
wire [MAX_SUM_WDTH_L-1:0]        Id1bc8bf048edb72a3564f864e8fb8671;
wire [MAX_SUM_WDTH_L-1:0]        Ibe502ebbb366f54a8f8fda4e361308e3;
wire [flogtanh_WDTH -1:0]        Id3da7061c05091ffc520d4480058e8e9;
wire [MAX_SUM_WDTH_L-1:0]        I7aa45db0b1c7bd90b21c438b91070a16;
wire [MAX_SUM_WDTH_L-1:0]        Ifce70fefde8f5ea4d2c1857236f66d65;
wire [flogtanh_WDTH -1:0]        Ie63d649228270b34d8ed25e7c4b09883;
wire [MAX_SUM_WDTH_L-1:0]        I4673a5950ad69c59f3cf4001a1dc93d2;
wire [MAX_SUM_WDTH_L-1:0]        Ice2c390d296e09b117d60905343e9098;
wire [flogtanh_WDTH -1:0]        I8eed3f7b36c046fff1e41dd52a300d29;
wire [MAX_SUM_WDTH_L-1:0]        Iffb8eaecd6bd058181a4532d83f674a5;
wire [MAX_SUM_WDTH_L-1:0]        I4b94402a53d981e953c21ef316c709b7;
wire [flogtanh_WDTH -1:0]        Iefcebe38e0c2d6d570017e165d70d3b1;
wire [MAX_SUM_WDTH_L-1:0]        I0a7e192f836bc8f7c0ea6bd7a66adaa7;
wire [MAX_SUM_WDTH_L-1:0]        I450c0d6ad5d3b1f18bb28e3a432b5442;
wire [flogtanh_WDTH -1:0]        Ia153222350357443978d7426663c3eaa;
wire [MAX_SUM_WDTH_L-1:0]        Ic38ac13f1b1f78c5e83379cabf407f5a;
wire [MAX_SUM_WDTH_L-1:0]        I2587a5800a5a9ffeabc4dca503e3d964;
wire [flogtanh_WDTH -1:0]        I06f0fd2d9d46a2fdb4221217ee2496d1;
wire [MAX_SUM_WDTH_L-1:0]        Ie9b7108feaaa1fd3e2dc5eeba3d6c4e5;
wire [MAX_SUM_WDTH_L-1:0]        I1182655739d7ab5bbe4a6546a5ca36fd;
wire [flogtanh_WDTH -1:0]        I9533ff0882ed01409795d7269329fd76;
wire [MAX_SUM_WDTH_L-1:0]        Iab83df9535036f6c0108658ebd03620a;
wire [MAX_SUM_WDTH_L-1:0]        I8110a5a62607093b21b7cd088b1d9ee0;
wire [flogtanh_WDTH -1:0]        Ia9eb9821e7dc31c23d7e60839949c1ff;
wire [MAX_SUM_WDTH_L-1:0]        I5dac976084afd52f5b0d21306bcbb511;
wire [MAX_SUM_WDTH_L-1:0]        I8b611f7c12ddd81de403ba74e212857f;
wire [flogtanh_WDTH -1:0]        I3663fc86620d6244a850819bd3ebe72c;
wire [MAX_SUM_WDTH_L-1:0]        I018c59ff182308d3ca739dbe309ba91e;
wire [MAX_SUM_WDTH_L-1:0]        I84a62a133dbceb5a32a7c907f371663d;
wire [flogtanh_WDTH -1:0]        I11293e7cdeddf352011d46abd6c3bb72;
wire [MAX_SUM_WDTH_L-1:0]        I9a117a38c8db8191f34cfe7a403aa135;
wire [MAX_SUM_WDTH_L-1:0]        Ia2fc8a1bbc3cb0dd7d89a7f05b04909c;
wire [flogtanh_WDTH -1:0]        Ic9339e415d0f756e34bcd930de63ad87;
wire [MAX_SUM_WDTH_L-1:0]        I60d5a8f56d1f22d535a53bbba3049a56;
wire [MAX_SUM_WDTH_L-1:0]        I2a3eb42a4402e873d081f94a14a99c20;
wire [flogtanh_WDTH -1:0]        Icf109f65e24d3a23ecad9e7d4cc54dc1;
wire [MAX_SUM_WDTH_L-1:0]        I270d4c8baa595241fcc0060b18749f4f;
wire [MAX_SUM_WDTH_L-1:0]        I58447d6ae49a6be2d043477a06f83df0;
wire [flogtanh_WDTH -1:0]        Idf7dd0ff83b2d56693e729a1a375fabb;
wire [MAX_SUM_WDTH_L-1:0]        I765d0dd290e34cee0116f45ce9527117;
wire [MAX_SUM_WDTH_L-1:0]        I83292bcda4645233d8e8a1dfe8e5f60b;
wire [flogtanh_WDTH -1:0]        I312a248019372261c0959cdc9378ec93;
wire [MAX_SUM_WDTH_L-1:0]        I9ef68d76daf35fa29a0c4168baf64516;
wire [MAX_SUM_WDTH_L-1:0]        Ic5e0a84cf1a2ef907b2456559ea26c75;
wire [flogtanh_WDTH -1:0]        I8e311b9891dda272762da2c640019e8c;
wire [MAX_SUM_WDTH_L-1:0]        Icc9faf407342c704a8f33b49c1ad8063;
wire [MAX_SUM_WDTH_L-1:0]        I2cefbf897bb7f6f67ca500727e85c683;
wire [flogtanh_WDTH -1:0]        I1874dd9f7c0a93310873173561402912;
wire [MAX_SUM_WDTH_L-1:0]        Ibdfcf91a62d88e9b8d011a22c8100106;
wire [MAX_SUM_WDTH_L-1:0]        If47be2ca4617a426258c51f8d977ba3f;
wire [flogtanh_WDTH -1:0]        I04adb3964e739a106098a6c4d2f49e94;
wire [MAX_SUM_WDTH_L-1:0]        I6ff243d4d70ead40034f55f7b0c49557;
wire [MAX_SUM_WDTH_L-1:0]        I7c68e0ae30efc4ca4d68b6047119c6c3;
wire [flogtanh_WDTH -1:0]        I9135b709c3c802a42c7186087b5664cc;
wire [MAX_SUM_WDTH_L-1:0]        I6fe27a172bfa6cd64ae70b8a22f66e4a;
wire [MAX_SUM_WDTH_L-1:0]        Iccca1936f4c1c9496205e77b588e9985;
wire [flogtanh_WDTH -1:0]        Ia236dfe34ff4938456d76f787d2db945;
wire [MAX_SUM_WDTH_L-1:0]        I20b96db33a7f876f9b37e0dd13d39630;
wire [MAX_SUM_WDTH_L-1:0]        I59d4567d3355fdae5660a1364d1b8d00;
wire [flogtanh_WDTH -1:0]        I41c98bae5fbdb31bac0913930573e80c;
wire [MAX_SUM_WDTH_L-1:0]        Ic1c711155cf28a3491f52352d5fbd05a;
wire [MAX_SUM_WDTH_L-1:0]        I4600963866dcb9bbea2515c805f885cb;
wire [flogtanh_WDTH -1:0]        I226befd72285893998aca87fe34d9aaf;
wire [MAX_SUM_WDTH_L-1:0]        Ic99fca70349dfdfdbec515ab163ad20f;
wire [MAX_SUM_WDTH_L-1:0]        If26d90629e70c5a871e6f5b14471b8cf;
wire [flogtanh_WDTH -1:0]        I20ab7c6174af39aee99492f704b2748c;
wire [MAX_SUM_WDTH_L-1:0]        I71db278548cbf6a478f5f2d7de410dc9;
wire [MAX_SUM_WDTH_L-1:0]        Iedb9bb14951bf67bc8865b0983490c14;
wire [flogtanh_WDTH -1:0]        I0a1c5724ffa14df653142a1f8bcf44a4;
wire [MAX_SUM_WDTH_L-1:0]        I67f75dfd3165ca969119ededc4c25b1d;
wire [MAX_SUM_WDTH_L-1:0]        I6a3854ed571e8c262aa3ec377c247778;
wire [flogtanh_WDTH -1:0]        I481973954b81accf069dd80830fba3bc;
wire [MAX_SUM_WDTH_L-1:0]        Ia4f05220e30b257689f831feaa0125e9;
wire [MAX_SUM_WDTH_L-1:0]        I05028975b49ec0c089bd981696f85a8b;
wire [flogtanh_WDTH -1:0]        Ia6825c3edc9d2a6832db7a7d684faf98;
wire [MAX_SUM_WDTH_L-1:0]        Ieeaf2a662a0f9295b3c3d6454f731098;
wire [MAX_SUM_WDTH_L-1:0]        Ife732309efcc740cfff5c747aab2e3d6;
wire [flogtanh_WDTH -1:0]        I5c964036207f47629302e282d56fef7b;
wire [MAX_SUM_WDTH_L-1:0]        Id7e4f0f2bded6e1d39467d074348b324;
wire [MAX_SUM_WDTH_L-1:0]        Idcef10a0465614cf38e0d6f503b5174a;
wire [flogtanh_WDTH -1:0]        I00b74ed4d6730b37c6fbfd42dee42584;
wire [MAX_SUM_WDTH_L-1:0]        I4c556e88e578d8f5d2d529b33a00b9eb;
wire [MAX_SUM_WDTH_L-1:0]        Ibd4aaf02982068ffbfd1b8b3795d9217;
wire [flogtanh_WDTH -1:0]        I0345fc4a507f9e3be3e1d46b71693de1;
wire [MAX_SUM_WDTH_L-1:0]        I25facb36e0360a4ca4ac5803101984c7;
wire [MAX_SUM_WDTH_L-1:0]        I788c64785b992c675fe348a1fa181525;
wire [flogtanh_WDTH -1:0]        I9f0735c1cf5d1af7c82a251ef4886f9c;
wire [MAX_SUM_WDTH_L-1:0]        Iab18a2d81fc63ba2b35df1cdf08621af;
wire [MAX_SUM_WDTH_L-1:0]        Ib235af5b28d56f24372d3f0af816f2c2;
wire [flogtanh_WDTH -1:0]        I861cf5dffb18c84953013dc4026bd08a;
wire [MAX_SUM_WDTH_L-1:0]        Icd609cdfdfa1ecb62bba040a015b8de5;
wire [MAX_SUM_WDTH_L-1:0]        I4c03a6569d1b954d088053e38827e811;
wire [flogtanh_WDTH -1:0]        I19722ceada71cc9cc06edde39142ff17;
wire [MAX_SUM_WDTH_L-1:0]        I00c895c62ee2842ad86d01beab41e900;
wire [MAX_SUM_WDTH_L-1:0]        Idda26504e422367082caeafbb29871f9;
wire [flogtanh_WDTH -1:0]        Id8349128e2c391df008828494da928c6;
wire [MAX_SUM_WDTH_L-1:0]        Idd279726169e173c111b7c490a2c4037;
wire [MAX_SUM_WDTH_L-1:0]        I195c3a82123142d509886ee37dc6fc98;
wire [flogtanh_WDTH -1:0]        I27209805df490a07f1726875a7b69922;
wire [MAX_SUM_WDTH_L-1:0]        I125a005c7f9d37d5365496513fef1893;
wire [MAX_SUM_WDTH_L-1:0]        I1abb512ca0383c9e7104418e07281841;
wire [flogtanh_WDTH -1:0]        I7532c1f0624a2d5a94321c89c73e38df;
wire [MAX_SUM_WDTH_L-1:0]        I62802ceb2a05dc315e7137f31590cc72;
wire [MAX_SUM_WDTH_L-1:0]        I00ff1331b1900bb031ee81d2a58c1bd5;
wire [flogtanh_WDTH -1:0]        Ife892846e66e2522c06b170811a11ada;
wire [MAX_SUM_WDTH_L-1:0]        I5b0fda1e3b1829738e08b1de1d934a1c;
wire [MAX_SUM_WDTH_L-1:0]        If65eb5e743a7b1878fb232ef2fe13cb0;
wire [flogtanh_WDTH -1:0]        Ib905ede2830f7e3c8cf993075f07345c;
wire [MAX_SUM_WDTH_L-1:0]        I0f86873fc1d12c964a3757bec70ad780;
wire [MAX_SUM_WDTH_L-1:0]        I24ae7de3549a84f4f88f561b6017b7a8;
wire [flogtanh_WDTH -1:0]        Ibf169f844d9e00eca8f3821ddc952ef0;
wire [MAX_SUM_WDTH_L-1:0]        I6f41f58cfeab93cd06c32cd2537426dd;
wire [MAX_SUM_WDTH_L-1:0]        I449c77140475475b138d839a74078337;
wire [flogtanh_WDTH -1:0]        I3137f75629e72f78abdac088e18608d5;
wire [MAX_SUM_WDTH_L-1:0]        Ibf529f3a5b5f9d44d2e072b2cfb0c987;
wire [MAX_SUM_WDTH_L-1:0]        Ia9e102d8679943c079f16c0228f0f0d1;
wire [flogtanh_WDTH -1:0]        I8fbcabc2f5c30fcf1c5b46de5dfe887d;
wire [MAX_SUM_WDTH_L-1:0]        I189af406b34e849a5700be4ea8d7a22b;
wire [MAX_SUM_WDTH_L-1:0]        Ibf1c9d86665f696d91c554db748ff42b;
wire [flogtanh_WDTH -1:0]        Ie7acfb624aa6242b558481350c85fda3;
wire [MAX_SUM_WDTH_L-1:0]        I2e6d80f71d9e42ef5e32d8e43c9ad77e;
wire [MAX_SUM_WDTH_L-1:0]        Ieb0336a1974a2aec0966f4f59f460802;
wire [flogtanh_WDTH -1:0]        I11e0b915338d5d649c800455b9a7695f;
wire [MAX_SUM_WDTH_L-1:0]        I8a8379ec2c6c9c360b2c32c34e63902d;
wire [MAX_SUM_WDTH_L-1:0]        Ic0819ccefe784a6379716b3633ae0196;
wire [flogtanh_WDTH -1:0]        Ia9e4e68dcd3d0281decde939eed0c3bd;
wire [MAX_SUM_WDTH_L-1:0]        Ic89ee3a7462610019feee4023e1ab63e;
wire [MAX_SUM_WDTH_L-1:0]        I0c4bbd1827b1859caabb067e864ce4b3;
wire [flogtanh_WDTH -1:0]        Id508f63a381fc565a28fe4e662b33efb;
wire [MAX_SUM_WDTH_L-1:0]        I49b0d9feed7042dc0551398d48b36f7f;
wire [MAX_SUM_WDTH_L-1:0]        I004c98da87996b77b5761d366210f782;
wire [flogtanh_WDTH -1:0]        I33582dc83370e68b0ae7b22b553276b4;
wire [MAX_SUM_WDTH_L-1:0]        Icfbd9d5dfe741fd84977d13887a54dee;
wire [MAX_SUM_WDTH_L-1:0]        Ia457938da4efe847cb06f645f2a54a52;
wire [flogtanh_WDTH -1:0]        I8aeca996ad6820edcc6fcbaa8a0f15ce;
wire [MAX_SUM_WDTH_L-1:0]        Ib2b669872ca023cf13754a529eab5ad5;
wire [MAX_SUM_WDTH_L-1:0]        I7e0474089ebc1c34747be1bc17a81d72;
wire [flogtanh_WDTH -1:0]        Ica86e8037319b868c8cb89f3cb02b136;
wire [MAX_SUM_WDTH_L-1:0]        Ife9a683c5c06abb98e9a9da56244cadf;
wire [MAX_SUM_WDTH_L-1:0]        Ib0b46b99e61d724ae664d9d1fec1e29f;
wire [flogtanh_WDTH -1:0]        Ia95013b19d9fc12d19ff9924007113d4;
wire [MAX_SUM_WDTH_L-1:0]        Ic2a2da3827248989cad50ff9fcc8822e;
wire [MAX_SUM_WDTH_L-1:0]        I56d1025271f1f7704a40dd7f0df02b0b;
wire [flogtanh_WDTH -1:0]        Ifcf979b713b014f22c1c8ce1d42132c2;
wire [MAX_SUM_WDTH_L-1:0]        Ifcbb960ba610a378b0472f005bea218a;
wire [MAX_SUM_WDTH_L-1:0]        I72c2256ba47cf03f95143df8f741fd83;
wire [flogtanh_WDTH -1:0]        I973b3306021532f286cf248084398c26;
wire [MAX_SUM_WDTH_L-1:0]        I9527b33b0941a515601b7fb75c0eba34;
wire [MAX_SUM_WDTH_L-1:0]        I733c3fa4d84e5680792b16a70bb1a51d;
wire [flogtanh_WDTH -1:0]        Iea7940bb396d1a436f56806fc533edee;
wire [MAX_SUM_WDTH_L-1:0]        Ia65e331b9f0ec80ee7860b2c4a6c1e55;
wire [MAX_SUM_WDTH_L-1:0]        If367d63311c96726517240de13bd2a4b;
wire [flogtanh_WDTH -1:0]        Ied55045b003302c294591a8d2a6a39fd;
wire [MAX_SUM_WDTH_L-1:0]        I2cbdbbf07d938e2f4847fdf594a010c8;
wire [MAX_SUM_WDTH_L-1:0]        Icc6d895d943e14f2801c22e79ce190e8;
wire [flogtanh_WDTH -1:0]        Ib64e948413d5dce1d9309fe95c0919ab;
wire [MAX_SUM_WDTH_L-1:0]        I260ec6308196983b8aeaddcac953709d;
wire [MAX_SUM_WDTH_L-1:0]        Ieb664ac9be65fba2e25960141f7fb4b6;
wire [flogtanh_WDTH -1:0]        I682fe6c6c621db5dd867574e8573d8ed;
wire [MAX_SUM_WDTH_L-1:0]        I456482f0ce8cb6c76d2b19b69cd0f4fc;
wire [MAX_SUM_WDTH_L-1:0]        I66071f20991b414140869a2e3b750471;
wire [flogtanh_WDTH -1:0]        I508b57f6ebc45eb70aa7b114096a7d12;
wire [MAX_SUM_WDTH_L-1:0]        Ie9d6a3cf41e366e12a6d90a61163fb48;
wire [MAX_SUM_WDTH_L-1:0]        Iffeefa89a2ba7d032db5db64cbf05e20;
wire [flogtanh_WDTH -1:0]        I8e82b8914260669ed1d88a690467a7b4;
wire [MAX_SUM_WDTH_L-1:0]        Ieb526cf88e7ac70a26f05c0f56d37c91;
wire [MAX_SUM_WDTH_L-1:0]        I9ab3cea6ee8d8473221da21bae06066b;
wire [flogtanh_WDTH -1:0]        I525feb94b558fb4bb8db8eead9f05afa;
wire [MAX_SUM_WDTH_L-1:0]        If4ccf2222e01f9418f342054b342412f;
wire [MAX_SUM_WDTH_L-1:0]        I3403ce6e697b523a9f441d8fd5e2d420;
wire [flogtanh_WDTH -1:0]        Ie5e4cf2b42054822a9091f5ef67cd968;
wire [MAX_SUM_WDTH_L-1:0]        I0875d93243187e274b27f729a86dd9fa;
wire [MAX_SUM_WDTH_L-1:0]        Ia98a70144e466b356d2998948dc4b602;
wire [flogtanh_WDTH -1:0]        I0d08d26e31c8b69ed8c089cdcd055a50;
wire [MAX_SUM_WDTH_L-1:0]        Ibd4f6d59420fe37742ef3ae1f22c152c;
wire [MAX_SUM_WDTH_L-1:0]        Ie4ca0836695d951ee09622892ee35928;
wire [flogtanh_WDTH -1:0]        I877f44c880a781381bfa8a8f8471d697;
wire [MAX_SUM_WDTH_L-1:0]        I2f726cba2feffeaeeadff790c6909402;
wire [MAX_SUM_WDTH_L-1:0]        I485a48b4ff4da08f977425fd10e6d392;
wire [flogtanh_WDTH -1:0]        I7fc78273dc765cf1c03b3c1a043b35f8;
wire [MAX_SUM_WDTH_L-1:0]        Id8d5b7c74ba1b051e3e4eb87d812e028;
wire [MAX_SUM_WDTH_L-1:0]        Ie8c79e6a5378808c0ead5a4b24319ce9;
wire [flogtanh_WDTH -1:0]        Ie67275a4b3fdc050f0f6e7ac7d1eebfc;
wire [MAX_SUM_WDTH_L-1:0]        I2c853ac0b4a3ac567a4db08ba5e9e26d;
wire [MAX_SUM_WDTH_L-1:0]        I9ca81c841a75a9ac242835956509e0fe;
wire [flogtanh_WDTH -1:0]        I41f9acc96650353174155a5f378d5cc5;
wire [MAX_SUM_WDTH_L-1:0]        Ifa2b0aa146869b9f6238969c5649acc7;
wire [MAX_SUM_WDTH_L-1:0]        Id50f18f642f3b00ffa34986f78a0eae6;
wire [flogtanh_WDTH -1:0]        I0d73c905b2ed777acd71d560928dcf0b;
wire [MAX_SUM_WDTH_L-1:0]        Ib4322244b363748db4a0543933452669;
wire [MAX_SUM_WDTH_L-1:0]        I75838ca09e301b8e1301cbf603a1f8c2;
wire [flogtanh_WDTH -1:0]        I2b6b1c25caf8b00d19ccc98156a8ca2b;
wire [MAX_SUM_WDTH_L-1:0]        Idbd452a90ce7a7c82d5d2d7f57fbd72c;
wire [MAX_SUM_WDTH_L-1:0]        Id968b34075e351ab01d65abcb4ed8cca;
wire [flogtanh_WDTH -1:0]        I28ea2b207bcd3518a85ff150466a6a08;
wire [MAX_SUM_WDTH_L-1:0]        I28ceab58b644f619bb359f153087cb9b;
wire [MAX_SUM_WDTH_L-1:0]        I84da4ce7441e132e775167c1cd81dbe5;
wire [flogtanh_WDTH -1:0]        I7d0a1c64b2e85e1bf0bf99423321466b;
wire [MAX_SUM_WDTH_L-1:0]        Iaf75fbdcad76103a769669bc20d0c5b7;
wire [MAX_SUM_WDTH_L-1:0]        If19dc22d45cc4664c85a043ec4c00617;
wire [flogtanh_WDTH -1:0]        I3b9b9b41b54ff194314b572a15daf606;
wire [MAX_SUM_WDTH_L-1:0]        I4a34573ee0f529e4088f1b5969eee325;
wire [MAX_SUM_WDTH_L-1:0]        Ibf482db0f5058be72061267c42ebc292;
wire [flogtanh_WDTH -1:0]        Ic914f847e623d9c52e2d9ae5076c21c3;
wire [MAX_SUM_WDTH_L-1:0]        I0602ea657e22176e268c3f005b327c5f;
wire [MAX_SUM_WDTH_L-1:0]        I6d2dbb953a58b91dafa7f0d34d41bdc3;
wire [flogtanh_WDTH -1:0]        I46fc20938dd554b23b5af5f7c3e39480;
wire [MAX_SUM_WDTH_L-1:0]        I48ef1d4bacb30b7602392e7298e88c40;
wire [MAX_SUM_WDTH_L-1:0]        Ib393146d81d3cf031466543311cee2ad;
wire [flogtanh_WDTH -1:0]        I1fa8b37b4697ae60cf399285d9524b8d;
wire [MAX_SUM_WDTH_L-1:0]        I36272af5470aa53e7c61cbc896f26290;
wire [MAX_SUM_WDTH_L-1:0]        I42564ec6a794ea803795f0b5b3523a93;
wire [flogtanh_WDTH -1:0]        I66c8261df769288836e188ecb32b6dc6;
wire [MAX_SUM_WDTH_L-1:0]        I146bdc684c432e98b5e1c3b274f3272c;
wire [MAX_SUM_WDTH_L-1:0]        I4a0033a180d7edce81fcfef603532e28;
wire [flogtanh_WDTH -1:0]        I267714c8a5aa14bae9c74da272a60aa5;
wire [MAX_SUM_WDTH_L-1:0]        I723e72d69796cee0c174c82c2514cd7c;
wire [MAX_SUM_WDTH_L-1:0]        Ic7a21921e2716fba55aad2e351f4498a;
wire [flogtanh_WDTH -1:0]        I47a34c8d2174c12f96041e82ad835db2;
wire [MAX_SUM_WDTH_L-1:0]        I305b258a587eb0f55a48679ab7ddcf91;
wire [MAX_SUM_WDTH_L-1:0]        I9a3f0b4867087790c78f674b719dbf7b;
wire [flogtanh_WDTH -1:0]        If99ca487495a015063fd8dc54ae596aa;
wire [MAX_SUM_WDTH_L-1:0]        Ia8a328c524c386c6008d76d6c920ab03;
wire [MAX_SUM_WDTH_L-1:0]        I138f008a6206a1067bb0e22ce3d90990;
wire [flogtanh_WDTH -1:0]        I1043f1b92b49a8c304a23c0b5c615def;
wire [MAX_SUM_WDTH_L-1:0]        I5269f5ff21c0c874811b85f6a028c113;
wire [MAX_SUM_WDTH_L-1:0]        I48ad9b737892d7c49340ed679f46e034;
wire [flogtanh_WDTH -1:0]        Icafa102383ef33455236ba268b1b7460;
wire [MAX_SUM_WDTH_L-1:0]        I93671d398af3e4f197eb71233121de97;
wire [MAX_SUM_WDTH_L-1:0]        I04a9c9765fd468a7e841577f09fc287b;
wire [flogtanh_WDTH -1:0]        I677fca8017154fed3e6cd54362e829db;
wire [MAX_SUM_WDTH_L-1:0]        Ia26b08bdae3e484e917194c100e1763d;
wire [MAX_SUM_WDTH_L-1:0]        I7b929c228c865112f00bc6b4dcc95b52;
wire [flogtanh_WDTH -1:0]        I826fe051a6b09d5cacf712431ce89b7c;
wire [MAX_SUM_WDTH_L-1:0]        I9fa2896c4dbd25ed089fce8d5ce372b2;
wire [MAX_SUM_WDTH_L-1:0]        I2b54a135e59945901e9c11580a29ee3d;
wire [flogtanh_WDTH -1:0]        I23f781ebfa449cec7975b94179d72259;
wire [MAX_SUM_WDTH_L-1:0]        I1e4586148b049d4493e1cafe947c3983;
wire [MAX_SUM_WDTH_L-1:0]        I566221060f06e724676ec9bec861d7de;
wire [flogtanh_WDTH -1:0]        Ia383b5dc3b7ce1bc7987926535639668;
wire [MAX_SUM_WDTH_L-1:0]        I375aeddea735459513ef97aec26fc8d1;
wire [MAX_SUM_WDTH_L-1:0]        Icd9a876a0feb16ea62bcad5be2004dac;
wire [flogtanh_WDTH -1:0]        I40ae857caffae41564c2ecb0c7e9777b;
wire [MAX_SUM_WDTH_L-1:0]        I683f128be784d4e752ea5881c1d483a8;
wire [MAX_SUM_WDTH_L-1:0]        I8f8273c4cb2a9ace8a09847efd4bdec7;
wire [flogtanh_WDTH -1:0]        I569d56a2673a104f3050d851d767af8a;
wire [MAX_SUM_WDTH_L-1:0]        Iacd3b2128fa021305b3de888d7612cf8;
wire [MAX_SUM_WDTH_L-1:0]        I96ef4b631a7f63e19f67f3920685f0e6;
wire [flogtanh_WDTH -1:0]        I2022005072d2979dae84b6e4491a3ce2;
wire [MAX_SUM_WDTH_L-1:0]        I0976b3262637cf38babc31162e3f6cea;
wire [MAX_SUM_WDTH_L-1:0]        I9e2de71442b8f504358e582087a6d19f;
wire [flogtanh_WDTH -1:0]        I98524ad028e4d832ebbcd92956dac08c;
wire [MAX_SUM_WDTH_L-1:0]        I484113b853de9a5684592b8318430da2;
wire [MAX_SUM_WDTH_L-1:0]        I1fb13d7500f5ac3821c424bd3688cf4e;
wire [flogtanh_WDTH -1:0]        I4d24e2ba47093eee6669f537374ecce7;
wire [MAX_SUM_WDTH_L-1:0]        I4b4a443a54b030b20a3e86ba0f63c1ee;
wire [MAX_SUM_WDTH_L-1:0]        I2aabda12ff89e708d04b4399472b5203;
wire [flogtanh_WDTH -1:0]        I227232e7189020459c16b3413e881b80;
wire [MAX_SUM_WDTH_L-1:0]        Ifb32581537c4402e5345932d83e1388f;
wire [MAX_SUM_WDTH_L-1:0]        I8c733a5d394e6b8d045eede5cc7451f6;
wire [flogtanh_WDTH -1:0]        If4359aebd4cc66c75cf2a44f681ccc72;
wire [MAX_SUM_WDTH_L-1:0]        Ib032b0c1073c1a3689b8f70a8a1f94b5;
wire [MAX_SUM_WDTH_L-1:0]        I4f45dd50d2825ab338b8a2a8264096c0;
wire [flogtanh_WDTH -1:0]        I8d2e10b8c474f1a915825ec78072ad56;
wire [MAX_SUM_WDTH_L-1:0]        I3ac6148b8dfcfb0816a01ff2a77b905d;
wire [MAX_SUM_WDTH_L-1:0]        Ib45caf6b563d22144be3e9225a99a1cd;
wire [flogtanh_WDTH -1:0]        Ie5b3748f3c81d9eeec767d546b29cbd8;
wire [MAX_SUM_WDTH_L-1:0]        Ie090d9460623450a9654f24bda1be1f7;
wire [MAX_SUM_WDTH_L-1:0]        I9d6730140c690037b5ca58aa30103f5b;
wire [flogtanh_WDTH -1:0]        Ib764a6d1978dc61cb4499b15c45cb1b4;
wire [MAX_SUM_WDTH_L-1:0]        I42979deb711e94d6a366a9c125277bc7;
wire [MAX_SUM_WDTH_L-1:0]        I9df5b63f66c162d517daa69f5d0e6095;
wire [flogtanh_WDTH -1:0]        I4fbe7db2d4288676183dc69ed56c9c68;
wire [MAX_SUM_WDTH_L-1:0]        I12b0827207c31ed0661711adddb9b59f;
wire [MAX_SUM_WDTH_L-1:0]        I1b40adfd6fa6c943dfa8d230d9e65514;
wire [flogtanh_WDTH -1:0]        I99f0cc5986099cb57fbebf9e5e262c56;
wire [MAX_SUM_WDTH_L-1:0]        If605c57ab8c22fa2cbb1e7f815274d80;
wire [MAX_SUM_WDTH_L-1:0]        I0eb3df4d4094e09e6c4b3c788baed61f;
wire [flogtanh_WDTH -1:0]        I4f5bb7e206563a334d7e2dd100b37c35;
wire [MAX_SUM_WDTH_L-1:0]        I82ed5aaddf52d30eba9c0116ef5e9a8c;
wire [MAX_SUM_WDTH_L-1:0]        Id6f7923a16cc5adc96a730083153ca6d;
wire [flogtanh_WDTH -1:0]        I59ecb14b5f34ebab3da4784709de66a4;
wire [MAX_SUM_WDTH_L-1:0]        I54e9afa2959a5a02f60ea11cfee788af;
wire [MAX_SUM_WDTH_L-1:0]        Idf8ebc0d747ae143aa61866e33d458c0;
wire [flogtanh_WDTH -1:0]        I54f5a8caf0e1c2df9477b37157d94995;
wire [MAX_SUM_WDTH_L-1:0]        I31b86d750f70d42455bd426e8d3e494f;
wire [MAX_SUM_WDTH_L-1:0]        Id682e531735437bc24abbf3d3d51e18b;
wire [flogtanh_WDTH -1:0]        I77e1bed2da0ccf1475dcfe908d64f82c;
wire [MAX_SUM_WDTH_L-1:0]        Ic2923e2c0a77b23dbe0724bf452ea190;
wire [MAX_SUM_WDTH_L-1:0]        I05ecce409cca00ea5b0df25de5a50cf2;
wire [flogtanh_WDTH -1:0]        I1a450ec193ccde2946f6ca20c0fa894c;
wire [MAX_SUM_WDTH_L-1:0]        Ie5fbbda327dbf0e90ad68ba42242fe21;
wire [MAX_SUM_WDTH_L-1:0]        I831d214dcb4f8d534b5ddaaeaeeb81ce;
wire [flogtanh_WDTH -1:0]        I01fbfc3b5c14733738f93a3487e54f35;
wire [MAX_SUM_WDTH_L-1:0]        I261e7001e9ca425607de438bef1f7f4d;
wire [MAX_SUM_WDTH_L-1:0]        Ia540866403683bc30504bace19bdda7b;
wire [flogtanh_WDTH -1:0]        Icff5d12020f78478c77210d9c692dfbe;
wire [MAX_SUM_WDTH_L-1:0]        I27aac717f95c8b5b7114810c77bb0761;
wire [MAX_SUM_WDTH_L-1:0]        I05fb1982415bd3fa78dd9a00af7a3d4a;
wire [flogtanh_WDTH -1:0]        I6eb28698ab4105a74c6510dbcfefbc3c;
wire [MAX_SUM_WDTH_L-1:0]        Id3820975eb9b8205aed04d02e9c21afb;
wire [MAX_SUM_WDTH_L-1:0]        I977864efb0d94149cce7dc4d165f11de;
wire [flogtanh_WDTH -1:0]        I7cc0f835ad7a18683e1fdb5bcbfb7f2f;
wire [MAX_SUM_WDTH_L-1:0]        Ifbd4c6cc29fdd08d49bd7fd9f68051b3;
wire [MAX_SUM_WDTH_L-1:0]        I9362b615a612599239e3b752a9334e8c;
wire [flogtanh_WDTH -1:0]        I9389a0dfe5a82a903c89e1a468f0ad57;
wire [MAX_SUM_WDTH_L-1:0]        I2e9993aa302580a47147469355f65dcf;
wire [MAX_SUM_WDTH_L-1:0]        I5d4fb4b5a5ad3dc48beebfa0e0cebbed;
wire [flogtanh_WDTH -1:0]        Idc4ce4afd846e212526d21a5e0cd1c14;
wire [MAX_SUM_WDTH_L-1:0]        I187d0d6496e96f11c9c2c241213d405e;
wire [MAX_SUM_WDTH_L-1:0]        Ifb9b29c43f435452cc761218c509f5df;
wire [flogtanh_WDTH -1:0]        I38a0ba1e69b467d4aed306e76ec3bfdb;
wire [MAX_SUM_WDTH_L-1:0]        I1fd12d5a4d0a5d8d08117f57f2f4880e;
wire [MAX_SUM_WDTH_L-1:0]        If2143db72bf9a02b64eb45b3a4faa39d;
wire [flogtanh_WDTH -1:0]        I66279b0fa707a272f43ee929cb297945;
wire [MAX_SUM_WDTH_L-1:0]        Iba9bee3dd12c2559872c8498e4cd6f2b;
wire [MAX_SUM_WDTH_L-1:0]        Ice780b1695a8e80607a03dee3c426ffe;
wire [flogtanh_WDTH -1:0]        Ib091954846c14743e01fd4e7bafda1b5;
wire [MAX_SUM_WDTH_L-1:0]        I8fecfe7601fa0d166db2b2fc9746129e;
wire [MAX_SUM_WDTH_L-1:0]        I90b0296f5ef87dfaa6110fc2e9d6ed9d;
wire [flogtanh_WDTH -1:0]        I3b8663f2adecb8da2c84dbb37341e25f;
wire [MAX_SUM_WDTH_L-1:0]        Ic3d6ada81005c125c29d8ff0abe88185;
wire [MAX_SUM_WDTH_L-1:0]        Icd37da8ea84a606529e32b2db4eb7f5f;
wire [flogtanh_WDTH -1:0]        I19bc03089c6c288e1778bd1f197a3ce3;
wire [MAX_SUM_WDTH_L-1:0]        Iddb333f6cb7253e92ba9e485a95c59c1;
wire [MAX_SUM_WDTH_L-1:0]        Ie626a24e3680f7d3995dd0c2ce60cbcc;
wire [flogtanh_WDTH -1:0]        I0988382a446b21da209d49d0d00bd6df;
wire [MAX_SUM_WDTH_L-1:0]        I64f8fb4dc07decbd4e91436847143c23;
wire [MAX_SUM_WDTH_L-1:0]        Iebee55168fb47664095b11c9f6641124;
wire [flogtanh_WDTH -1:0]        I19f5cb50b27b6c5e40012df9397aa288;
wire [MAX_SUM_WDTH_L-1:0]        I65c608dc3e2923360416cb08cfba6aeb;
wire [MAX_SUM_WDTH_L-1:0]        Ic0954671eb1dc893c3932e456800fadf;
wire [flogtanh_WDTH -1:0]        I706ca74386e5778b30eca35432429bc3;
wire [MAX_SUM_WDTH_L-1:0]        I70bae72ccecf63dd5a367bf40b4ac870;
wire [MAX_SUM_WDTH_L-1:0]        Ia4131464996aabab8aae1db85f6a50e4;
wire [flogtanh_WDTH -1:0]        If6af0cc7a120b2897c3a69d54a554e86;
wire [MAX_SUM_WDTH_L-1:0]        I32e73ad10e9df77b20d3eda78deeafac;
wire [MAX_SUM_WDTH_L-1:0]        I2de1ca2c390bdd3011fff4a359bb5332;
wire [flogtanh_WDTH -1:0]        I88ebe846173f486b07d2051a80bd055f;
wire [MAX_SUM_WDTH_L-1:0]        I4688025bd745934e70eaa03f3bb7d089;
wire [MAX_SUM_WDTH_L-1:0]        I6fb55222b69475b7168874423226ec9c;
wire [flogtanh_WDTH -1:0]        I2c577b130db6f4673704c858d454f3ea;
wire [MAX_SUM_WDTH_L-1:0]        I2c6ba69dd7827396366ce8e6513f8d4c;
wire [MAX_SUM_WDTH_L-1:0]        I9b09b800a9dcd8ac36f25cb0324e748d;
wire [flogtanh_WDTH -1:0]        I383f23d4e769bbdc1c8acd9c660a0b3e;
wire [MAX_SUM_WDTH_L-1:0]        Iecde1ff7e98a3f2aa847d1e55403f00f;
wire [MAX_SUM_WDTH_L-1:0]        I74ac0327175f50f508a5013df298df02;
wire [flogtanh_WDTH -1:0]        Iea20a6ecf4bbf907d1a102bde797284f;
wire [MAX_SUM_WDTH_L-1:0]        I28ae9c81892f556ffbc3ed65b7ec0fb5;
wire [MAX_SUM_WDTH_L-1:0]        Ica26f542586d50c56ce0f3c00f36b388;
wire [flogtanh_WDTH -1:0]        I77d655383c0c22b1af75d9308fab2e4f;
wire [MAX_SUM_WDTH_L-1:0]        I1bfb39b04609b92c72d95b724eb3cae0;
wire [MAX_SUM_WDTH_L-1:0]        I7c6862830daffc98cb2c1fc121d82c38;
wire [flogtanh_WDTH -1:0]        I4a4ebb2f3389d67c4b7671e12fc5cd92;
wire [MAX_SUM_WDTH_L-1:0]        I73ba173234b8583fa63ea947b5d2f957;
wire [MAX_SUM_WDTH_L-1:0]        Icf19dd665616a8c96146b3ab9f46c741;
wire [flogtanh_WDTH -1:0]        Ibc927d678e218397e23147b5c0654fd9;
wire [MAX_SUM_WDTH_L-1:0]        I9f0cce614937f873f39006b334729d72;
wire [MAX_SUM_WDTH_L-1:0]        I97f2813ec39bbf1513faf66b3e38838a;
wire [flogtanh_WDTH -1:0]        Ib0358b6f47edcd54971935de215203f8;
wire [MAX_SUM_WDTH_L-1:0]        I129867553993fbc89983071472910fa4;
wire [MAX_SUM_WDTH_L-1:0]        I716ee53e79883f69aa045380a357e913;
wire [flogtanh_WDTH -1:0]        Iaa6f2bbd8a343ebf878da57badb4572b;
wire [MAX_SUM_WDTH_L-1:0]        I2d6c9368bf6cc6e58ea202397528a736;
wire [MAX_SUM_WDTH_L-1:0]        I25c324feaca84e80f58075597e8c448f;
wire [flogtanh_WDTH -1:0]        I823f1a0d2d757d5ca83dc7b5ca08e0f8;
wire [MAX_SUM_WDTH_L-1:0]        I715eedae273662cb8417d53b77f280c2;
wire [MAX_SUM_WDTH_L-1:0]        I7fc190647082a3d71614f46f670167bc;
wire [flogtanh_WDTH -1:0]        I1a650234a61a3ff90ea079e29d322069;
wire [MAX_SUM_WDTH_L-1:0]        Iab6f27ce8700543dfb7a8005ae320445;
wire [MAX_SUM_WDTH_L-1:0]        Iebdf938a28594624f4d4a337356485cb;
wire [flogtanh_WDTH -1:0]        I70a7b1083c9593840759854430ee9d62;
wire [MAX_SUM_WDTH_L-1:0]        Iaf6ebea4db33923d6db2c721d1dcd0d4;
wire [MAX_SUM_WDTH_L-1:0]        I3fd068d55154441ffd005999ea823fd0;
wire [flogtanh_WDTH -1:0]        I99aa55a3e285e62e9a8b50174e84b68c;
wire [MAX_SUM_WDTH_L-1:0]        Ic17b627fb3201547b05b457648431ad5;
wire [MAX_SUM_WDTH_L-1:0]        Ic5ca74b66763c6e5591c7c2bfeeb0663;
wire [flogtanh_WDTH -1:0]        Ief099d2084b84e0e23599d98102a13b7;
wire [MAX_SUM_WDTH_L-1:0]        Iee1fb0a6e0aceddc45640b7ea4b4d0cd;
wire [MAX_SUM_WDTH_L-1:0]        I5ab556386d2973354a5551ba9823e4ba;
wire [flogtanh_WDTH -1:0]        I84aa89bab681c2fc7a8c7c6b47200dec;
wire [MAX_SUM_WDTH_L-1:0]        I851d25c73aa5ee6bb26c0435353af3b8;
wire [MAX_SUM_WDTH_L-1:0]        I64f65df774d29696425ba460dda09b68;
wire [flogtanh_WDTH -1:0]        I101b9397639b59fd53a88d17425e0c96;
wire [MAX_SUM_WDTH_L-1:0]        I35e97af89c2791175cc545646eb7ba92;
wire [MAX_SUM_WDTH_L-1:0]        I9e09c25be9f877c1e1aaf79bf12c7943;
wire [flogtanh_WDTH -1:0]        Ic302f050dba883d8f4bd20b1030ba14d;
wire [MAX_SUM_WDTH_L-1:0]        I99b5120e2171e49d3320913b9e372936;
wire [MAX_SUM_WDTH_L-1:0]        I42c1d469ff97913cbf15e3ebee6fdfa8;
wire [flogtanh_WDTH -1:0]        I848425f041888d7433b68900f259732a;
wire [MAX_SUM_WDTH_L-1:0]        Idb7353d31a0038c904c4e25c78be46a5;
wire [MAX_SUM_WDTH_L-1:0]        If9f2a53dbf6e9b9a335a7657b7a2b468;
wire [flogtanh_WDTH -1:0]        I2b4671193178503f5329954e74a399b3;
wire [MAX_SUM_WDTH_L-1:0]        I17ae1aa33db4ca2948befb43f1bd3d06;
wire [MAX_SUM_WDTH_L-1:0]        I495f8be463b15db906474c518e0741e2;
wire [flogtanh_WDTH -1:0]        I97b93c6d963d51a819b1dc9ab3bf28ea;
wire [MAX_SUM_WDTH_L-1:0]        Ida342ed2e96314bb7c0182b3d895b647;
wire [MAX_SUM_WDTH_L-1:0]        I3e265a7dcf29687248b9275df49771fb;
wire [flogtanh_WDTH -1:0]        I2593b1b30f4c97845a1f77c3f558b263;
wire [MAX_SUM_WDTH_L-1:0]        If1d8968112c433d9d9bb309cc916fec9;
wire [MAX_SUM_WDTH_L-1:0]        Iffd94cf3a8a4681ff3327c90bf89bd8b;
wire [flogtanh_WDTH -1:0]        I3a4695c79b62f6baa47cdc939c4e2974;
wire [MAX_SUM_WDTH_L-1:0]        I6a927fb5af8b12fcd5d5b1b2b4e1f4b5;
wire [MAX_SUM_WDTH_L-1:0]        Iea71417e738c6ca54c50aa014cc38627;
wire [flogtanh_WDTH -1:0]        Ibc577b2948aec87c0696c860d7efa1d7;
wire [MAX_SUM_WDTH_L-1:0]        Ic6b949621a3f4c61ac219919731f8f83;
wire [MAX_SUM_WDTH_L-1:0]        Ic8df04756f67e6dd29f3374c5f86d451;
wire [flogtanh_WDTH -1:0]        I08401e4e9a1766a0034f45933b5bb29a;
wire [MAX_SUM_WDTH_L-1:0]        Ie8bfce645fef58bf090818dce30d86e4;
wire [MAX_SUM_WDTH_L-1:0]        I546122346a22ad64a6ab2b4978cde095;
wire [flogtanh_WDTH -1:0]        I5e5bb0de4fe6682a6beaa86f6cd1ca32;
wire [MAX_SUM_WDTH_L-1:0]        Ide2a4d41e8d2871f7c52249a8cb48ac1;
wire [MAX_SUM_WDTH_L-1:0]        Icaae0fb0f460f68d690ab00697355a49;
wire [flogtanh_WDTH -1:0]        Ia487e80f0010e7cb34aa12471e62a62f;
wire [MAX_SUM_WDTH_L-1:0]        Ib58e63392e279cbb87c4e5be4e4b0109;
wire [MAX_SUM_WDTH_L-1:0]        I42455e7e4d0c63f97702d204d18a446e;
wire [flogtanh_WDTH -1:0]        I3bee9305e2f4456aae800bbb174b7843;
wire [MAX_SUM_WDTH_L-1:0]        Ic680a004d350df1379eddb3ed06be34e;
wire [MAX_SUM_WDTH_L-1:0]        Iaec2f15665e83416bc140890f3cdde9a;
wire [flogtanh_WDTH -1:0]        I14f1aa0dbf6f1f0fbf6b5f996e229a04;
wire [MAX_SUM_WDTH_L-1:0]        I8074f2ecf0e4178d0b8d58f4d6680282;
wire [MAX_SUM_WDTH_L-1:0]        I487391402b6aa27bf212724a37ea9c33;
wire [flogtanh_WDTH -1:0]        If87afc1cf342dca9986f798c38a69dab;
wire [MAX_SUM_WDTH_L-1:0]        I20b0882e61c68796b057b0a9d237a979;
wire [MAX_SUM_WDTH_L-1:0]        Ia9f375709014a9d553d46cff2799b59f;
wire [flogtanh_WDTH -1:0]        Ibb1c020ea255a966e54c00fc7cc745b5;
wire [MAX_SUM_WDTH_L-1:0]        I4c1ecb851699ea3c2642c78fa44b04e6;
wire [MAX_SUM_WDTH_L-1:0]        I34d428a56bd0142a9be9f627f1c3c87f;
wire [flogtanh_WDTH -1:0]        Icae8a2980dd7403caf72820ae508885b;
wire [MAX_SUM_WDTH_L-1:0]        I421cb46488584e6314f701cfe34d3e79;
wire [MAX_SUM_WDTH_L-1:0]        I57db98eb439d59a895dabe029c6a3a8b;
wire [flogtanh_WDTH -1:0]        Ic8f858d7f7a16b771933741d31679dc1;
wire [MAX_SUM_WDTH_L-1:0]        Ibed20c973d23c4058efffc1575d66478;
wire [MAX_SUM_WDTH_L-1:0]        I9937af6fcf9d834f308bc3683d524981;
wire [flogtanh_WDTH -1:0]        I9dcf19da38f352fe7fa27c22bff08c19;
wire [MAX_SUM_WDTH_L-1:0]        I2f5e17be80bab46917da109cf7ac3532;
wire [MAX_SUM_WDTH_L-1:0]        I463f4f370e1ecad71de44780eff10df4;
wire [flogtanh_WDTH -1:0]        I2bc787aa749db4a5f48bd917715a11d5;
wire [MAX_SUM_WDTH_L-1:0]        I43b6cac96c5c2236629f6ee87f13e0be;
wire [MAX_SUM_WDTH_L-1:0]        I53309409a6059c3bd39f037c23ec3458;
wire [flogtanh_WDTH -1:0]        I3d072e173fd12ac9d802a29a0ff4378c;
wire [MAX_SUM_WDTH_L-1:0]        I54a8f8a82aa219427914ca74da599696;
wire [MAX_SUM_WDTH_L-1:0]        I2603e0b8b93f6680e44c9c8883f6512c;
wire [flogtanh_WDTH -1:0]        I2115d62275a57ec7273e3631c0a32872;
wire [MAX_SUM_WDTH_L-1:0]        I23e89a266dd6a09d486b129eea48fae5;
wire [MAX_SUM_WDTH_L-1:0]        Iab354cc9ac1173335c0efeef694f3567;
wire [flogtanh_WDTH -1:0]        I91bc663fcd7f86a066b8b3f93b1dcfc2;
wire [MAX_SUM_WDTH_L-1:0]        I8b68b47c8e9b4055b176745aec55b3b2;
wire [MAX_SUM_WDTH_L-1:0]        I6c19936ca2edeb0e261e880a1055e964;
wire [flogtanh_WDTH -1:0]        I988c0d94f97329dd1cff7d913cb449e7;
wire [MAX_SUM_WDTH_L-1:0]        I1195ee9289f2afca25519bb6d493e73a;
wire [MAX_SUM_WDTH_L-1:0]        Ifebfa58419ecd22a334ed4b67f5c3581;
wire [flogtanh_WDTH -1:0]        If444a37a85774dcc2769ffd74b785e46;
wire [MAX_SUM_WDTH_L-1:0]        I2844ec353c6ac19013e7a64d350f0204;
wire [MAX_SUM_WDTH_L-1:0]        I71a28e8525f07dabeabe4b4f45f353d0;
wire [flogtanh_WDTH -1:0]        Idbb89639b8399b57b190efd898643328;
wire [MAX_SUM_WDTH_L-1:0]        Ie4848a127b84c06712bd2b40d80b214d;
wire [MAX_SUM_WDTH_L-1:0]        I514830acdad20c4ff3d078477e939b4b;
wire [flogtanh_WDTH -1:0]        Ib1d70f302858eb7c78fb834071616a9b;
wire [MAX_SUM_WDTH_L-1:0]        Id93016d32ebfabc6e464df96ae3aa74c;
wire [MAX_SUM_WDTH_L-1:0]        I036342f6be0f2e2f1f4927099a5c4a78;
wire [flogtanh_WDTH -1:0]        I82bd4ea32da7ae3a0d5938fc8a1424c5;
wire [MAX_SUM_WDTH_L-1:0]        I0ed0efac703623c9a35ffb79a57683dc;
wire [MAX_SUM_WDTH_L-1:0]        Iedb655aa25e5f0e35137ec6c3acdc527;
wire [flogtanh_WDTH -1:0]        I6964f2e681e9cdf63fbc0358cb6edcca;
wire [MAX_SUM_WDTH_L-1:0]        I2f1a1b3caf70a00d30678c22f68f9cfe;
wire [MAX_SUM_WDTH_L-1:0]        I0c59e8c82a31aacbf5977ff778a7ff49;
wire [flogtanh_WDTH -1:0]        I41aeb75239ce0d636288e8ceb0665b34;
wire [MAX_SUM_WDTH_L-1:0]        I8acdcab405f76f4bf751e8860a50e614;
wire [MAX_SUM_WDTH_L-1:0]        I1b6d20c64b9f23fb6c30f723546aa285;
wire [flogtanh_WDTH -1:0]        Ie0d3fd5e7c38c10fdcae3f1b217c28f4;
wire [MAX_SUM_WDTH_L-1:0]        I88ede5095d3876c7ca6dac02faa3eede;
wire [MAX_SUM_WDTH_L-1:0]        I0d66aa55747362354aa81d96057bc4c2;
wire [flogtanh_WDTH -1:0]        Ia8b7d74eaf227e697c3eb58b31eb355f;
wire [MAX_SUM_WDTH_L-1:0]        I68bc064fabdc9564021be1d29f3cbb7a;
wire [MAX_SUM_WDTH_L-1:0]        I1ea33707e40a2e41513fdb3118371437;
wire [flogtanh_WDTH -1:0]        I79034cd4180d03348de2c101927048a7;
wire [MAX_SUM_WDTH_L-1:0]        Idfd56dd8b81f3ec49acfa9131d4b78c4;
wire [MAX_SUM_WDTH_L-1:0]        I68c85727adecde0aa8aa66ed08c4b502;
wire [flogtanh_WDTH -1:0]        Id23895e0696cdd27e3087294fb52a65b;
wire [MAX_SUM_WDTH_L-1:0]        I777937fc3cbdcb60a10ee0c0d1f56dc5;
wire [MAX_SUM_WDTH_L-1:0]        Iebd050e29044153d5881ef80b2db8c28;
wire [flogtanh_WDTH -1:0]        I43939a168f9f5e476262ace39c6ae483;
wire [MAX_SUM_WDTH_L-1:0]        I2de42de0be5ebc2ee41fb217953cb823;
wire [MAX_SUM_WDTH_L-1:0]        I3c057d64cf4fca0238a874f0ced99c76;
wire [flogtanh_WDTH -1:0]        Ie5167faac3e6510d4b208a1bdc0cd44c;
wire [MAX_SUM_WDTH_L-1:0]        Ied21906ec121c7c7da1d0268e93ab0a6;
wire [MAX_SUM_WDTH_L-1:0]        I066cd52173ec5dbce9a3f470d73325af;
wire [flogtanh_WDTH -1:0]        I1cad8b885a541dd049093ce60c3f8a06;
wire [MAX_SUM_WDTH_L-1:0]        I074d42d6f79dd8786745ad7b0f59b3e5;
wire [MAX_SUM_WDTH_L-1:0]        Ic7ad59f6a232a997706d17b4098e0324;
wire [flogtanh_WDTH -1:0]        Icd2d69f12d4744ce7b09fce7f27ab830;
wire [MAX_SUM_WDTH_L-1:0]        I78cfd6df12d7b773c498ed763953c8a2;
wire [MAX_SUM_WDTH_L-1:0]        Icf8cfc800f0a2aa5140a7f83f035b0cc;
wire [flogtanh_WDTH -1:0]        Ic9ee0243e36f66f462eb3d4ce93fdde9;
wire [MAX_SUM_WDTH_L-1:0]        I3e452666c55d9b30beef77c58690c8fd;
wire [MAX_SUM_WDTH_L-1:0]        I6bfbf7ff79ff0a6facc9ba5031239644;
wire [flogtanh_WDTH -1:0]        I5353c3239ddb4d7fa7094e413b5303b1;
wire [MAX_SUM_WDTH_L-1:0]        I5524ea6d4e43842521569ba37425b387;
wire [MAX_SUM_WDTH_L-1:0]        I78ade92efd265027807c861be44a10af;
wire [flogtanh_WDTH -1:0]        Idfca1b1d8041e5808799499e8c8dcf5e;
wire [MAX_SUM_WDTH_L-1:0]        I8153350f4b99d2a42acc18f730911337;
wire [MAX_SUM_WDTH_L-1:0]        I2bc5a10c587d89d10021aa5eaafb490a;
wire [flogtanh_WDTH -1:0]        I4710d61c763098027934286c6a9f3714;
wire [MAX_SUM_WDTH_L-1:0]        I685829af9b536012f05d3a22e0d7651b;
wire [MAX_SUM_WDTH_L-1:0]        I30080cc6c03bbe933165d266558a822c;
wire [flogtanh_WDTH -1:0]        If6a04c29b7205c5db5f2ff3cf302c45f;
wire [MAX_SUM_WDTH_L-1:0]        Ibb607d3707048ec1dd1f126852667fcb;
wire [MAX_SUM_WDTH_L-1:0]        I7e28234bdf66ab5489d36d15678db797;
wire [flogtanh_WDTH -1:0]        Ib5d9348a114627a8b1f56aca968d20b1;
wire [MAX_SUM_WDTH_L-1:0]        Ib948458593df6c9b4bef35c88845492d;
wire [MAX_SUM_WDTH_L-1:0]        I74b3c9dd3a8168aacd4369b9ff68fdfd;
wire [flogtanh_WDTH -1:0]        I4e2b59a03731959106d469ffee7b7d33;
wire [MAX_SUM_WDTH_L-1:0]        Ifbebc06fa0ddc76aa8053ee669fda467;
wire [MAX_SUM_WDTH_L-1:0]        Ia7046faae1ab05978e4b32bd44049fb9;
wire [flogtanh_WDTH -1:0]        Ic6d519691c7543b1bd0707a8c9899088;
wire [MAX_SUM_WDTH_L-1:0]        I059d9b49b8c6de67643992e5ef74d939;
wire [MAX_SUM_WDTH_L-1:0]        I0c5250aaca86185fed5978438c8861b6;
wire [flogtanh_WDTH -1:0]        Icc6bde490bd8df2ce5efe8cfb24cf5f5;
wire [MAX_SUM_WDTH_L-1:0]        I141b6f8e6baa353f2527dc1171c95908;
wire [MAX_SUM_WDTH_L-1:0]        Ic78949e07e643f571f23df7e8f15d9fb;
wire [flogtanh_WDTH -1:0]        I861bd8df5caf968dc6edd7a05d690033;
wire [MAX_SUM_WDTH_L-1:0]        I891992837c6e3d393516506efec821e1;
wire [MAX_SUM_WDTH_L-1:0]        Ifb8b3586a5b69b20cf03eabf51344ab6;
wire [flogtanh_WDTH -1:0]        I6f44882493f9eadbdbe1ac46a3d2a43b;
wire [MAX_SUM_WDTH_L-1:0]        I9739e5853bd26c50167491b69e92ed6f;
wire [MAX_SUM_WDTH_L-1:0]        I9ea09f27ce4484f2e7fc3a6b6d6ecb7c;
wire [flogtanh_WDTH -1:0]        I5a3ec39885fba8d015009d671a1cb544;
wire [MAX_SUM_WDTH_L-1:0]        I80c41a49bba592ec70c6ca394bb48845;
wire [MAX_SUM_WDTH_L-1:0]        If0b9225e759438be175c4128c78605ea;
wire [flogtanh_WDTH -1:0]        Ic4e6d76148a8170d1af0c95f370367a5;
wire [MAX_SUM_WDTH_L-1:0]        Ia96cc576fbc424161dcc350151e4476d;
wire [MAX_SUM_WDTH_L-1:0]        I33d941ad9d4858fcfb77f0f6cf99d2ec;
wire [flogtanh_WDTH -1:0]        I244bd772f9d750b4e1800e0b0ca67d63;
wire [MAX_SUM_WDTH_L-1:0]        I3abbd492752bc871096dac47e3208d01;
wire [MAX_SUM_WDTH_L-1:0]        Ia0868eee7e7e0640ce1a4d3ca9c001cb;
wire [flogtanh_WDTH -1:0]        I00c203d60e09f1cccdadb8ebff2de650;
wire [MAX_SUM_WDTH_L-1:0]        Iff5e7ff31a18e5a3947f16c456cb4bf2;
wire [MAX_SUM_WDTH_L-1:0]        Icb3ab2c67a87b2ee158e0021b72fc186;
wire [flogtanh_WDTH -1:0]        I20c7780e77b49d31808e59cae58968a9;
wire [MAX_SUM_WDTH_L-1:0]        I6f437a921b54934b3a5d13eb2d8e4b5e;
wire [MAX_SUM_WDTH_L-1:0]        I5b64997d083769666741c794dd92fb7f;
wire [flogtanh_WDTH -1:0]        Ia332fad029505e5975156f8e13910358;
wire [MAX_SUM_WDTH_L-1:0]        Ieb8e5fdc6ac722d69775b46b0f081bf7;
wire [MAX_SUM_WDTH_L-1:0]        I0a3323aac825506435068f6746aee974;
wire [flogtanh_WDTH -1:0]        I9cc95185621ad5718a905092c03315f8;
wire [MAX_SUM_WDTH_L-1:0]        I8b60818e4831ff872dd58accdbe94b30;
wire [MAX_SUM_WDTH_L-1:0]        Ibec442c099da091afcf75a7c970bf8ea;
wire [flogtanh_WDTH -1:0]        Iba2a341076f0506aeac3769e71b91f43;
wire [MAX_SUM_WDTH_L-1:0]        I9e1401baae9fab762f3ac1382b4658ed;
wire [MAX_SUM_WDTH_L-1:0]        If3a79ede332c39a8d2a276de833242f6;
wire [flogtanh_WDTH -1:0]        Ic9e82f153d0e690d5ea47ee159523b72;
wire [MAX_SUM_WDTH_L-1:0]        I19e98430858ce2db7853b31e4a8409f0;
wire [MAX_SUM_WDTH_L-1:0]        I49ccb3e14fe61618806e791ecb4f4eae;
wire [flogtanh_WDTH -1:0]        Ia265b95249953a7867c611d475d01169;
wire [MAX_SUM_WDTH_L-1:0]        I58ed96e69f7ce8d98d44b992f52fe7ca;
wire [MAX_SUM_WDTH_L-1:0]        I461ebbf3a02ae63e2eb27531b1370f24;
wire [flogtanh_WDTH -1:0]        I5ef2899606d7f08aa6d0028f9f113e38;
wire [MAX_SUM_WDTH_L-1:0]        Ie2b3c1982842e9b4f2befd0fce03a1cf;
wire [MAX_SUM_WDTH_L-1:0]        Ice66c108aa66981051df71e226cb0e4d;
wire [flogtanh_WDTH -1:0]        Idf3a6723fec1ef62c1e37a419590122c;
wire [MAX_SUM_WDTH_L-1:0]        I1a66d7f556b0f90b7f7c1321d1998cc3;
wire [MAX_SUM_WDTH_L-1:0]        I645ff0d8c0a87ba7f792fc83f342b958;
wire [flogtanh_WDTH -1:0]        I0bde2fc197586c74374ffb402956baf5;
wire [MAX_SUM_WDTH_L-1:0]        I87ace9b2a7e2e5ced87a85ad45c0b0c9;
wire [MAX_SUM_WDTH_L-1:0]        Ica94017f26e96fb22a47add326ee126e;
wire [flogtanh_WDTH -1:0]        I9182b3349816b6ddaffde1cbec78339e;
wire [MAX_SUM_WDTH_L-1:0]        Ia51a22a9b78f5e3e8b6e86b919ceb13d;
wire [MAX_SUM_WDTH_L-1:0]        Id32e7ad5b1aa825732d9b26d0fa02ca1;
wire [flogtanh_WDTH -1:0]        I5bf9702e2afd6c791b28c76c84aeb886;
wire [MAX_SUM_WDTH_L-1:0]        Ibb6b016405d27b6863c2d182e9465a5e;
wire [MAX_SUM_WDTH_L-1:0]        I51b5e641856239367cf43f9b5679b268;
wire [flogtanh_WDTH -1:0]        Ifbd7b868d9cb7e04bf2189922bcb9c92;
wire [MAX_SUM_WDTH_L-1:0]        I2bd977c2b670677802c6486507b0672f;
wire [MAX_SUM_WDTH_L-1:0]        I2d1a5645b126761fc7fb70d24e37189a;
wire [flogtanh_WDTH -1:0]        Ib78e7602e521bc064d5cd9efe10ec6b1;
wire [MAX_SUM_WDTH_L-1:0]        Ie9cd522fdd4e6e94287e7a8ce329c31e;
wire [MAX_SUM_WDTH_L-1:0]        I49f5f87662fbb540d72c94bfd1acd060;
wire [flogtanh_WDTH -1:0]        I0497115b3dd67c6538039969368e03ae;
wire [MAX_SUM_WDTH_L-1:0]        I1330526fdd2ffaa0137d4735167961b5;
wire [MAX_SUM_WDTH_L-1:0]        I30253dc91301ca27b5732312c01145e0;
wire [flogtanh_WDTH -1:0]        Ieba8e28ee660b8e2d78909d61ced3233;
wire [MAX_SUM_WDTH_L-1:0]        Ib9939f977a24ec96a60403bc4e8d4ef3;
wire [MAX_SUM_WDTH_L-1:0]        I143f5e324716a94d24ada126886bf895;
wire [flogtanh_WDTH -1:0]        I12e6fe32f6159ce6bb8be6411af2b7bb;
wire [MAX_SUM_WDTH_L-1:0]        I6d268ba2240ef4c0ac98f5e771964820;
wire [MAX_SUM_WDTH_L-1:0]        If64aa8c220b9ab6652e081da7e404e80;
wire [flogtanh_WDTH -1:0]        I03392e42f99b06cb65b38122c1e4dc81;
wire [MAX_SUM_WDTH_L-1:0]        If6639d10ed80985c8e322a85cfe65887;
wire [MAX_SUM_WDTH_L-1:0]        I1092325b801600fa7ec85fa640167da9;
wire [flogtanh_WDTH -1:0]        I32270eb6cf0594020ee19abb2edfe93d;
wire [MAX_SUM_WDTH_L-1:0]        I5d4d3b9363d24d988468d1782347a41c;
wire [MAX_SUM_WDTH_L-1:0]        Ib028686da9c849e827cf249a744b7db3;
wire [flogtanh_WDTH -1:0]        Ib135d3d7d338f5ff3a1f504aec754bbd;
wire [MAX_SUM_WDTH_L-1:0]        I6461781f905b7694ad26c54d6f8cb062;
wire [MAX_SUM_WDTH_L-1:0]        I5f3ff7fa8686f7a380302d71b88cfb4b;
wire [flogtanh_WDTH -1:0]        Id9cbc2e4b0f437840f028c7273d49416;
wire [MAX_SUM_WDTH_L-1:0]        I731ddcd050cee04fdfd5724c7236e9fb;
wire [MAX_SUM_WDTH_L-1:0]        Ic01904f7c518990eff2dc1de127676c4;
wire [flogtanh_WDTH -1:0]        I98b5a84c247422b51abf63a705fbb5f7;
wire [MAX_SUM_WDTH_L-1:0]        I0306fc584747e83ab0f2be50b228a1ad;
wire [MAX_SUM_WDTH_L-1:0]        I43f2ddd9780f86af489f8deae51168ec;
wire [flogtanh_WDTH -1:0]        I0ae39e89061b4f8c5c0e56eba2f48889;
wire [MAX_SUM_WDTH_L-1:0]        I7b2920a709b708955c261faa5ffda88c;
wire [MAX_SUM_WDTH_L-1:0]        I0a013fff6c792363bd7feb03d9691db8;
wire [flogtanh_WDTH -1:0]        If612cf94a3cefcfb844d6e975ba4aada;
wire [MAX_SUM_WDTH_L-1:0]        Iae6e4e88f9136c6c09f4fe0c9825e2e0;
wire [MAX_SUM_WDTH_L-1:0]        I7cf8401bf6893eab0b9f33a0f91ddd05;
wire [flogtanh_WDTH -1:0]        I3dab04eb1045e1b3b6bb47e0f4c390ad;
wire [MAX_SUM_WDTH_L-1:0]        Ic729485a48ee429c62eab4aef90b03b8;
wire [MAX_SUM_WDTH_L-1:0]        Ic7ccbeaf4ab94d0660eb7a0533723e24;
wire [flogtanh_WDTH -1:0]        I447db5cb14c9588418037bbb793a6274;
wire [MAX_SUM_WDTH_L-1:0]        I009290dfe067ac2cc190b53a07374b34;
wire [MAX_SUM_WDTH_L-1:0]        I08043393cb7f2558c145a698ea6652c9;
wire [flogtanh_WDTH -1:0]        Ic1227b130f19411495bed64035ea317b;
wire [MAX_SUM_WDTH_L-1:0]        I97455c455bbd84f8085f827abe335a75;
wire [MAX_SUM_WDTH_L-1:0]        I84865c4f872c0845124b78fabf695c2c;
wire [flogtanh_WDTH -1:0]        I6861b48d33277dd057c6f09ba630d700;
wire [MAX_SUM_WDTH_L-1:0]        I89efdab57b5f47e1ff25b260a26b7ce0;
wire [MAX_SUM_WDTH_L-1:0]        I57b9dd7a7deea6695dcd03439c9723cf;
wire [flogtanh_WDTH -1:0]        I022bebca44e2f0b8f9877dd0e709b29f;
wire [MAX_SUM_WDTH_L-1:0]        I9f27d55531f208c5e3b038a7e263fc48;
wire [MAX_SUM_WDTH_L-1:0]        I1cd6b35bcdfd461db69a4c1bdb1d387f;
wire [flogtanh_WDTH -1:0]        I8e3d5a48955fe19e24975579d55f4e14;
wire [MAX_SUM_WDTH_L-1:0]        Ib61c6917f61d77ed3c4a7cccf800147a;
wire [MAX_SUM_WDTH_L-1:0]        I40a1ecabded8add5bffe316f2d8beda9;
wire [flogtanh_WDTH -1:0]        I7ee915ffb1c7b8985788c5e6af532ce3;
wire [MAX_SUM_WDTH_L-1:0]        Id6b11b9d84008c2444e2d5bd86e5415d;
wire [MAX_SUM_WDTH_L-1:0]        I7c52ae4af926267b5e27a530202fcce0;
wire [flogtanh_WDTH -1:0]        Ia897087d82c2deac4697755c31766241;
wire [MAX_SUM_WDTH_L-1:0]        I3ee69feaef543b025d4267eb09c2cde9;
wire [MAX_SUM_WDTH_L-1:0]        I1a5c6c50817db8bde279d5f0b5095d76;
wire [flogtanh_WDTH -1:0]        I4c23326dc80b54231289f9f18c4db711;
wire [MAX_SUM_WDTH_L-1:0]        I7ebbfe102249fcdd69f0088cd52a1fbb;
wire [MAX_SUM_WDTH_L-1:0]        Idf0c1b85712fcbbbcc12915158ebff62;
wire [flogtanh_WDTH -1:0]        I8326b063a9b9688fb3014667c49ada1b;
wire [MAX_SUM_WDTH_L-1:0]        Ic50e81e4594d56cfd739f7f9791b1e15;
wire [MAX_SUM_WDTH_L-1:0]        I6b32298e8c61e75d0a38bca3084c0528;
wire [flogtanh_WDTH -1:0]        Ic41133a438fcea4a1cad9f5e5ee05a03;
wire [MAX_SUM_WDTH_L-1:0]        I2968c281ccf212e6a4d456ef3e6a820e;
wire [MAX_SUM_WDTH_L-1:0]        I5b0d72cedc120406402076148e2d30b0;
wire [flogtanh_WDTH -1:0]        I1ac5e426032b874b250cb8adad5b345a;
wire [MAX_SUM_WDTH_L-1:0]        Idd368451dfa1cd543cc66f44f3def824;
wire [MAX_SUM_WDTH_L-1:0]        Iaf624549f73b0d13c1a73c850b99f810;
wire [flogtanh_WDTH -1:0]        If9aca7e28f987bf6c7f2fb9b6f11962f;
wire [MAX_SUM_WDTH_L-1:0]        Ib979f9151b0b4c7c6e850780ce01cd5c;
wire [MAX_SUM_WDTH_L-1:0]        Iaaf7efeae9f6dc9e8222dc2b10122000;
wire [flogtanh_WDTH -1:0]        Id98a58cd8017fd149ea4f5b295f7ec80;
wire [MAX_SUM_WDTH_L-1:0]        Ie3b60e864d739cc4d2c015bc0e4d85ed;
wire [MAX_SUM_WDTH_L-1:0]        Iea1cd2321d2ac9b891b344e2ba2363d3;
wire [flogtanh_WDTH -1:0]        Ib9e45e75ce8cdd3b548eaf3e41a091ce;
wire [MAX_SUM_WDTH_L-1:0]        Id80fb022cc3ea4d663506b98ead354a4;
wire [MAX_SUM_WDTH_L-1:0]        Ia544fa24b953fe91800978895e3e610e;
wire [flogtanh_WDTH -1:0]        I9fcedcbd532cefe1e66ec94b22457cf4;
wire [MAX_SUM_WDTH_L-1:0]        I25fc15d8cb0faffee2dd7aadf733ac0e;
wire [MAX_SUM_WDTH_L-1:0]        I7fa710c37f5f96c3cdc35612a702a71c;
wire [flogtanh_WDTH -1:0]        Ic627802cf228a709638c14adf83091f8;
wire [MAX_SUM_WDTH_L-1:0]        I343f01a96adfc2286191f40a13d92ebf;
wire [MAX_SUM_WDTH_L-1:0]        I98fd105696fca11c1075f9bd30013747;
wire [flogtanh_WDTH -1:0]        Ib6bd27a683e11d238fcb775bb44dd913;
wire [MAX_SUM_WDTH_L-1:0]        Iab18cb1f98768ce17f46117b9a72090a;
wire [MAX_SUM_WDTH_L-1:0]        I61345963ceabdaa0f25f8a463fc9fe5d;
wire [flogtanh_WDTH -1:0]        I3affcbe66b25dc7f11f98b4e444937a2;
wire [MAX_SUM_WDTH_L-1:0]        Icd8c66b0c9d66db6764cc3566a14cf06;
wire [MAX_SUM_WDTH_L-1:0]        I9e8375af6af10f4bac3e87e416d430ee;
wire [flogtanh_WDTH -1:0]        Ib537657951962c85ad92d43777458588;
wire [MAX_SUM_WDTH_L-1:0]        I51c808cc77479f221a7c60486b75f6ed;
wire [MAX_SUM_WDTH_L-1:0]        Ida1cd844022bbf1b8431225e66b2b78f;
wire [flogtanh_WDTH -1:0]        Id0af2b1d8b0aa3ba9764ea6a22fafc8c;
wire [MAX_SUM_WDTH_L-1:0]        I18a65513ce78aa9c77275103956df746;
wire [MAX_SUM_WDTH_L-1:0]        I30e9ab592e97dbc5fb6ab58d2ffbf8d4;
wire [flogtanh_WDTH -1:0]        I3f934c17beeba9f2d2ca58b3677fe1f3;
wire [MAX_SUM_WDTH_L-1:0]        I004491418434bb0a6a307d305df7dab0;
wire [MAX_SUM_WDTH_L-1:0]        I2ec2a6de2be39b1bc259b0be72e35a0f;
wire [flogtanh_WDTH -1:0]        Ie3e094ae62dc2a694777f4792c78c886;
wire [MAX_SUM_WDTH_L-1:0]        Ia74f2ce0e44e31217be3962f40588238;
wire [MAX_SUM_WDTH_L-1:0]        Ic32e349efae2ca419e095ee5e15a501d;
wire [flogtanh_WDTH -1:0]        Idea1d2f5e910ebadc99d356dee8646bd;
wire [MAX_SUM_WDTH_L-1:0]        Ic92636db4722431041a6b48e99b5924d;
wire [MAX_SUM_WDTH_L-1:0]        I1befb935ee9cb871c9a7476c1fc0da3f;
wire [flogtanh_WDTH -1:0]        I7cf160bea55d67417a4ee9ce9b252871;
wire [MAX_SUM_WDTH_L-1:0]        Ib525e226298f02a92a49a6fe5fcf6527;
wire [MAX_SUM_WDTH_L-1:0]        I01c57f697f2af7d2c6ae904319f10725;
wire [flogtanh_WDTH -1:0]        I196915263bfb62cc21659f81572438b4;
wire [MAX_SUM_WDTH_L-1:0]        Icefd1ea8daf4aaf25abd3b31256dcaa5;
wire [MAX_SUM_WDTH_L-1:0]        Id580f8a2748efff9b6b747c497c16e9c;
wire [flogtanh_WDTH -1:0]        I548af5c4ccd2816978de565c0c02f176;
wire [MAX_SUM_WDTH_L-1:0]        I6f9a280cf50379308d67506d6d6a5c61;
wire [MAX_SUM_WDTH_L-1:0]        I77b54488bd26318f14b4364035cd1836;
wire [flogtanh_WDTH -1:0]        Ifb7004286169cd9b229b083aea58a408;
wire [MAX_SUM_WDTH_L-1:0]        Ia4e1d880c6b384bd3b315ab453e03326;
wire [MAX_SUM_WDTH_L-1:0]        I786338397f55073dce91e1c8c5f8e298;
wire [flogtanh_WDTH -1:0]        Ib04408fcc6f4d26fcdb5599b03b1b534;
wire [MAX_SUM_WDTH_L-1:0]        Icc8d6c731fe2502a4d041cc5aefcc9d8;
wire [MAX_SUM_WDTH_L-1:0]        I0e5931219d94c8e8e1f4af081404dcab;
wire [flogtanh_WDTH -1:0]        Ifda1a58a6f54318a30faa98dc1982e8e;
wire [MAX_SUM_WDTH_L-1:0]        I311ca38028cb07e4d7a8f3914aec47cc;
wire [MAX_SUM_WDTH_L-1:0]        I8d96b419b010f8076311420d7b9c8a18;
wire [flogtanh_WDTH -1:0]        I799ce64e6df49e2b62dc6beda4500146;
wire [MAX_SUM_WDTH_L-1:0]        I68dc05646fbd91403f254c5de1bc3c70;
wire [MAX_SUM_WDTH_L-1:0]        Ife13f962c7a8df3845cde104a959f678;
wire [flogtanh_WDTH -1:0]        Ia592b65aa89be2fcd981cf144683a298;
wire [MAX_SUM_WDTH_L-1:0]        I2550505d6e2fe478dd0c789bc3b823cf;
wire [MAX_SUM_WDTH_L-1:0]        I7f701ff37ad3fc34d2f4efafe5ff5351;
wire [flogtanh_WDTH -1:0]        Ib52365bf14aedf524bb23a4a6fe10551;
wire [MAX_SUM_WDTH_L-1:0]        Idc3ffe555b7641f987c8cc2cc2f7cb59;
wire [MAX_SUM_WDTH_L-1:0]        I43c815a8ce0b2df9744a525328969691;
wire [flogtanh_WDTH -1:0]        Ieba74e8bf3d692612c544af3ce6046fd;
wire [MAX_SUM_WDTH_L-1:0]        Ie9ab765b69fae4069793331ca0e0e5f7;
wire [MAX_SUM_WDTH_L-1:0]        I6c4a1ded9bf39091cf302ebe0103e2f0;
wire [flogtanh_WDTH -1:0]        I6cc1587e659f3f97d636485b708b1eeb;
wire [MAX_SUM_WDTH_L-1:0]        I371fef521a66e4761eb7b3e950d6ed5c;
wire [MAX_SUM_WDTH_L-1:0]        Icd4ff8d14af2699db2b5168027894ebb;
wire [flogtanh_WDTH -1:0]        I84b09aba55d2335f19faa5762aeedb89;
wire [MAX_SUM_WDTH_L-1:0]        I6dc9b65102f0ca4eccc76b6c0321beba;
wire [MAX_SUM_WDTH_L-1:0]        Ia79d52fe2130426c07890fcaa50137db;
wire [flogtanh_WDTH -1:0]        I3c4b9082ba72cade4d52924eff135135;
wire [MAX_SUM_WDTH_L-1:0]        If4ac2065f0165f0a22d459e53b74ba91;
wire [MAX_SUM_WDTH_L-1:0]        I308aaa8ac500b5589aa4af533a9062bf;
wire [flogtanh_WDTH -1:0]        I65f6c14ae4e7139fd858d7637ec3fd46;
wire [MAX_SUM_WDTH_L-1:0]        I9ee4045d22e1e23f26f255e747bc2c25;
wire [MAX_SUM_WDTH_L-1:0]        Iac91f4037e542d9fda30fadafe7e79ac;
wire [flogtanh_WDTH -1:0]        I02425810db970e5ef0b791dc4be103a9;
wire [MAX_SUM_WDTH_L-1:0]        Ia356c2d6982d65670b4c3b276950011a;
wire [MAX_SUM_WDTH_L-1:0]        I8cd5970682bc84881489c12ff073212c;
wire [flogtanh_WDTH -1:0]        Id0bc7b00dec58136a8016979d8a9faad;
wire [MAX_SUM_WDTH_L-1:0]        I711a3fd75980a579031be60aa25e1da4;
wire [MAX_SUM_WDTH_L-1:0]        I1ee27be7e1a38aff0039b21c45f406d1;
wire [flogtanh_WDTH -1:0]        I7c61892052c3c32343ed172d4ae354cc;
wire [MAX_SUM_WDTH_L-1:0]        I75a05a0c3ecaf5a582e01297b8dde431;
wire [MAX_SUM_WDTH_L-1:0]        Idf90f01353ad1057e11fd060442f4e53;
wire [flogtanh_WDTH -1:0]        I7cd312338aa5a86e1b05cc28ab7a2b23;
wire [MAX_SUM_WDTH_L-1:0]        Ib50109a1e4490b3bdaefc5bf87674df2;
wire [MAX_SUM_WDTH_L-1:0]        Id45f4e0f142b6c3925f24a37dcf7c0ae;
wire [flogtanh_WDTH -1:0]        I88d4372b4f7bfddd2af726c2df391287;
wire [MAX_SUM_WDTH_L-1:0]        I5717425e31d5707f3f1c7010cc261651;
wire [MAX_SUM_WDTH_L-1:0]        I52a9bcfbd2d3a763671f19cfeaf7bb8b;
wire [flogtanh_WDTH -1:0]        Ic8978ad86275ac6f4a0cf80ebefc5b27;
wire [MAX_SUM_WDTH_L-1:0]        Ie8244d4913aa3720080a883429b5f2e3;
wire [MAX_SUM_WDTH_L-1:0]        Ia3cc6acf2cae41e560e09993007ffd2b;
wire [flogtanh_WDTH -1:0]        I99745124c45f37d3882064590394a0aa;
wire [MAX_SUM_WDTH_L-1:0]        I32bcd4d63f2064e8b6058defcddf1523;
wire [MAX_SUM_WDTH_L-1:0]        Iba0d2f08788f2208a648ae7b5414195d;
wire [flogtanh_WDTH -1:0]        I33fe34f9be3c51b4b93f89c3f862e332;
wire [MAX_SUM_WDTH_L-1:0]        I3d765cb8f72daad8ad6fd19b230ef2e1;
wire [MAX_SUM_WDTH_L-1:0]        I9f7df6ad60284c812aeb522974578e0b;
wire [flogtanh_WDTH -1:0]        Iecda9a183e74f78b9fd5ce34e80d712e;
wire [MAX_SUM_WDTH_L-1:0]        I6c50eab3042fbe8d0a9c1f13b891ca3b;
wire [MAX_SUM_WDTH_L-1:0]        Iab1fb7006598181bd8749ed90c519b13;
wire [flogtanh_WDTH -1:0]        I5293b996bbf152abf110df1205ad4856;
wire [MAX_SUM_WDTH_L-1:0]        I7a87da6d33b578f6bc60ca0c4ee59cf5;
wire [MAX_SUM_WDTH_L-1:0]        Ieef3b299ec35075c71ef9fb10525bfc4;
wire [flogtanh_WDTH -1:0]        Ia99c08ee345bdc1489ce82a62481ef3b;
wire [MAX_SUM_WDTH_L-1:0]        I6ba6d7a611d9e209c8888454e1a9650e;
wire [MAX_SUM_WDTH_L-1:0]        I58a7c08adf48d0737c5803e2a818c045;
wire [flogtanh_WDTH -1:0]        Iaa314530e04145eb73672ebb150858af;
wire [MAX_SUM_WDTH_L-1:0]        I7b6878abc6b5d1bc713bb9128c238d9d;
wire [MAX_SUM_WDTH_L-1:0]        I30a1c8fcd9a510a6ed559f07dd809b90;
wire [flogtanh_WDTH -1:0]        I05f7363bfcc34691280079e82f6f5449;
wire [MAX_SUM_WDTH_L-1:0]        I3debbdfea21b3d4d975aff74df6a89a4;
wire [MAX_SUM_WDTH_L-1:0]        Ic4f5e9d49419e1c57cfa387761ab643d;
wire [flogtanh_WDTH -1:0]        Ica5ce135e77ed1d7cbc8277344ffeaeb;
wire [MAX_SUM_WDTH_L-1:0]        Ie21e2ff26b0c30eea53233d9142ec128;
wire [MAX_SUM_WDTH_L-1:0]        Id3dd71ea0bf0f2996fbe42b8c3318762;
wire [flogtanh_WDTH -1:0]        Iac98c702c4d9d78460fc7c212bce7841;
wire [MAX_SUM_WDTH_L-1:0]        I9134717dde036edd9737f695d9c791ae;
wire [MAX_SUM_WDTH_L-1:0]        Ib834b91bf81067e8efa9d470023e8b9d;
wire [flogtanh_WDTH -1:0]        I1fe269380ba03e78a8e41c17aa4bd757;
wire [MAX_SUM_WDTH_L-1:0]        Ic492036079044fd3af487ee7c84e68d0;
wire [MAX_SUM_WDTH_L-1:0]        Ic6ead78ed741442f17a15a157cd6ef9c;
wire [flogtanh_WDTH -1:0]        Ib19549130ee3307413b69c50042f7302;
wire [MAX_SUM_WDTH_L-1:0]        Ib6e42f1caafaddc1c964b5b04862f5c1;
wire [MAX_SUM_WDTH_L-1:0]        I4e257dbd6f196a02dc0f5a2e5f6047d7;
wire [flogtanh_WDTH -1:0]        Iad6acaf97d307fdbe0f20bf010acb468;
wire [MAX_SUM_WDTH_L-1:0]        I54e99c231380749e3d48384c78fbf0e8;
wire [MAX_SUM_WDTH_L-1:0]        I3dbfbd34d1fdfd4f422d900154123b6b;
wire [flogtanh_WDTH -1:0]        I67c9882f9e19df5a7b9bd0d900bb2f75;
wire [MAX_SUM_WDTH_L-1:0]        I4acf64c7b000236974dc1762d0d7223e;
wire [MAX_SUM_WDTH_L-1:0]        I529b763dace1924613d184c6c70c2708;
wire [flogtanh_WDTH -1:0]        I3099768bc986a11350656e472fc21ac1;
wire [MAX_SUM_WDTH_L-1:0]        Ib5f05c310200a5759e4dd169a9b3ca8c;
wire [MAX_SUM_WDTH_L-1:0]        I7a600aeb6cf8c3311c10afa4d82767a1;
wire [flogtanh_WDTH -1:0]        Ifba5972f9d38199dbc675432a29934e4;
wire [MAX_SUM_WDTH_L-1:0]        Ibeef99739eace0ce4d691cd2b4075571;
wire [MAX_SUM_WDTH_L-1:0]        I8c7aab31f8cb705ea13a41a5bd349303;
wire [flogtanh_WDTH -1:0]        I0934fb292b19451a050fb3374a7bd1a7;
wire [MAX_SUM_WDTH_L-1:0]        Iea5ee3bf75ed967ef2dfc8ed8d9bbc2f;
wire [MAX_SUM_WDTH_L-1:0]        I171149dcaab2c0f0e2a10547ad95084d;
wire [flogtanh_WDTH -1:0]        I9a3d1741c77fb1bbc1a54383874de82a;
wire [MAX_SUM_WDTH_L-1:0]        Ib10b3fb9882f1a07acee84ad15ad21f1;
wire [MAX_SUM_WDTH_L-1:0]        I23b60ca4da2df0ec40c1df62d058deef;
wire [flogtanh_WDTH -1:0]        If89f2ce813bab91af88f73ddc570d5a1;
wire [MAX_SUM_WDTH_L-1:0]        I7a74e6f3e2acbd05e92ff91cc8771f91;
wire [MAX_SUM_WDTH_L-1:0]        I7978d2d800b4438d0644ae3df6bcac9c;
wire [flogtanh_WDTH -1:0]        Ibc0dfcffac26f4898d42808534f6588f;
wire [MAX_SUM_WDTH_L-1:0]        I8f718fbf0d8b43af7002b67f6e0ef202;
wire [MAX_SUM_WDTH_L-1:0]        Ibc4eddc0f1768e9ec7e38e951a28ec42;
wire [flogtanh_WDTH -1:0]        I3a0a6f3d0141e8ad04d89c4bf306a96f;
wire [MAX_SUM_WDTH_L-1:0]        I3bf775756dc497fa91654eb7cf0657e9;
wire [MAX_SUM_WDTH_L-1:0]        I1c97fd1d21a31af8b5498a79b1a3e7b6;
wire [flogtanh_WDTH -1:0]        I1c875571dd1be1bb28aa15554964b485;
wire [MAX_SUM_WDTH_L-1:0]        I7c6d4cac0d6ff029d636fa006aa59912;
wire [MAX_SUM_WDTH_L-1:0]        Ie4f063eeaf7ee3f033e2a01ffaca623e;
wire [flogtanh_WDTH -1:0]        Ide5d5fdcf86b369b015890030a222a0a;
wire [MAX_SUM_WDTH_L-1:0]        I46249ffce3ba1abfbaaf1447070c1990;
wire [MAX_SUM_WDTH_L-1:0]        Ibb3d57d510cad00064a331f61f6400a2;
wire [flogtanh_WDTH -1:0]        I7cf6e8d40e7bd7685a7260638523690c;
wire [MAX_SUM_WDTH_L-1:0]        I13b24152d7160e4e4c0b8de8ca43ce6a;
wire [MAX_SUM_WDTH_L-1:0]        I9485ae915474a31562ce358666d66245;
wire [flogtanh_WDTH -1:0]        I52ccac771cc9a1c1797862bc781e1f58;
wire [MAX_SUM_WDTH_L-1:0]        If1d125c997fc331af17a03fa647c3a1e;
wire [MAX_SUM_WDTH_L-1:0]        Ia54b6f7044a831020e49f1bf48bc063a;
wire [flogtanh_WDTH -1:0]        I9db2090916f2535b14ed3292e78baa32;
wire [MAX_SUM_WDTH_L-1:0]        Id02c9cea3b4048f89cdb011325b5f874;
wire [MAX_SUM_WDTH_L-1:0]        Ie71c7babb5d17378d40444b6bbd4e7a6;
wire [flogtanh_WDTH -1:0]        I5b77a8ce7f495ae61315d1590bfd71b8;
wire [MAX_SUM_WDTH_L-1:0]        Iaabab9f3f0c05d0d5fba679bbcb14b3d;
wire [MAX_SUM_WDTH_L-1:0]        Ia0977b79857bdbf058535c30e338c38a;
wire [flogtanh_WDTH -1:0]        I4e4bb795cf09757c8ad3933c9ce4686f;
wire [MAX_SUM_WDTH_L-1:0]        I2bfaf258762bbc682298a56d3092d369;
wire [MAX_SUM_WDTH_L-1:0]        I600ea1371a2be66430ac9534583b512b;
wire [flogtanh_WDTH -1:0]        I78c29808e737dab48b5144b232dd02f6;
wire [MAX_SUM_WDTH_L-1:0]        If15b5be646c24f6e8ab29b0b7646ebe0;
wire [MAX_SUM_WDTH_L-1:0]        Ife5b9afdbb30c122b84d5378f9cb366d;
wire [flogtanh_WDTH -1:0]        Ie2ae83a457d79fbddc640d49d626171c;
wire [MAX_SUM_WDTH_L-1:0]        I58a4e50090f1a5028e267e31bf7c2e00;
wire [MAX_SUM_WDTH_L-1:0]        I27556d599dd1a27ee8f49e819ccbf29a;
wire [flogtanh_WDTH -1:0]        I3711e49a4eec517e47897fb731d75958;
wire [MAX_SUM_WDTH_L-1:0]        I2f87ae03574e521a6911a4dcd3dc4ec3;
wire [MAX_SUM_WDTH_L-1:0]        Icce595233ce089eafcca3eae5e71e5f8;
wire [flogtanh_WDTH -1:0]        Ifda4e727eb6275266f583badb6d4a9ed;
wire [MAX_SUM_WDTH_L-1:0]        I84e1a5675d75723d7c5fd8ec7a8bd093;
wire [MAX_SUM_WDTH_L-1:0]        Icc3cadf40c09be1a8c2847caf0e3e63c;
wire [flogtanh_WDTH -1:0]        I2be66a82c7b58e3c14b5816522b46969;
wire [MAX_SUM_WDTH_L-1:0]        I905aab3b31d9dd6fecb74ede9f4c56c0;
wire [MAX_SUM_WDTH_L-1:0]        Ib43886d923b8c683004713ff25b2f90d;
wire [flogtanh_WDTH -1:0]        I826fe7ad9e67061800d5d6543d779864;
wire [MAX_SUM_WDTH_L-1:0]        I66d3f7876f1fdc9a4d753a3bbd462300;
wire [MAX_SUM_WDTH_L-1:0]        I132d9671c582876568c0f7f5335f5227;
wire [flogtanh_WDTH -1:0]        Ic0c9069041758b53f56a46da81dd2d60;
wire [MAX_SUM_WDTH_L-1:0]        I3cd15e755f29b592bf2c1532e86d8f33;
wire [MAX_SUM_WDTH_L-1:0]        I0859c80b42a8c60dade8f05d58ee3701;
wire [flogtanh_WDTH -1:0]        I6f4c5a8de7690fec959861f43c134915;
wire [MAX_SUM_WDTH_L-1:0]        I14423aefbe6d66dbd2f518ae34f43f61;
wire [MAX_SUM_WDTH_L-1:0]        Ib3690ec149adde94343d3e617931a287;
wire [flogtanh_WDTH -1:0]        I14f1005a8c0fbdc5ca02c032b8891c2b;
wire [MAX_SUM_WDTH_L-1:0]        Ib1331d92ac9a84842b3e1b81968f241c;
wire [MAX_SUM_WDTH_L-1:0]        I41f2bf9ff00f983ad1298c8c83b041cb;
wire [flogtanh_WDTH -1:0]        Iacd30dfb96f6572ec56eff0a4094ec04;
wire [MAX_SUM_WDTH_L-1:0]        If5d175d3ad99e5f1a37ca02c5b72b550;
wire [MAX_SUM_WDTH_L-1:0]        Ib5414585cd6976cfce42e42190cc08d7;
wire [flogtanh_WDTH -1:0]        I1c748b8fe4979331bc3fe5aff4b6f9f4;
wire [MAX_SUM_WDTH_L-1:0]        I44e3174343cfa4f55b79f77e80005fbb;
wire [MAX_SUM_WDTH_L-1:0]        I1ca59325ff30db83df5bf0a2cd9706b6;
wire [flogtanh_WDTH -1:0]        I158c7973974f36c2793127964e50d1bd;
wire [MAX_SUM_WDTH_L-1:0]        I7d917703c26558414d5fb997398a8757;
wire [MAX_SUM_WDTH_L-1:0]        Ie2f5b03f3b136e651b8aba92a30d298a;
wire [flogtanh_WDTH -1:0]        Id5ea6ba2402275cb925a1848b31ec2e1;
wire [MAX_SUM_WDTH_L-1:0]        I5ff9bb8ef0620b2a968cc99b709723c7;
wire [MAX_SUM_WDTH_L-1:0]        I312ce79a8dd2ce3d37c930d42640509b;
wire [flogtanh_WDTH -1:0]        I3862f7017bc2bc69844b73f2a79f47f5;
wire [MAX_SUM_WDTH_L-1:0]        Icb83a6adcf84370776ad71a9f5a8735b;
wire [MAX_SUM_WDTH_L-1:0]        I467d5e2554ef25873e0b44e947ee0011;
wire [flogtanh_WDTH -1:0]        I4ed41fde5449b7112baf000a05484ac4;
wire [MAX_SUM_WDTH_L-1:0]        Ieaa23d9c0997f273064a57b8071c64c1;
wire [MAX_SUM_WDTH_L-1:0]        Ice73b514709469fd21cd254bf4ceadd9;
wire [flogtanh_WDTH -1:0]        I40c4db2872b602bf9d6a4fc4ba5ac34d;
wire [MAX_SUM_WDTH_L-1:0]        I69b89cf26b64d319f7796610e92caec9;
wire [MAX_SUM_WDTH_L-1:0]        I45ba06a6d6f00c174b1439a6f226a085;
wire [flogtanh_WDTH -1:0]        Ibe5ab52bd0f220f7a6aac244c0e3867e;
wire [MAX_SUM_WDTH_L-1:0]        I6bf4038fafaa59349f73aa011149067e;
wire [MAX_SUM_WDTH_L-1:0]        Ic8a272f82736fd599fb3250e970edf9b;
wire [flogtanh_WDTH -1:0]        I36668064f280c70f9143ee9f39973015;
wire [MAX_SUM_WDTH_L-1:0]        Idbe16e45feac2ab46cd58d32eb0e3113;
wire [MAX_SUM_WDTH_L-1:0]        I5b9710b16effc8bf0695517c6e651836;
wire [flogtanh_WDTH -1:0]        Ief92462253c5a03a42d46ed7087caf9a;
wire [MAX_SUM_WDTH_L-1:0]        I11eb91a1ff576ec2787ec76b0787977c;
wire [MAX_SUM_WDTH_L-1:0]        I038b42a83025f5eaebf45799d1ebe7b0;
wire [flogtanh_WDTH -1:0]        Idf196345491ff3290796ba7827d31c17;
wire [MAX_SUM_WDTH_L-1:0]        Ie45dede493b6ce54a123db34cfedcefe;
wire [MAX_SUM_WDTH_L-1:0]        I73ddd7cf9272ceab5a663e2244e72d7e;
wire [flogtanh_WDTH -1:0]        I2230f0e48899877bc2bcb3538be81bfa;
wire [MAX_SUM_WDTH_L-1:0]        I69df2773462a5c7a2802176217eeee01;
wire [MAX_SUM_WDTH_L-1:0]        I16507fab8f9076bfeb419896fa7cdc1d;
wire [flogtanh_WDTH -1:0]        Ibc0ec83d6b8e6be89ddc88ef83f0b03d;
wire [MAX_SUM_WDTH_L-1:0]        Id8a3ef0da815bdd206d02be6d7b82c89;
wire [MAX_SUM_WDTH_L-1:0]        I3dd1f28cf199299aba54e47a429c9b11;
wire [flogtanh_WDTH -1:0]        Ifc59c1b26ec09b3a7fe5a2b90511c93b;
wire [MAX_SUM_WDTH_L-1:0]        I9f74767b10d0981465160f7f9c915826;
wire [MAX_SUM_WDTH_L-1:0]        I49d9203dc6f8c17f17383e8f7e01f005;
wire [flogtanh_WDTH -1:0]        I9c6fc8e09cd63551f40accc98d784a44;
wire [MAX_SUM_WDTH_L-1:0]        I6340b82b10836e90efc17d3d8ce27aa4;
wire [MAX_SUM_WDTH_L-1:0]        Ibeec86c75d950ee00dd63a2930f08a24;
wire [flogtanh_WDTH -1:0]        I26692a6aab1d81d71219a436bee5e10b;
wire [MAX_SUM_WDTH_L-1:0]        Ief2d5177fa9a28016b5da2def9de4050;
wire [MAX_SUM_WDTH_L-1:0]        I47b2438c3680b2d816168df37d7c491c;
wire [flogtanh_WDTH -1:0]        Ieb50592e17305d0f74cbf216be947862;
wire [MAX_SUM_WDTH_L-1:0]        I49214ecffd1e025db688d04119248a84;
wire [MAX_SUM_WDTH_L-1:0]        I5983bf2c6c90b872ee6cf58b5e520311;
wire [flogtanh_WDTH -1:0]        I0071f023f1be4400541c13bc68278417;
wire [MAX_SUM_WDTH_L-1:0]        Icb84682ddc30efd01dcfe2d96a84ba9d;
wire [MAX_SUM_WDTH_L-1:0]        I6745cacecb7ee86cf3c7ad7eeee6048f;
wire [flogtanh_WDTH -1:0]        Ib2f1635b38ca6090e5ff633cbfa13273;
wire [MAX_SUM_WDTH_L-1:0]        I7f99c71ccc1918b7ee0ca2e9ed84ea17;
wire [MAX_SUM_WDTH_L-1:0]        Ib9672d20643d856ff31905ab14c0ac87;
wire [flogtanh_WDTH -1:0]        Id2c0bc90fd26e82fe91b5aef7bdd3a29;
wire [MAX_SUM_WDTH_L-1:0]        Ifbc9e59e2ea7b320ad2ec483bd58c1c4;
wire [MAX_SUM_WDTH_L-1:0]        Ib9dfea1f34a120eda30d5bd919365a6a;
wire [flogtanh_WDTH -1:0]        If4a723ce836f5327b85e234ebd195bd9;
wire [MAX_SUM_WDTH_L-1:0]        I98a7d5627114777569c3ad29fbdf33ce;
wire [MAX_SUM_WDTH_L-1:0]        Ia7bf82c9e5ca4467b5e50beeaeb975e9;
wire [flogtanh_WDTH -1:0]        If63dd5997e033817126a9ebaf38c1955;
wire [MAX_SUM_WDTH_L-1:0]        Ic3cf4882216f4f3c63524154ca5bf020;
wire [MAX_SUM_WDTH_L-1:0]        I327c9acb8934729b4ea5486787afa2e8;
wire [flogtanh_WDTH -1:0]        Ie2ee6baf8ec357f6131dff92fb480e42;
wire [MAX_SUM_WDTH_L-1:0]        Iaa2e0df90fb601ebaddcf0d4afaeedd2;
wire [MAX_SUM_WDTH_L-1:0]        Ieddef08050c38d07e5d38f5bb7b099c0;
wire [flogtanh_WDTH -1:0]        Ibff4d4fca3681fe10807414ed84e4157;
wire [MAX_SUM_WDTH_L-1:0]        I0f5bf0ab35c2588426d461588a882388;
wire [MAX_SUM_WDTH_L-1:0]        I39f9e8430db114991bfb27cc46ef3e39;
wire [flogtanh_WDTH -1:0]        I4540d74c919f50e9b6e40ef6b8cfd279;
wire [MAX_SUM_WDTH_L-1:0]        Ic7fc2a5137184b1908cb1293341fcf26;
wire [MAX_SUM_WDTH_L-1:0]        I56aa548618a4a15e9a35e04f5eeb823f;
wire [flogtanh_WDTH -1:0]        I01637ffca829d72accbb5dcee48817ca;
wire [MAX_SUM_WDTH_L-1:0]        I0e1b866232599fcb497ce38c2c68f32a;
wire [MAX_SUM_WDTH_L-1:0]        I1908897b529ca04df7e7da395be4a8ce;
wire [flogtanh_WDTH -1:0]        I7e8af960e934c7cc3cb163d6f8e7d597;
wire [MAX_SUM_WDTH_L-1:0]        Id526a3d6594056c40bd5c1ee1f109925;
wire [MAX_SUM_WDTH_L-1:0]        Ib2bbd59cd6098608ed53ac556036534f;
wire [flogtanh_WDTH -1:0]        Ifd80d371c8851b9e16193a3e62ddf79a;
wire [MAX_SUM_WDTH_L-1:0]        Ia75d451c04e28eb476104090e9f952b2;
wire [MAX_SUM_WDTH_L-1:0]        If004552b2047ab1cf23bb50375460b01;
wire [flogtanh_WDTH -1:0]        I19d2c4bc969133fa59d22f7f2d8cfd4a;
wire [MAX_SUM_WDTH_L-1:0]        Ib30ec3e9a870536690a38fe069018f42;
wire [MAX_SUM_WDTH_L-1:0]        If97092e1e2147de199c94a23831cf6b9;
wire [flogtanh_WDTH -1:0]        I532326ad245909d441134296dae9a5d4;
wire [MAX_SUM_WDTH_L-1:0]        I00edc092e1c7c9738943465938a693bd;
wire [MAX_SUM_WDTH_L-1:0]        Ibf74a4dfaab7f7f538d2b5fac7394b63;
wire [flogtanh_WDTH -1:0]        I6ca7199e28b480ac5816bf5b4cfb1eef;
wire [MAX_SUM_WDTH_L-1:0]        I4dc8aa3d45b1cbb2a926179a5cccdf57;
wire [MAX_SUM_WDTH_L-1:0]        I991a7a7d562eb0a8b4b8d8f008ef2225;
wire [flogtanh_WDTH -1:0]        I0d5b26d24fbce6b236120b5697d0db6b;
wire [MAX_SUM_WDTH_L-1:0]        I4a60dfcad5fab348684831c1c5301d02;
wire [MAX_SUM_WDTH_L-1:0]        I64c3d7be41abaa17d6992f9af8e72789;
wire [flogtanh_WDTH -1:0]        I618d329f2b0f18617d80aa350b79601c;
wire [MAX_SUM_WDTH_L-1:0]        I6d9fce52b1224fa10ee9bd3e5a02b68b;
wire [MAX_SUM_WDTH_L-1:0]        Icb91e63ebabc7a75a54eb7c731df4fa0;
wire [flogtanh_WDTH -1:0]        I58e3a5e842e14d09de91959839798a67;
wire [MAX_SUM_WDTH_L-1:0]        Ifcc8638ec8cc700bfafedd844eabe861;
wire [MAX_SUM_WDTH_L-1:0]        I673d1d0d0daab99bd940c46cc14ef55a;
wire [flogtanh_WDTH -1:0]        Icdecd5095ef818a0915ff3fcb395db5b;
wire [MAX_SUM_WDTH_L-1:0]        I60914917663174bf0a5f6b1b16a0a1ce;
wire [MAX_SUM_WDTH_L-1:0]        I62cadbd70b07a6a7a2974c7c392696b3;
wire [flogtanh_WDTH -1:0]        I236f843994d3065b6ee70c41f390a3d0;
wire [MAX_SUM_WDTH_L-1:0]        I4ef6d192effc3fb6d583b0370194cd62;
wire [MAX_SUM_WDTH_L-1:0]        Icd8257d7f53d93db989eb56eaeb7e593;
wire [flogtanh_WDTH -1:0]        I7a9001d6c1d1aa8af79d9b152e596b70;
wire [MAX_SUM_WDTH_L-1:0]        I9fe9281eeaac31b7c9499f5c3e8bfe9a;
wire [MAX_SUM_WDTH_L-1:0]        I05931ceae6eff26e5a66a44a54d628ae;
wire [flogtanh_WDTH -1:0]        I56a43a072d463792d9e676c4907b3e76;
wire [MAX_SUM_WDTH_L-1:0]        I80bc60c27d0ebfc778d59b578732f07e;
wire [MAX_SUM_WDTH_L-1:0]        I306fec0aa68a0396053a6e0fa1cda38f;
wire [flogtanh_WDTH -1:0]        I336a86e85d3a8a42c4b6458ccb92ae05;
wire [MAX_SUM_WDTH_L-1:0]        Id371abee85a8611bc9f15cb475c76169;
wire [MAX_SUM_WDTH_L-1:0]        Idee8c8144207d676d1f2f9064bbdff45;
wire [flogtanh_WDTH -1:0]        Id97f66b78f1e3b6bf0b962b85ca1cde7;
wire [MAX_SUM_WDTH_L-1:0]        Ida40585da3f7140c84ef2d0088d42977;
wire [MAX_SUM_WDTH_L-1:0]        I5855124d566af739caa6511f8598f2c5;
wire [flogtanh_WDTH -1:0]        I52c7f0a8f9b4533052b5acd1b5bd5e17;
wire [MAX_SUM_WDTH_L-1:0]        Ib175445b5c07a6fd6e4ea0dc6e6952fe;
wire [MAX_SUM_WDTH_L-1:0]        I50729db4a8e04f18979707df14cb2419;
wire [flogtanh_WDTH -1:0]        I3b1db672b1a94502b90451260062a274;
wire [MAX_SUM_WDTH_L-1:0]        Idb001650555c8e77733c2cae7b6f099f;
wire [MAX_SUM_WDTH_L-1:0]        Ia3cb3ea64576a3e7332e1fb55953aa3e;
wire [flogtanh_WDTH -1:0]        I1a83f91eb1262911ae8d99e305294bf8;
wire [MAX_SUM_WDTH_L-1:0]        Icfa6a05bc48790590b66ff78773cc9a6;
wire [MAX_SUM_WDTH_L-1:0]        I3cb1f233951d49f985b0deac6e052bfd;
wire [flogtanh_WDTH -1:0]        Id01bfbd86b6321a843e239ca97cec514;
wire [MAX_SUM_WDTH_L-1:0]        Ib953adc95f33e5f0f97545b7ac0e6a82;
wire [MAX_SUM_WDTH_L-1:0]        I7015def91103398e54f446ce3e43af01;
wire [flogtanh_WDTH -1:0]        I26b769b58e1c21b68dd95c9f38c0362b;
wire [MAX_SUM_WDTH_L-1:0]        I3e379d83cf4dae9968eaadd4da9e2b4c;
wire [MAX_SUM_WDTH_L-1:0]        I04874bd1bf257f205b5189c8c20e5a12;
wire [flogtanh_WDTH -1:0]        Ic86f9988281398adfe43152beb722c1b;
wire [MAX_SUM_WDTH_L-1:0]        I51508292b5316d23e45d217d48eb623d;
wire [MAX_SUM_WDTH_L-1:0]        I937e3a8ede2305ea7c1750283224a870;
wire [flogtanh_WDTH -1:0]        I9d8ac6c29c2f5df7c2d124dface59e35;
wire [MAX_SUM_WDTH_L-1:0]        I36d727f90d4a830f79443b4941c9df9c;
wire [MAX_SUM_WDTH_L-1:0]        Ia7206430a739a11af4d860096eedd6c3;
wire [flogtanh_WDTH -1:0]        I56b46c426895409b40c3be9b79365a8a;
wire [MAX_SUM_WDTH_L-1:0]        I519b932add092db1a149df22a471d04e;
wire [MAX_SUM_WDTH_L-1:0]        Ibf4c2c00f8e012e9498361bfd3c5b06e;
wire [flogtanh_WDTH -1:0]        Ic63de8464f79ae05f27f05c935dbf495;
wire [MAX_SUM_WDTH_L-1:0]        I44395e9b406cd0ae7b3672e8ff86af4d;
wire [MAX_SUM_WDTH_L-1:0]        I899e5f03cd1d52d11f898959559aaeea;
wire [flogtanh_WDTH -1:0]        I4d21ee443e5921532d5bf1db7ef93f82;
wire [MAX_SUM_WDTH_L-1:0]        I08955fcfabffed0ad0c5e398e7872be1;
wire [MAX_SUM_WDTH_L-1:0]        I59c80c7ec26f43308b1a646c47160568;
wire [flogtanh_WDTH -1:0]        Ieb5fa20abbdb29a7f75021b7afafea31;
wire [MAX_SUM_WDTH_L-1:0]        I99252b9918c30f2ba5611abc79e08fbb;
wire [MAX_SUM_WDTH_L-1:0]        I8a954a331d36266465a0813d2e8b319b;
wire [flogtanh_WDTH -1:0]        I16a12326344aadf4226bd149424a53a8;
wire [MAX_SUM_WDTH_L-1:0]        I9cb632c1ab546359ef5a787a4bc3aaa6;
wire [MAX_SUM_WDTH_L-1:0]        Ib49e53ca8efd9564ee9572eb3089bb51;
wire [flogtanh_WDTH -1:0]        I07f36b533b48344c13dbb133739712f4;
wire [MAX_SUM_WDTH_L-1:0]        Ia4ee264b162c3ab4fec78ddb3a4fc6da;
wire [MAX_SUM_WDTH_L-1:0]        Icbde2c6230e9cc67ef12031e38bb344f;
wire [flogtanh_WDTH -1:0]        I7a0072bf1e5fb0c4de85c6e4447878a4;
wire [MAX_SUM_WDTH_L-1:0]        I116d3b804a2077edec9cf686b7cf5737;
wire [MAX_SUM_WDTH_L-1:0]        I2e22e867f6f84a7807b82f64a147022e;
wire [flogtanh_WDTH -1:0]        I320bafc5a1775d6933bcb9f2d2c84576;
wire [MAX_SUM_WDTH_L-1:0]        I5f89382f736f2688bc2c3696e0796002;
wire [MAX_SUM_WDTH_L-1:0]        Id9704e1d8096cd28577c5c357d30b7a4;
wire [flogtanh_WDTH -1:0]        I5ec61756ff7237146f2d83f17eb5bb3a;
wire [MAX_SUM_WDTH_L-1:0]        Ie139e712a1c886d4452735c1cd51af2e;
wire [MAX_SUM_WDTH_L-1:0]        I4b8554cab486a4fc1e14884a6495016e;
wire [flogtanh_WDTH -1:0]        I382008a17338641e68fa859ac2af1d20;
wire [MAX_SUM_WDTH_L-1:0]        Ic3137e053b8e22028a8ccdeb9c573170;
wire [MAX_SUM_WDTH_L-1:0]        Iaa235d085a5916a3b0814c3ed2a9026f;
wire [flogtanh_WDTH -1:0]        Ifd375ad8038ea2455c0e3b1463b83b7e;
wire [MAX_SUM_WDTH_L-1:0]        I8e15864be74893cd89bc56c0c2df858a;
wire [MAX_SUM_WDTH_L-1:0]        I5d86ce0b58c0b281d747116a9069ef33;
wire [flogtanh_WDTH -1:0]        I0b75763235278d8eca6ca72fc97fb83c;
wire [MAX_SUM_WDTH_L-1:0]        I015b6b916b0b84ddbfded84bca8f849f;
wire [MAX_SUM_WDTH_L-1:0]        Id20394136fb036435bb4680aac64581f;
wire [flogtanh_WDTH -1:0]        I9bc4c3b77a9635bb77ad31527d961952;
wire [MAX_SUM_WDTH_L-1:0]        I7ee0d250f9a3166db6bd3f366059804a;
wire [MAX_SUM_WDTH_L-1:0]        I8a16afac6e470ca69634d7fe9656387a;
wire [flogtanh_WDTH -1:0]        Ief93f4a7eaaa1f43ea1788dc4629c093;
wire [MAX_SUM_WDTH_L-1:0]        I6fc4b3ab1858416a94ce844cd92277ce;
wire [MAX_SUM_WDTH_L-1:0]        Ic4e7f690bc050f1d1f84eae7ca193e1c;
wire [flogtanh_WDTH -1:0]        I34b86fbc3949cb2083931ad8edd2444d;
wire [MAX_SUM_WDTH_L-1:0]        I9035dc3d53fc938d0927370681b669b3;
wire [MAX_SUM_WDTH_L-1:0]        Ia60421aa427236540b4d0d08d52ff507;
wire [flogtanh_WDTH -1:0]        I560c163fb55aa4b56da25f96e9b8ef6c;
wire [MAX_SUM_WDTH_L-1:0]        I162c001a328c8bbc178403bc97725ed6;
wire [MAX_SUM_WDTH_L-1:0]        Icace650ee3865bd7bbddd2d9435c5561;
wire [flogtanh_WDTH -1:0]        Ib3c46d34c5bc3d2651147b3e764d9786;
wire [MAX_SUM_WDTH_L-1:0]        I5fac1be3058558fcba4ae7c095138a07;
wire [MAX_SUM_WDTH_L-1:0]        I7d27d070b96b7810f667e1d1845342d3;
wire [flogtanh_WDTH -1:0]        Ie5e2ba4fe22870afc81d6cfc708570be;
wire [MAX_SUM_WDTH_L-1:0]        I0e7ff238062811c5a3d3549bbf3bec52;
wire [MAX_SUM_WDTH_L-1:0]        Ida7ec09c913caa0e78a2c4cbaae517c8;
wire [flogtanh_WDTH -1:0]        Ibf3bde181da4f960537516d6c0b2a72c;
wire [MAX_SUM_WDTH_L-1:0]        Ie6509743f0bbe16d5f0aae9039db3d21;
wire [MAX_SUM_WDTH_L-1:0]        Ic5eba898858be1f768841ead792d6d86;
wire [flogtanh_WDTH -1:0]        Ia93f96aa0718f8755e9ebb8cc5d8f405;
wire [MAX_SUM_WDTH_L-1:0]        I2b807f3aaa37eaddf34d61f95d436d48;
wire [MAX_SUM_WDTH_L-1:0]        I72197797a307c611fa8952533e63d7bf;

reg                              start_d2;
reg                              start_d3;
reg                              start_d4;
reg                              start_d5;
reg                              start_d6;
reg                              start_d7;
reg                              start_d8;
reg                              start_d9;


wire [fgallag_WDTH-1:0]          fgallag_00000_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00000_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00000_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00000_00000;
wire [fgallag_WDTH-1:0]          fgallag_00000_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00000_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00000_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00000_00001;
wire [fgallag_WDTH-1:0]          fgallag_00000_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00000_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00000_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00000_00002;
wire [fgallag_WDTH-1:0]          fgallag_00000_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00000_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00000_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00000_00003;
wire [fgallag_WDTH-1:0]          fgallag_00000_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00000_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00000_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00000_00004;
wire [fgallag_WDTH-1:0]          fgallag_00000_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00000_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00000_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00000_00005;
wire [fgallag_WDTH-1:0]          fgallag_00000_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00000_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00000_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00000_00006;
wire [fgallag_WDTH-1:0]          fgallag_00000_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00000_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00000_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00000_00007;
wire [fgallag_WDTH-1:0]          fgallag_00001_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00001_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00001_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00001_00000;
wire [fgallag_WDTH-1:0]          fgallag_00001_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00001_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00001_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00001_00001;
wire [fgallag_WDTH-1:0]          fgallag_00001_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00001_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00001_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00001_00002;
wire [fgallag_WDTH-1:0]          fgallag_00001_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00001_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00001_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00001_00003;
wire [fgallag_WDTH-1:0]          fgallag_00001_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00001_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00001_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00001_00004;
wire [fgallag_WDTH-1:0]          fgallag_00001_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00001_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00001_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00001_00005;
wire [fgallag_WDTH-1:0]          fgallag_00001_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00001_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00001_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00001_00006;
wire [fgallag_WDTH-1:0]          fgallag_00001_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00001_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00001_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00001_00007;
wire [fgallag_WDTH-1:0]          fgallag_00002_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00002_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00002_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00002_00000;
wire [fgallag_WDTH-1:0]          fgallag_00002_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00002_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00002_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00002_00001;
wire [fgallag_WDTH-1:0]          fgallag_00002_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00002_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00002_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00002_00002;
wire [fgallag_WDTH-1:0]          fgallag_00002_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00002_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00002_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00002_00003;
wire [fgallag_WDTH-1:0]          fgallag_00002_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00002_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00002_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00002_00004;
wire [fgallag_WDTH-1:0]          fgallag_00002_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00002_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00002_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00002_00005;
wire [fgallag_WDTH-1:0]          fgallag_00002_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00002_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00002_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00002_00006;
wire [fgallag_WDTH-1:0]          fgallag_00002_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00002_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00002_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00002_00007;
wire [fgallag_WDTH-1:0]          fgallag_00003_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00003_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00003_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00003_00000;
wire [fgallag_WDTH-1:0]          fgallag_00003_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00003_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00003_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00003_00001;
wire [fgallag_WDTH-1:0]          fgallag_00003_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00003_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00003_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00003_00002;
wire [fgallag_WDTH-1:0]          fgallag_00003_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00003_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00003_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00003_00003;
wire [fgallag_WDTH-1:0]          fgallag_00003_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00003_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00003_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00003_00004;
wire [fgallag_WDTH-1:0]          fgallag_00003_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00003_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00003_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00003_00005;
wire [fgallag_WDTH-1:0]          fgallag_00003_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00003_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00003_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00003_00006;
wire [fgallag_WDTH-1:0]          fgallag_00003_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00003_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00003_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00003_00007;
wire [fgallag_WDTH-1:0]          fgallag_00004_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00004_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00004_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00004_00000;
wire [fgallag_WDTH-1:0]          fgallag_00004_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00004_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00004_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00004_00001;
wire [fgallag_WDTH-1:0]          fgallag_00004_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00004_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00004_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00004_00002;
wire [fgallag_WDTH-1:0]          fgallag_00004_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00004_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00004_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00004_00003;
wire [fgallag_WDTH-1:0]          fgallag_00004_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00004_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00004_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00004_00004;
wire [fgallag_WDTH-1:0]          fgallag_00004_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00004_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00004_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00004_00005;
wire [fgallag_WDTH-1:0]          fgallag_00004_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00004_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00004_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00004_00006;
wire [fgallag_WDTH-1:0]          fgallag_00004_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00004_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00004_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00004_00007;
wire [fgallag_WDTH-1:0]          fgallag_00004_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00004_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00004_00008;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00004_00008;
wire [fgallag_WDTH-1:0]          fgallag_00004_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00004_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00004_00009;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00004_00009;
wire [fgallag_WDTH-1:0]          fgallag_00005_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00005_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00005_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00005_00000;
wire [fgallag_WDTH-1:0]          fgallag_00005_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00005_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00005_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00005_00001;
wire [fgallag_WDTH-1:0]          fgallag_00005_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00005_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00005_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00005_00002;
wire [fgallag_WDTH-1:0]          fgallag_00005_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00005_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00005_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00005_00003;
wire [fgallag_WDTH-1:0]          fgallag_00005_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00005_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00005_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00005_00004;
wire [fgallag_WDTH-1:0]          fgallag_00005_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00005_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00005_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00005_00005;
wire [fgallag_WDTH-1:0]          fgallag_00005_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00005_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00005_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00005_00006;
wire [fgallag_WDTH-1:0]          fgallag_00005_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00005_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00005_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00005_00007;
wire [fgallag_WDTH-1:0]          fgallag_00005_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00005_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00005_00008;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00005_00008;
wire [fgallag_WDTH-1:0]          fgallag_00005_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00005_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00005_00009;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00005_00009;
wire [fgallag_WDTH-1:0]          fgallag_00006_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00006_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00006_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00006_00000;
wire [fgallag_WDTH-1:0]          fgallag_00006_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00006_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00006_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00006_00001;
wire [fgallag_WDTH-1:0]          fgallag_00006_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00006_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00006_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00006_00002;
wire [fgallag_WDTH-1:0]          fgallag_00006_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00006_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00006_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00006_00003;
wire [fgallag_WDTH-1:0]          fgallag_00006_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00006_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00006_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00006_00004;
wire [fgallag_WDTH-1:0]          fgallag_00006_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00006_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00006_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00006_00005;
wire [fgallag_WDTH-1:0]          fgallag_00006_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00006_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00006_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00006_00006;
wire [fgallag_WDTH-1:0]          fgallag_00006_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00006_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00006_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00006_00007;
wire [fgallag_WDTH-1:0]          fgallag_00006_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00006_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00006_00008;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00006_00008;
wire [fgallag_WDTH-1:0]          fgallag_00006_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00006_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00006_00009;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00006_00009;
wire [fgallag_WDTH-1:0]          fgallag_00007_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00007_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00007_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00007_00000;
wire [fgallag_WDTH-1:0]          fgallag_00007_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00007_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00007_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00007_00001;
wire [fgallag_WDTH-1:0]          fgallag_00007_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00007_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00007_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00007_00002;
wire [fgallag_WDTH-1:0]          fgallag_00007_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00007_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00007_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00007_00003;
wire [fgallag_WDTH-1:0]          fgallag_00007_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00007_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00007_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00007_00004;
wire [fgallag_WDTH-1:0]          fgallag_00007_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00007_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00007_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00007_00005;
wire [fgallag_WDTH-1:0]          fgallag_00007_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00007_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00007_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00007_00006;
wire [fgallag_WDTH-1:0]          fgallag_00007_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00007_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00007_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00007_00007;
wire [fgallag_WDTH-1:0]          fgallag_00007_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00007_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00007_00008;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00007_00008;
wire [fgallag_WDTH-1:0]          fgallag_00007_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00007_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00007_00009;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00007_00009;
wire [fgallag_WDTH-1:0]          fgallag_00008_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00008_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00008_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00008_00000;
wire [fgallag_WDTH-1:0]          fgallag_00008_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00008_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00008_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00008_00001;
wire [fgallag_WDTH-1:0]          fgallag_00008_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00008_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00008_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00008_00002;
wire [fgallag_WDTH-1:0]          fgallag_00008_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00008_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00008_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00008_00003;
wire [fgallag_WDTH-1:0]          fgallag_00008_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00008_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00008_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00008_00004;
wire [fgallag_WDTH-1:0]          fgallag_00008_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00008_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00008_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00008_00005;
wire [fgallag_WDTH-1:0]          fgallag_00008_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00008_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00008_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00008_00006;
wire [fgallag_WDTH-1:0]          fgallag_00008_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00008_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00008_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00008_00007;
wire [fgallag_WDTH-1:0]          fgallag_00009_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00009_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00009_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00009_00000;
wire [fgallag_WDTH-1:0]          fgallag_00009_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00009_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00009_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00009_00001;
wire [fgallag_WDTH-1:0]          fgallag_00009_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00009_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00009_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00009_00002;
wire [fgallag_WDTH-1:0]          fgallag_00009_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00009_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00009_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00009_00003;
wire [fgallag_WDTH-1:0]          fgallag_00009_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00009_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00009_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00009_00004;
wire [fgallag_WDTH-1:0]          fgallag_00009_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00009_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00009_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00009_00005;
wire [fgallag_WDTH-1:0]          fgallag_00009_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00009_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00009_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00009_00006;
wire [fgallag_WDTH-1:0]          fgallag_00009_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00009_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00009_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00009_00007;
wire [fgallag_WDTH-1:0]          fgallag_00010_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00010_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00010_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00010_00000;
wire [fgallag_WDTH-1:0]          fgallag_00010_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00010_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00010_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00010_00001;
wire [fgallag_WDTH-1:0]          fgallag_00010_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00010_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00010_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00010_00002;
wire [fgallag_WDTH-1:0]          fgallag_00010_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00010_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00010_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00010_00003;
wire [fgallag_WDTH-1:0]          fgallag_00010_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00010_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00010_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00010_00004;
wire [fgallag_WDTH-1:0]          fgallag_00010_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00010_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00010_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00010_00005;
wire [fgallag_WDTH-1:0]          fgallag_00010_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00010_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00010_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00010_00006;
wire [fgallag_WDTH-1:0]          fgallag_00010_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00010_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00010_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00010_00007;
wire [fgallag_WDTH-1:0]          fgallag_00011_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00011_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00011_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00011_00000;
wire [fgallag_WDTH-1:0]          fgallag_00011_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00011_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00011_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00011_00001;
wire [fgallag_WDTH-1:0]          fgallag_00011_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00011_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00011_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00011_00002;
wire [fgallag_WDTH-1:0]          fgallag_00011_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00011_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00011_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00011_00003;
wire [fgallag_WDTH-1:0]          fgallag_00011_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00011_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00011_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00011_00004;
wire [fgallag_WDTH-1:0]          fgallag_00011_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00011_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00011_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00011_00005;
wire [fgallag_WDTH-1:0]          fgallag_00011_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00011_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00011_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00011_00006;
wire [fgallag_WDTH-1:0]          fgallag_00011_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00011_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00011_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00011_00007;
wire [fgallag_WDTH-1:0]          fgallag_00012_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00012_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00012_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00012_00000;
wire [fgallag_WDTH-1:0]          fgallag_00012_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00012_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00012_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00012_00001;
wire [fgallag_WDTH-1:0]          fgallag_00012_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00012_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00012_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00012_00002;
wire [fgallag_WDTH-1:0]          fgallag_00012_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00012_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00012_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00012_00003;
wire [fgallag_WDTH-1:0]          fgallag_00012_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00012_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00012_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00012_00004;
wire [fgallag_WDTH-1:0]          fgallag_00012_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00012_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00012_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00012_00005;
wire [fgallag_WDTH-1:0]          fgallag_00012_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00012_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00012_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00012_00006;
wire [fgallag_WDTH-1:0]          fgallag_00012_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00012_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00012_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00012_00007;
wire [fgallag_WDTH-1:0]          fgallag_00012_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00012_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00012_00008;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00012_00008;
wire [fgallag_WDTH-1:0]          fgallag_00012_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00012_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00012_00009;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00012_00009;
wire [fgallag_WDTH-1:0]          fgallag_00013_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00013_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00013_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00013_00000;
wire [fgallag_WDTH-1:0]          fgallag_00013_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00013_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00013_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00013_00001;
wire [fgallag_WDTH-1:0]          fgallag_00013_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00013_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00013_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00013_00002;
wire [fgallag_WDTH-1:0]          fgallag_00013_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00013_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00013_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00013_00003;
wire [fgallag_WDTH-1:0]          fgallag_00013_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00013_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00013_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00013_00004;
wire [fgallag_WDTH-1:0]          fgallag_00013_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00013_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00013_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00013_00005;
wire [fgallag_WDTH-1:0]          fgallag_00013_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00013_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00013_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00013_00006;
wire [fgallag_WDTH-1:0]          fgallag_00013_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00013_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00013_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00013_00007;
wire [fgallag_WDTH-1:0]          fgallag_00013_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00013_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00013_00008;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00013_00008;
wire [fgallag_WDTH-1:0]          fgallag_00013_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00013_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00013_00009;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00013_00009;
wire [fgallag_WDTH-1:0]          fgallag_00014_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00014_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00014_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00014_00000;
wire [fgallag_WDTH-1:0]          fgallag_00014_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00014_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00014_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00014_00001;
wire [fgallag_WDTH-1:0]          fgallag_00014_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00014_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00014_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00014_00002;
wire [fgallag_WDTH-1:0]          fgallag_00014_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00014_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00014_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00014_00003;
wire [fgallag_WDTH-1:0]          fgallag_00014_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00014_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00014_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00014_00004;
wire [fgallag_WDTH-1:0]          fgallag_00014_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00014_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00014_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00014_00005;
wire [fgallag_WDTH-1:0]          fgallag_00014_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00014_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00014_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00014_00006;
wire [fgallag_WDTH-1:0]          fgallag_00014_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00014_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00014_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00014_00007;
wire [fgallag_WDTH-1:0]          fgallag_00014_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00014_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00014_00008;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00014_00008;
wire [fgallag_WDTH-1:0]          fgallag_00014_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00014_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00014_00009;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00014_00009;
wire [fgallag_WDTH-1:0]          fgallag_00015_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00015_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00015_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00015_00000;
wire [fgallag_WDTH-1:0]          fgallag_00015_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00015_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00015_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00015_00001;
wire [fgallag_WDTH-1:0]          fgallag_00015_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00015_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00015_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00015_00002;
wire [fgallag_WDTH-1:0]          fgallag_00015_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00015_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00015_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00015_00003;
wire [fgallag_WDTH-1:0]          fgallag_00015_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00015_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00015_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00015_00004;
wire [fgallag_WDTH-1:0]          fgallag_00015_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00015_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00015_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00015_00005;
wire [fgallag_WDTH-1:0]          fgallag_00015_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00015_00006;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00015_00006;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00015_00006;
wire [fgallag_WDTH-1:0]          fgallag_00015_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00015_00007;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00015_00007;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00015_00007;
wire [fgallag_WDTH-1:0]          fgallag_00015_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00015_00008;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00015_00008;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00015_00008;
wire [fgallag_WDTH-1:0]          fgallag_00015_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00015_00009;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00015_00009;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00015_00009;
wire [fgallag_WDTH-1:0]          fgallag_00016_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00016_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00016_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00016_00000;
wire [fgallag_WDTH-1:0]          fgallag_00016_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00016_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00016_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00016_00001;
wire [fgallag_WDTH-1:0]          fgallag_00016_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00016_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00016_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00016_00002;
wire [fgallag_WDTH-1:0]          fgallag_00016_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00016_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00016_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00016_00003;
wire [fgallag_WDTH-1:0]          fgallag_00017_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00017_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00017_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00017_00000;
wire [fgallag_WDTH-1:0]          fgallag_00017_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00017_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00017_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00017_00001;
wire [fgallag_WDTH-1:0]          fgallag_00017_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00017_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00017_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00017_00002;
wire [fgallag_WDTH-1:0]          fgallag_00017_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00017_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00017_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00017_00003;
wire [fgallag_WDTH-1:0]          fgallag_00018_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00018_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00018_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00018_00000;
wire [fgallag_WDTH-1:0]          fgallag_00018_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00018_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00018_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00018_00001;
wire [fgallag_WDTH-1:0]          fgallag_00018_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00018_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00018_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00018_00002;
wire [fgallag_WDTH-1:0]          fgallag_00018_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00018_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00018_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00018_00003;
wire [fgallag_WDTH-1:0]          fgallag_00019_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00019_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00019_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00019_00000;
wire [fgallag_WDTH-1:0]          fgallag_00019_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00019_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00019_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00019_00001;
wire [fgallag_WDTH-1:0]          fgallag_00019_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00019_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00019_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00019_00002;
wire [fgallag_WDTH-1:0]          fgallag_00019_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00019_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00019_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00019_00003;
wire [fgallag_WDTH-1:0]          fgallag_00020_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00020_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00020_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00020_00000;
wire [fgallag_WDTH-1:0]          fgallag_00020_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00020_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00020_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00020_00001;
wire [fgallag_WDTH-1:0]          fgallag_00020_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00020_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00020_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00020_00002;
wire [fgallag_WDTH-1:0]          fgallag_00020_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00020_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00020_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00020_00003;
wire [fgallag_WDTH-1:0]          fgallag_00020_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00020_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00020_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00020_00004;
wire [fgallag_WDTH-1:0]          fgallag_00020_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00020_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00020_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00020_00005;
wire [fgallag_WDTH-1:0]          fgallag_00021_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00021_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00021_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00021_00000;
wire [fgallag_WDTH-1:0]          fgallag_00021_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00021_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00021_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00021_00001;
wire [fgallag_WDTH-1:0]          fgallag_00021_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00021_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00021_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00021_00002;
wire [fgallag_WDTH-1:0]          fgallag_00021_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00021_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00021_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00021_00003;
wire [fgallag_WDTH-1:0]          fgallag_00021_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00021_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00021_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00021_00004;
wire [fgallag_WDTH-1:0]          fgallag_00021_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00021_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00021_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00021_00005;
wire [fgallag_WDTH-1:0]          fgallag_00022_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00022_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00022_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00022_00000;
wire [fgallag_WDTH-1:0]          fgallag_00022_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00022_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00022_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00022_00001;
wire [fgallag_WDTH-1:0]          fgallag_00022_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00022_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00022_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00022_00002;
wire [fgallag_WDTH-1:0]          fgallag_00022_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00022_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00022_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00022_00003;
wire [fgallag_WDTH-1:0]          fgallag_00022_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00022_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00022_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00022_00004;
wire [fgallag_WDTH-1:0]          fgallag_00022_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00022_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00022_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00022_00005;
wire [fgallag_WDTH-1:0]          fgallag_00023_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00023_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00023_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00023_00000;
wire [fgallag_WDTH-1:0]          fgallag_00023_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00023_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00023_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00023_00001;
wire [fgallag_WDTH-1:0]          fgallag_00023_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00023_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00023_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00023_00002;
wire [fgallag_WDTH-1:0]          fgallag_00023_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00023_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00023_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00023_00003;
wire [fgallag_WDTH-1:0]          fgallag_00023_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00023_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00023_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00023_00004;
wire [fgallag_WDTH-1:0]          fgallag_00023_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00023_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00023_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00023_00005;
wire [fgallag_WDTH-1:0]          fgallag_00024_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00024_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00024_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00024_00000;
wire [fgallag_WDTH-1:0]          fgallag_00024_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00024_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00024_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00024_00001;
wire [fgallag_WDTH-1:0]          fgallag_00024_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00024_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00024_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00024_00002;
wire [fgallag_WDTH-1:0]          fgallag_00024_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00024_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00024_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00024_00003;
wire [fgallag_WDTH-1:0]          fgallag_00024_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00024_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00024_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00024_00004;
wire [fgallag_WDTH-1:0]          fgallag_00024_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00024_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00024_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00024_00005;
wire [fgallag_WDTH-1:0]          fgallag_00025_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00025_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00025_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00025_00000;
wire [fgallag_WDTH-1:0]          fgallag_00025_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00025_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00025_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00025_00001;
wire [fgallag_WDTH-1:0]          fgallag_00025_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00025_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00025_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00025_00002;
wire [fgallag_WDTH-1:0]          fgallag_00025_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00025_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00025_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00025_00003;
wire [fgallag_WDTH-1:0]          fgallag_00025_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00025_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00025_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00025_00004;
wire [fgallag_WDTH-1:0]          fgallag_00025_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00025_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00025_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00025_00005;
wire [fgallag_WDTH-1:0]          fgallag_00026_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00026_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00026_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00026_00000;
wire [fgallag_WDTH-1:0]          fgallag_00026_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00026_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00026_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00026_00001;
wire [fgallag_WDTH-1:0]          fgallag_00026_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00026_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00026_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00026_00002;
wire [fgallag_WDTH-1:0]          fgallag_00026_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00026_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00026_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00026_00003;
wire [fgallag_WDTH-1:0]          fgallag_00026_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00026_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00026_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00026_00004;
wire [fgallag_WDTH-1:0]          fgallag_00026_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00026_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00026_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00026_00005;
wire [fgallag_WDTH-1:0]          fgallag_00027_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00027_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00027_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00027_00000;
wire [fgallag_WDTH-1:0]          fgallag_00027_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00027_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00027_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00027_00001;
wire [fgallag_WDTH-1:0]          fgallag_00027_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00027_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00027_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00027_00002;
wire [fgallag_WDTH-1:0]          fgallag_00027_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00027_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00027_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00027_00003;
wire [fgallag_WDTH-1:0]          fgallag_00027_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00027_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00027_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00027_00004;
wire [fgallag_WDTH-1:0]          fgallag_00027_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00027_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00027_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00027_00005;
wire [fgallag_WDTH-1:0]          fgallag_00028_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00028_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00028_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00028_00000;
wire [fgallag_WDTH-1:0]          fgallag_00028_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00028_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00028_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00028_00001;
wire [fgallag_WDTH-1:0]          fgallag_00028_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00028_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00028_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00028_00002;
wire [fgallag_WDTH-1:0]          fgallag_00028_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00028_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00028_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00028_00003;
wire [fgallag_WDTH-1:0]          fgallag_00028_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00028_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00028_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00028_00004;
wire [fgallag_WDTH-1:0]          fgallag_00028_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00028_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00028_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00028_00005;
wire [fgallag_WDTH-1:0]          fgallag_00029_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00029_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00029_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00029_00000;
wire [fgallag_WDTH-1:0]          fgallag_00029_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00029_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00029_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00029_00001;
wire [fgallag_WDTH-1:0]          fgallag_00029_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00029_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00029_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00029_00002;
wire [fgallag_WDTH-1:0]          fgallag_00029_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00029_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00029_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00029_00003;
wire [fgallag_WDTH-1:0]          fgallag_00029_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00029_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00029_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00029_00004;
wire [fgallag_WDTH-1:0]          fgallag_00029_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00029_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00029_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00029_00005;
wire [fgallag_WDTH-1:0]          fgallag_00030_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00030_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00030_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00030_00000;
wire [fgallag_WDTH-1:0]          fgallag_00030_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00030_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00030_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00030_00001;
wire [fgallag_WDTH-1:0]          fgallag_00030_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00030_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00030_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00030_00002;
wire [fgallag_WDTH-1:0]          fgallag_00030_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00030_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00030_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00030_00003;
wire [fgallag_WDTH-1:0]          fgallag_00030_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00030_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00030_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00030_00004;
wire [fgallag_WDTH-1:0]          fgallag_00030_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00030_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00030_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00030_00005;
wire [fgallag_WDTH-1:0]          fgallag_00031_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00031_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00031_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00031_00000;
wire [fgallag_WDTH-1:0]          fgallag_00031_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00031_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00031_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00031_00001;
wire [fgallag_WDTH-1:0]          fgallag_00031_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00031_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00031_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00031_00002;
wire [fgallag_WDTH-1:0]          fgallag_00031_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00031_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00031_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00031_00003;
wire [fgallag_WDTH-1:0]          fgallag_00031_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00031_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00031_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00031_00004;
wire [fgallag_WDTH-1:0]          fgallag_00031_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00031_00005;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00031_00005;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00031_00005;
wire [fgallag_WDTH-1:0]          fgallag_00032_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00032_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00032_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00032_00000;
wire [fgallag_WDTH-1:0]          fgallag_00032_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00032_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00032_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00032_00001;
wire [fgallag_WDTH-1:0]          fgallag_00032_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00032_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00032_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00032_00002;
wire [fgallag_WDTH-1:0]          fgallag_00032_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00032_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00032_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00032_00003;
wire [fgallag_WDTH-1:0]          fgallag_00033_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00033_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00033_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00033_00000;
wire [fgallag_WDTH-1:0]          fgallag_00033_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00033_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00033_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00033_00001;
wire [fgallag_WDTH-1:0]          fgallag_00033_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00033_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00033_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00033_00002;
wire [fgallag_WDTH-1:0]          fgallag_00033_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00033_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00033_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00033_00003;
wire [fgallag_WDTH-1:0]          fgallag_00034_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00034_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00034_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00034_00000;
wire [fgallag_WDTH-1:0]          fgallag_00034_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00034_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00034_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00034_00001;
wire [fgallag_WDTH-1:0]          fgallag_00034_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00034_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00034_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00034_00002;
wire [fgallag_WDTH-1:0]          fgallag_00034_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00034_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00034_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00034_00003;
wire [fgallag_WDTH-1:0]          fgallag_00035_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00035_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00035_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00035_00000;
wire [fgallag_WDTH-1:0]          fgallag_00035_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00035_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00035_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00035_00001;
wire [fgallag_WDTH-1:0]          fgallag_00035_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00035_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00035_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00035_00002;
wire [fgallag_WDTH-1:0]          fgallag_00035_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00035_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00035_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00035_00003;
wire [fgallag_WDTH-1:0]          fgallag_00036_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00036_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00036_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00036_00000;
wire [fgallag_WDTH-1:0]          fgallag_00036_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00036_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00036_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00036_00001;
wire [fgallag_WDTH-1:0]          fgallag_00036_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00036_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00036_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00036_00002;
wire [fgallag_WDTH-1:0]          fgallag_00036_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00036_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00036_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00036_00003;
wire [fgallag_WDTH-1:0]          fgallag_00036_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00036_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00036_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00036_00004;
wire [fgallag_WDTH-1:0]          fgallag_00037_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00037_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00037_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00037_00000;
wire [fgallag_WDTH-1:0]          fgallag_00037_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00037_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00037_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00037_00001;
wire [fgallag_WDTH-1:0]          fgallag_00037_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00037_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00037_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00037_00002;
wire [fgallag_WDTH-1:0]          fgallag_00037_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00037_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00037_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00037_00003;
wire [fgallag_WDTH-1:0]          fgallag_00037_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00037_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00037_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00037_00004;
wire [fgallag_WDTH-1:0]          fgallag_00038_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00038_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00038_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00038_00000;
wire [fgallag_WDTH-1:0]          fgallag_00038_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00038_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00038_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00038_00001;
wire [fgallag_WDTH-1:0]          fgallag_00038_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00038_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00038_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00038_00002;
wire [fgallag_WDTH-1:0]          fgallag_00038_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00038_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00038_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00038_00003;
wire [fgallag_WDTH-1:0]          fgallag_00038_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00038_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00038_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00038_00004;
wire [fgallag_WDTH-1:0]          fgallag_00039_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00039_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00039_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00039_00000;
wire [fgallag_WDTH-1:0]          fgallag_00039_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00039_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00039_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00039_00001;
wire [fgallag_WDTH-1:0]          fgallag_00039_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00039_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00039_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00039_00002;
wire [fgallag_WDTH-1:0]          fgallag_00039_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00039_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00039_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00039_00003;
wire [fgallag_WDTH-1:0]          fgallag_00039_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00039_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00039_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00039_00004;
wire [fgallag_WDTH-1:0]          fgallag_00040_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00040_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00040_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00040_00000;
wire [fgallag_WDTH-1:0]          fgallag_00040_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00040_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00040_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00040_00001;
wire [fgallag_WDTH-1:0]          fgallag_00040_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00040_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00040_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00040_00002;
wire [fgallag_WDTH-1:0]          fgallag_00040_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00040_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00040_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00040_00003;
wire [fgallag_WDTH-1:0]          fgallag_00040_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00040_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00040_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00040_00004;
wire [fgallag_WDTH-1:0]          fgallag_00041_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00041_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00041_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00041_00000;
wire [fgallag_WDTH-1:0]          fgallag_00041_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00041_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00041_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00041_00001;
wire [fgallag_WDTH-1:0]          fgallag_00041_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00041_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00041_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00041_00002;
wire [fgallag_WDTH-1:0]          fgallag_00041_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00041_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00041_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00041_00003;
wire [fgallag_WDTH-1:0]          fgallag_00041_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00041_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00041_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00041_00004;
wire [fgallag_WDTH-1:0]          fgallag_00042_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00042_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00042_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00042_00000;
wire [fgallag_WDTH-1:0]          fgallag_00042_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00042_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00042_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00042_00001;
wire [fgallag_WDTH-1:0]          fgallag_00042_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00042_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00042_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00042_00002;
wire [fgallag_WDTH-1:0]          fgallag_00042_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00042_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00042_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00042_00003;
wire [fgallag_WDTH-1:0]          fgallag_00042_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00042_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00042_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00042_00004;
wire [fgallag_WDTH-1:0]          fgallag_00043_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00043_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00043_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00043_00000;
wire [fgallag_WDTH-1:0]          fgallag_00043_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00043_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00043_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00043_00001;
wire [fgallag_WDTH-1:0]          fgallag_00043_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00043_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00043_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00043_00002;
wire [fgallag_WDTH-1:0]          fgallag_00043_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00043_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00043_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00043_00003;
wire [fgallag_WDTH-1:0]          fgallag_00043_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00043_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00043_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00043_00004;
wire [fgallag_WDTH-1:0]          fgallag_00044_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00044_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00044_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00044_00000;
wire [fgallag_WDTH-1:0]          fgallag_00044_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00044_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00044_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00044_00001;
wire [fgallag_WDTH-1:0]          fgallag_00044_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00044_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00044_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00044_00002;
wire [fgallag_WDTH-1:0]          fgallag_00044_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00044_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00044_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00044_00003;
wire [fgallag_WDTH-1:0]          fgallag_00044_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00044_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00044_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00044_00004;
wire [fgallag_WDTH-1:0]          fgallag_00045_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00045_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00045_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00045_00000;
wire [fgallag_WDTH-1:0]          fgallag_00045_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00045_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00045_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00045_00001;
wire [fgallag_WDTH-1:0]          fgallag_00045_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00045_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00045_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00045_00002;
wire [fgallag_WDTH-1:0]          fgallag_00045_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00045_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00045_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00045_00003;
wire [fgallag_WDTH-1:0]          fgallag_00045_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00045_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00045_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00045_00004;
wire [fgallag_WDTH-1:0]          fgallag_00046_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00046_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00046_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00046_00000;
wire [fgallag_WDTH-1:0]          fgallag_00046_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00046_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00046_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00046_00001;
wire [fgallag_WDTH-1:0]          fgallag_00046_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00046_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00046_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00046_00002;
wire [fgallag_WDTH-1:0]          fgallag_00046_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00046_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00046_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00046_00003;
wire [fgallag_WDTH-1:0]          fgallag_00046_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00046_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00046_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00046_00004;
wire [fgallag_WDTH-1:0]          fgallag_00047_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00047_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00047_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00047_00000;
wire [fgallag_WDTH-1:0]          fgallag_00047_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00047_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00047_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00047_00001;
wire [fgallag_WDTH-1:0]          fgallag_00047_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00047_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00047_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00047_00002;
wire [fgallag_WDTH-1:0]          fgallag_00047_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00047_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00047_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00047_00003;
wire [fgallag_WDTH-1:0]          fgallag_00047_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00047_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00047_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00047_00004;
wire [fgallag_WDTH-1:0]          fgallag_00048_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00048_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00048_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00048_00000;
wire [fgallag_WDTH-1:0]          fgallag_00048_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00048_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00048_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00048_00001;
wire [fgallag_WDTH-1:0]          fgallag_00048_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00048_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00048_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00048_00002;
wire [fgallag_WDTH-1:0]          fgallag_00048_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00048_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00048_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00048_00003;
wire [fgallag_WDTH-1:0]          fgallag_00049_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00049_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00049_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00049_00000;
wire [fgallag_WDTH-1:0]          fgallag_00049_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00049_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00049_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00049_00001;
wire [fgallag_WDTH-1:0]          fgallag_00049_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00049_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00049_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00049_00002;
wire [fgallag_WDTH-1:0]          fgallag_00049_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00049_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00049_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00049_00003;
wire [fgallag_WDTH-1:0]          fgallag_00050_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00050_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00050_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00050_00000;
wire [fgallag_WDTH-1:0]          fgallag_00050_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00050_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00050_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00050_00001;
wire [fgallag_WDTH-1:0]          fgallag_00050_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00050_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00050_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00050_00002;
wire [fgallag_WDTH-1:0]          fgallag_00050_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00050_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00050_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00050_00003;
wire [fgallag_WDTH-1:0]          fgallag_00051_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00051_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00051_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00051_00000;
wire [fgallag_WDTH-1:0]          fgallag_00051_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00051_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00051_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00051_00001;
wire [fgallag_WDTH-1:0]          fgallag_00051_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00051_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00051_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00051_00002;
wire [fgallag_WDTH-1:0]          fgallag_00051_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00051_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00051_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00051_00003;
wire [fgallag_WDTH-1:0]          fgallag_00052_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00052_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00052_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00052_00000;
wire [fgallag_WDTH-1:0]          fgallag_00052_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00052_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00052_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00052_00001;
wire [fgallag_WDTH-1:0]          fgallag_00052_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00052_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00052_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00052_00002;
wire [fgallag_WDTH-1:0]          fgallag_00052_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00052_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00052_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00052_00003;
wire [fgallag_WDTH-1:0]          fgallag_00052_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00052_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00052_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00052_00004;
wire [fgallag_WDTH-1:0]          fgallag_00053_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00053_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00053_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00053_00000;
wire [fgallag_WDTH-1:0]          fgallag_00053_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00053_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00053_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00053_00001;
wire [fgallag_WDTH-1:0]          fgallag_00053_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00053_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00053_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00053_00002;
wire [fgallag_WDTH-1:0]          fgallag_00053_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00053_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00053_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00053_00003;
wire [fgallag_WDTH-1:0]          fgallag_00053_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00053_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00053_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00053_00004;
wire [fgallag_WDTH-1:0]          fgallag_00054_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00054_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00054_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00054_00000;
wire [fgallag_WDTH-1:0]          fgallag_00054_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00054_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00054_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00054_00001;
wire [fgallag_WDTH-1:0]          fgallag_00054_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00054_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00054_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00054_00002;
wire [fgallag_WDTH-1:0]          fgallag_00054_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00054_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00054_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00054_00003;
wire [fgallag_WDTH-1:0]          fgallag_00054_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00054_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00054_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00054_00004;
wire [fgallag_WDTH-1:0]          fgallag_00055_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00055_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00055_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00055_00000;
wire [fgallag_WDTH-1:0]          fgallag_00055_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00055_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00055_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00055_00001;
wire [fgallag_WDTH-1:0]          fgallag_00055_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00055_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00055_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00055_00002;
wire [fgallag_WDTH-1:0]          fgallag_00055_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00055_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00055_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00055_00003;
wire [fgallag_WDTH-1:0]          fgallag_00055_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00055_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00055_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00055_00004;
wire [fgallag_WDTH-1:0]          fgallag_00056_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00056_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00056_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00056_00000;
wire [fgallag_WDTH-1:0]          fgallag_00056_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00056_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00056_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00056_00001;
wire [fgallag_WDTH-1:0]          fgallag_00056_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00056_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00056_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00056_00002;
wire [fgallag_WDTH-1:0]          fgallag_00056_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00056_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00056_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00056_00003;
wire [fgallag_WDTH-1:0]          fgallag_00056_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00056_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00056_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00056_00004;
wire [fgallag_WDTH-1:0]          fgallag_00057_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00057_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00057_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00057_00000;
wire [fgallag_WDTH-1:0]          fgallag_00057_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00057_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00057_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00057_00001;
wire [fgallag_WDTH-1:0]          fgallag_00057_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00057_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00057_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00057_00002;
wire [fgallag_WDTH-1:0]          fgallag_00057_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00057_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00057_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00057_00003;
wire [fgallag_WDTH-1:0]          fgallag_00057_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00057_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00057_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00057_00004;
wire [fgallag_WDTH-1:0]          fgallag_00058_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00058_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00058_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00058_00000;
wire [fgallag_WDTH-1:0]          fgallag_00058_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00058_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00058_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00058_00001;
wire [fgallag_WDTH-1:0]          fgallag_00058_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00058_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00058_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00058_00002;
wire [fgallag_WDTH-1:0]          fgallag_00058_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00058_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00058_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00058_00003;
wire [fgallag_WDTH-1:0]          fgallag_00058_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00058_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00058_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00058_00004;
wire [fgallag_WDTH-1:0]          fgallag_00059_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00059_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00059_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00059_00000;
wire [fgallag_WDTH-1:0]          fgallag_00059_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00059_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00059_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00059_00001;
wire [fgallag_WDTH-1:0]          fgallag_00059_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00059_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00059_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00059_00002;
wire [fgallag_WDTH-1:0]          fgallag_00059_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00059_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00059_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00059_00003;
wire [fgallag_WDTH-1:0]          fgallag_00059_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00059_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00059_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00059_00004;
wire [fgallag_WDTH-1:0]          fgallag_00060_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00060_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00060_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00060_00000;
wire [fgallag_WDTH-1:0]          fgallag_00060_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00060_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00060_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00060_00001;
wire [fgallag_WDTH-1:0]          fgallag_00060_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00060_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00060_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00060_00002;
wire [fgallag_WDTH-1:0]          fgallag_00060_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00060_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00060_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00060_00003;
wire [fgallag_WDTH-1:0]          fgallag_00061_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00061_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00061_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00061_00000;
wire [fgallag_WDTH-1:0]          fgallag_00061_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00061_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00061_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00061_00001;
wire [fgallag_WDTH-1:0]          fgallag_00061_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00061_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00061_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00061_00002;
wire [fgallag_WDTH-1:0]          fgallag_00061_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00061_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00061_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00061_00003;
wire [fgallag_WDTH-1:0]          fgallag_00062_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00062_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00062_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00062_00000;
wire [fgallag_WDTH-1:0]          fgallag_00062_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00062_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00062_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00062_00001;
wire [fgallag_WDTH-1:0]          fgallag_00062_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00062_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00062_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00062_00002;
wire [fgallag_WDTH-1:0]          fgallag_00062_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00062_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00062_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00062_00003;
wire [fgallag_WDTH-1:0]          fgallag_00063_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00063_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00063_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00063_00000;
wire [fgallag_WDTH-1:0]          fgallag_00063_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00063_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00063_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00063_00001;
wire [fgallag_WDTH-1:0]          fgallag_00063_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00063_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00063_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00063_00002;
wire [fgallag_WDTH-1:0]          fgallag_00063_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00063_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00063_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00063_00003;
wire [fgallag_WDTH-1:0]          fgallag_00064_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00064_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00064_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00064_00000;
wire [fgallag_WDTH-1:0]          fgallag_00064_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00064_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00064_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00064_00001;
wire [fgallag_WDTH-1:0]          fgallag_00064_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00064_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00064_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00064_00002;
wire [fgallag_WDTH-1:0]          fgallag_00064_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00064_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00064_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00064_00003;
wire [fgallag_WDTH-1:0]          fgallag_00064_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00064_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00064_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00064_00004;
wire [fgallag_WDTH-1:0]          fgallag_00065_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00065_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00065_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00065_00000;
wire [fgallag_WDTH-1:0]          fgallag_00065_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00065_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00065_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00065_00001;
wire [fgallag_WDTH-1:0]          fgallag_00065_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00065_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00065_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00065_00002;
wire [fgallag_WDTH-1:0]          fgallag_00065_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00065_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00065_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00065_00003;
wire [fgallag_WDTH-1:0]          fgallag_00065_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00065_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00065_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00065_00004;
wire [fgallag_WDTH-1:0]          fgallag_00066_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00066_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00066_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00066_00000;
wire [fgallag_WDTH-1:0]          fgallag_00066_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00066_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00066_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00066_00001;
wire [fgallag_WDTH-1:0]          fgallag_00066_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00066_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00066_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00066_00002;
wire [fgallag_WDTH-1:0]          fgallag_00066_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00066_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00066_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00066_00003;
wire [fgallag_WDTH-1:0]          fgallag_00066_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00066_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00066_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00066_00004;
wire [fgallag_WDTH-1:0]          fgallag_00067_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00067_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00067_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00067_00000;
wire [fgallag_WDTH-1:0]          fgallag_00067_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00067_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00067_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00067_00001;
wire [fgallag_WDTH-1:0]          fgallag_00067_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00067_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00067_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00067_00002;
wire [fgallag_WDTH-1:0]          fgallag_00067_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00067_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00067_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00067_00003;
wire [fgallag_WDTH-1:0]          fgallag_00067_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00067_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00067_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00067_00004;
wire [fgallag_WDTH-1:0]          fgallag_00068_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00068_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00068_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00068_00000;
wire [fgallag_WDTH-1:0]          fgallag_00068_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00068_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00068_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00068_00001;
wire [fgallag_WDTH-1:0]          fgallag_00068_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00068_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00068_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00068_00002;
wire [fgallag_WDTH-1:0]          fgallag_00068_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00068_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00068_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00068_00003;
wire [fgallag_WDTH-1:0]          fgallag_00068_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00068_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00068_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00068_00004;
wire [fgallag_WDTH-1:0]          fgallag_00069_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00069_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00069_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00069_00000;
wire [fgallag_WDTH-1:0]          fgallag_00069_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00069_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00069_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00069_00001;
wire [fgallag_WDTH-1:0]          fgallag_00069_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00069_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00069_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00069_00002;
wire [fgallag_WDTH-1:0]          fgallag_00069_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00069_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00069_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00069_00003;
wire [fgallag_WDTH-1:0]          fgallag_00069_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00069_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00069_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00069_00004;
wire [fgallag_WDTH-1:0]          fgallag_00070_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00070_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00070_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00070_00000;
wire [fgallag_WDTH-1:0]          fgallag_00070_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00070_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00070_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00070_00001;
wire [fgallag_WDTH-1:0]          fgallag_00070_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00070_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00070_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00070_00002;
wire [fgallag_WDTH-1:0]          fgallag_00070_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00070_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00070_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00070_00003;
wire [fgallag_WDTH-1:0]          fgallag_00070_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00070_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00070_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00070_00004;
wire [fgallag_WDTH-1:0]          fgallag_00071_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00071_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00071_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00071_00000;
wire [fgallag_WDTH-1:0]          fgallag_00071_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00071_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00071_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00071_00001;
wire [fgallag_WDTH-1:0]          fgallag_00071_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00071_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00071_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00071_00002;
wire [fgallag_WDTH-1:0]          fgallag_00071_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00071_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00071_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00071_00003;
wire [fgallag_WDTH-1:0]          fgallag_00071_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00071_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00071_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00071_00004;
wire [fgallag_WDTH-1:0]          fgallag_00072_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00072_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00072_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00072_00000;
wire [fgallag_WDTH-1:0]          fgallag_00072_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00072_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00072_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00072_00001;
wire [fgallag_WDTH-1:0]          fgallag_00072_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00072_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00072_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00072_00002;
wire [fgallag_WDTH-1:0]          fgallag_00072_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00072_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00072_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00072_00003;
wire [fgallag_WDTH-1:0]          fgallag_00073_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00073_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00073_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00073_00000;
wire [fgallag_WDTH-1:0]          fgallag_00073_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00073_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00073_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00073_00001;
wire [fgallag_WDTH-1:0]          fgallag_00073_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00073_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00073_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00073_00002;
wire [fgallag_WDTH-1:0]          fgallag_00073_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00073_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00073_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00073_00003;
wire [fgallag_WDTH-1:0]          fgallag_00074_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00074_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00074_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00074_00000;
wire [fgallag_WDTH-1:0]          fgallag_00074_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00074_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00074_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00074_00001;
wire [fgallag_WDTH-1:0]          fgallag_00074_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00074_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00074_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00074_00002;
wire [fgallag_WDTH-1:0]          fgallag_00074_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00074_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00074_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00074_00003;
wire [fgallag_WDTH-1:0]          fgallag_00075_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00075_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00075_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00075_00000;
wire [fgallag_WDTH-1:0]          fgallag_00075_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00075_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00075_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00075_00001;
wire [fgallag_WDTH-1:0]          fgallag_00075_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00075_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00075_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00075_00002;
wire [fgallag_WDTH-1:0]          fgallag_00075_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00075_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00075_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00075_00003;
wire [fgallag_WDTH-1:0]          fgallag_00076_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00076_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00076_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00076_00000;
wire [fgallag_WDTH-1:0]          fgallag_00076_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00076_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00076_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00076_00001;
wire [fgallag_WDTH-1:0]          fgallag_00076_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00076_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00076_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00076_00002;
wire [fgallag_WDTH-1:0]          fgallag_00076_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00076_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00076_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00076_00003;
wire [fgallag_WDTH-1:0]          fgallag_00077_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00077_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00077_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00077_00000;
wire [fgallag_WDTH-1:0]          fgallag_00077_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00077_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00077_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00077_00001;
wire [fgallag_WDTH-1:0]          fgallag_00077_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00077_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00077_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00077_00002;
wire [fgallag_WDTH-1:0]          fgallag_00077_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00077_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00077_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00077_00003;
wire [fgallag_WDTH-1:0]          fgallag_00078_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00078_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00078_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00078_00000;
wire [fgallag_WDTH-1:0]          fgallag_00078_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00078_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00078_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00078_00001;
wire [fgallag_WDTH-1:0]          fgallag_00078_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00078_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00078_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00078_00002;
wire [fgallag_WDTH-1:0]          fgallag_00078_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00078_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00078_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00078_00003;
wire [fgallag_WDTH-1:0]          fgallag_00079_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00079_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00079_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00079_00000;
wire [fgallag_WDTH-1:0]          fgallag_00079_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00079_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00079_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00079_00001;
wire [fgallag_WDTH-1:0]          fgallag_00079_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00079_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00079_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00079_00002;
wire [fgallag_WDTH-1:0]          fgallag_00079_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00079_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00079_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00079_00003;
wire [fgallag_WDTH-1:0]          fgallag_00080_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00080_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00080_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00080_00000;
wire [fgallag_WDTH-1:0]          fgallag_00080_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00080_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00080_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00080_00001;
wire [fgallag_WDTH-1:0]          fgallag_00080_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00080_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00080_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00080_00002;
wire [fgallag_WDTH-1:0]          fgallag_00080_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00080_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00080_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00080_00003;
wire [fgallag_WDTH-1:0]          fgallag_00081_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00081_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00081_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00081_00000;
wire [fgallag_WDTH-1:0]          fgallag_00081_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00081_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00081_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00081_00001;
wire [fgallag_WDTH-1:0]          fgallag_00081_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00081_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00081_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00081_00002;
wire [fgallag_WDTH-1:0]          fgallag_00081_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00081_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00081_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00081_00003;
wire [fgallag_WDTH-1:0]          fgallag_00082_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00082_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00082_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00082_00000;
wire [fgallag_WDTH-1:0]          fgallag_00082_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00082_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00082_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00082_00001;
wire [fgallag_WDTH-1:0]          fgallag_00082_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00082_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00082_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00082_00002;
wire [fgallag_WDTH-1:0]          fgallag_00082_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00082_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00082_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00082_00003;
wire [fgallag_WDTH-1:0]          fgallag_00083_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00083_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00083_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00083_00000;
wire [fgallag_WDTH-1:0]          fgallag_00083_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00083_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00083_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00083_00001;
wire [fgallag_WDTH-1:0]          fgallag_00083_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00083_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00083_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00083_00002;
wire [fgallag_WDTH-1:0]          fgallag_00083_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00083_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00083_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00083_00003;
wire [fgallag_WDTH-1:0]          fgallag_00084_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00084_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00084_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00084_00000;
wire [fgallag_WDTH-1:0]          fgallag_00084_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00084_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00084_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00084_00001;
wire [fgallag_WDTH-1:0]          fgallag_00084_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00084_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00084_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00084_00002;
wire [fgallag_WDTH-1:0]          fgallag_00084_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00084_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00084_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00084_00003;
wire [fgallag_WDTH-1:0]          fgallag_00085_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00085_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00085_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00085_00000;
wire [fgallag_WDTH-1:0]          fgallag_00085_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00085_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00085_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00085_00001;
wire [fgallag_WDTH-1:0]          fgallag_00085_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00085_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00085_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00085_00002;
wire [fgallag_WDTH-1:0]          fgallag_00085_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00085_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00085_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00085_00003;
wire [fgallag_WDTH-1:0]          fgallag_00086_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00086_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00086_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00086_00000;
wire [fgallag_WDTH-1:0]          fgallag_00086_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00086_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00086_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00086_00001;
wire [fgallag_WDTH-1:0]          fgallag_00086_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00086_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00086_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00086_00002;
wire [fgallag_WDTH-1:0]          fgallag_00086_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00086_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00086_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00086_00003;
wire [fgallag_WDTH-1:0]          fgallag_00087_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00087_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00087_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00087_00000;
wire [fgallag_WDTH-1:0]          fgallag_00087_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00087_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00087_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00087_00001;
wire [fgallag_WDTH-1:0]          fgallag_00087_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00087_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00087_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00087_00002;
wire [fgallag_WDTH-1:0]          fgallag_00087_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00087_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00087_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00087_00003;
wire [fgallag_WDTH-1:0]          fgallag_00088_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00088_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00088_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00088_00000;
wire [fgallag_WDTH-1:0]          fgallag_00088_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00088_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00088_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00088_00001;
wire [fgallag_WDTH-1:0]          fgallag_00088_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00088_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00088_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00088_00002;
wire [fgallag_WDTH-1:0]          fgallag_00089_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00089_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00089_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00089_00000;
wire [fgallag_WDTH-1:0]          fgallag_00089_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00089_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00089_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00089_00001;
wire [fgallag_WDTH-1:0]          fgallag_00089_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00089_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00089_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00089_00002;
wire [fgallag_WDTH-1:0]          fgallag_00090_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00090_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00090_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00090_00000;
wire [fgallag_WDTH-1:0]          fgallag_00090_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00090_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00090_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00090_00001;
wire [fgallag_WDTH-1:0]          fgallag_00090_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00090_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00090_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00090_00002;
wire [fgallag_WDTH-1:0]          fgallag_00091_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00091_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00091_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00091_00000;
wire [fgallag_WDTH-1:0]          fgallag_00091_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00091_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00091_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00091_00001;
wire [fgallag_WDTH-1:0]          fgallag_00091_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00091_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00091_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00091_00002;
wire [fgallag_WDTH-1:0]          fgallag_00092_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00092_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00092_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00092_00000;
wire [fgallag_WDTH-1:0]          fgallag_00092_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00092_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00092_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00092_00001;
wire [fgallag_WDTH-1:0]          fgallag_00092_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00092_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00092_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00092_00002;
wire [fgallag_WDTH-1:0]          fgallag_00092_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00092_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00092_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00092_00003;
wire [fgallag_WDTH-1:0]          fgallag_00093_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00093_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00093_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00093_00000;
wire [fgallag_WDTH-1:0]          fgallag_00093_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00093_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00093_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00093_00001;
wire [fgallag_WDTH-1:0]          fgallag_00093_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00093_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00093_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00093_00002;
wire [fgallag_WDTH-1:0]          fgallag_00093_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00093_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00093_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00093_00003;
wire [fgallag_WDTH-1:0]          fgallag_00094_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00094_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00094_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00094_00000;
wire [fgallag_WDTH-1:0]          fgallag_00094_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00094_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00094_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00094_00001;
wire [fgallag_WDTH-1:0]          fgallag_00094_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00094_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00094_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00094_00002;
wire [fgallag_WDTH-1:0]          fgallag_00094_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00094_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00094_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00094_00003;
wire [fgallag_WDTH-1:0]          fgallag_00095_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00095_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00095_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00095_00000;
wire [fgallag_WDTH-1:0]          fgallag_00095_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00095_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00095_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00095_00001;
wire [fgallag_WDTH-1:0]          fgallag_00095_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00095_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00095_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00095_00002;
wire [fgallag_WDTH-1:0]          fgallag_00095_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00095_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00095_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00095_00003;
wire [fgallag_WDTH-1:0]          fgallag_00096_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00096_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00096_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00096_00000;
wire [fgallag_WDTH-1:0]          fgallag_00096_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00096_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00096_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00096_00001;
wire [fgallag_WDTH-1:0]          fgallag_00096_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00096_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00096_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00096_00002;
wire [fgallag_WDTH-1:0]          fgallag_00096_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00096_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00096_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00096_00003;
wire [fgallag_WDTH-1:0]          fgallag_00097_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00097_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00097_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00097_00000;
wire [fgallag_WDTH-1:0]          fgallag_00097_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00097_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00097_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00097_00001;
wire [fgallag_WDTH-1:0]          fgallag_00097_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00097_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00097_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00097_00002;
wire [fgallag_WDTH-1:0]          fgallag_00097_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00097_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00097_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00097_00003;
wire [fgallag_WDTH-1:0]          fgallag_00098_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00098_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00098_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00098_00000;
wire [fgallag_WDTH-1:0]          fgallag_00098_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00098_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00098_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00098_00001;
wire [fgallag_WDTH-1:0]          fgallag_00098_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00098_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00098_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00098_00002;
wire [fgallag_WDTH-1:0]          fgallag_00098_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00098_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00098_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00098_00003;
wire [fgallag_WDTH-1:0]          fgallag_00099_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00099_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00099_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00099_00000;
wire [fgallag_WDTH-1:0]          fgallag_00099_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00099_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00099_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00099_00001;
wire [fgallag_WDTH-1:0]          fgallag_00099_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00099_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00099_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00099_00002;
wire [fgallag_WDTH-1:0]          fgallag_00099_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00099_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00099_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00099_00003;
wire [fgallag_WDTH-1:0]          fgallag_00100_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00100_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00100_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00100_00000;
wire [fgallag_WDTH-1:0]          fgallag_00100_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00100_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00100_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00100_00001;
wire [fgallag_WDTH-1:0]          fgallag_00100_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00100_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00100_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00100_00002;
wire [fgallag_WDTH-1:0]          fgallag_00101_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00101_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00101_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00101_00000;
wire [fgallag_WDTH-1:0]          fgallag_00101_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00101_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00101_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00101_00001;
wire [fgallag_WDTH-1:0]          fgallag_00101_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00101_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00101_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00101_00002;
wire [fgallag_WDTH-1:0]          fgallag_00102_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00102_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00102_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00102_00000;
wire [fgallag_WDTH-1:0]          fgallag_00102_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00102_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00102_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00102_00001;
wire [fgallag_WDTH-1:0]          fgallag_00102_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00102_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00102_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00102_00002;
wire [fgallag_WDTH-1:0]          fgallag_00103_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00103_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00103_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00103_00000;
wire [fgallag_WDTH-1:0]          fgallag_00103_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00103_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00103_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00103_00001;
wire [fgallag_WDTH-1:0]          fgallag_00103_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00103_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00103_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00103_00002;
wire [fgallag_WDTH-1:0]          fgallag_00104_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00104_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00104_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00104_00000;
wire [fgallag_WDTH-1:0]          fgallag_00104_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00104_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00104_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00104_00001;
wire [fgallag_WDTH-1:0]          fgallag_00104_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00104_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00104_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00104_00002;
wire [fgallag_WDTH-1:0]          fgallag_00104_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00104_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00104_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00104_00003;
wire [fgallag_WDTH-1:0]          fgallag_00104_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00104_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00104_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00104_00004;
wire [fgallag_WDTH-1:0]          fgallag_00105_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00105_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00105_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00105_00000;
wire [fgallag_WDTH-1:0]          fgallag_00105_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00105_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00105_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00105_00001;
wire [fgallag_WDTH-1:0]          fgallag_00105_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00105_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00105_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00105_00002;
wire [fgallag_WDTH-1:0]          fgallag_00105_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00105_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00105_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00105_00003;
wire [fgallag_WDTH-1:0]          fgallag_00105_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00105_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00105_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00105_00004;
wire [fgallag_WDTH-1:0]          fgallag_00106_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00106_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00106_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00106_00000;
wire [fgallag_WDTH-1:0]          fgallag_00106_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00106_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00106_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00106_00001;
wire [fgallag_WDTH-1:0]          fgallag_00106_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00106_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00106_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00106_00002;
wire [fgallag_WDTH-1:0]          fgallag_00106_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00106_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00106_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00106_00003;
wire [fgallag_WDTH-1:0]          fgallag_00106_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00106_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00106_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00106_00004;
wire [fgallag_WDTH-1:0]          fgallag_00107_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00107_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00107_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00107_00000;
wire [fgallag_WDTH-1:0]          fgallag_00107_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00107_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00107_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00107_00001;
wire [fgallag_WDTH-1:0]          fgallag_00107_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00107_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00107_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00107_00002;
wire [fgallag_WDTH-1:0]          fgallag_00107_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00107_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00107_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00107_00003;
wire [fgallag_WDTH-1:0]          fgallag_00107_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00107_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00107_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00107_00004;
wire [fgallag_WDTH-1:0]          fgallag_00108_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00108_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00108_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00108_00000;
wire [fgallag_WDTH-1:0]          fgallag_00108_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00108_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00108_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00108_00001;
wire [fgallag_WDTH-1:0]          fgallag_00108_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00108_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00108_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00108_00002;
wire [fgallag_WDTH-1:0]          fgallag_00109_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00109_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00109_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00109_00000;
wire [fgallag_WDTH-1:0]          fgallag_00109_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00109_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00109_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00109_00001;
wire [fgallag_WDTH-1:0]          fgallag_00109_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00109_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00109_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00109_00002;
wire [fgallag_WDTH-1:0]          fgallag_00110_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00110_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00110_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00110_00000;
wire [fgallag_WDTH-1:0]          fgallag_00110_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00110_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00110_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00110_00001;
wire [fgallag_WDTH-1:0]          fgallag_00110_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00110_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00110_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00110_00002;
wire [fgallag_WDTH-1:0]          fgallag_00111_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00111_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00111_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00111_00000;
wire [fgallag_WDTH-1:0]          fgallag_00111_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00111_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00111_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00111_00001;
wire [fgallag_WDTH-1:0]          fgallag_00111_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00111_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00111_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00111_00002;
wire [fgallag_WDTH-1:0]          fgallag_00112_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00112_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00112_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00112_00000;
wire [fgallag_WDTH-1:0]          fgallag_00112_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00112_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00112_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00112_00001;
wire [fgallag_WDTH-1:0]          fgallag_00112_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00112_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00112_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00112_00002;
wire [fgallag_WDTH-1:0]          fgallag_00112_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00112_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00112_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00112_00003;
wire [fgallag_WDTH-1:0]          fgallag_00113_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00113_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00113_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00113_00000;
wire [fgallag_WDTH-1:0]          fgallag_00113_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00113_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00113_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00113_00001;
wire [fgallag_WDTH-1:0]          fgallag_00113_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00113_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00113_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00113_00002;
wire [fgallag_WDTH-1:0]          fgallag_00113_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00113_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00113_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00113_00003;
wire [fgallag_WDTH-1:0]          fgallag_00114_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00114_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00114_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00114_00000;
wire [fgallag_WDTH-1:0]          fgallag_00114_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00114_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00114_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00114_00001;
wire [fgallag_WDTH-1:0]          fgallag_00114_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00114_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00114_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00114_00002;
wire [fgallag_WDTH-1:0]          fgallag_00114_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00114_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00114_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00114_00003;
wire [fgallag_WDTH-1:0]          fgallag_00115_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00115_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00115_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00115_00000;
wire [fgallag_WDTH-1:0]          fgallag_00115_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00115_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00115_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00115_00001;
wire [fgallag_WDTH-1:0]          fgallag_00115_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00115_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00115_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00115_00002;
wire [fgallag_WDTH-1:0]          fgallag_00115_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00115_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00115_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00115_00003;
wire [fgallag_WDTH-1:0]          fgallag_00116_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00116_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00116_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00116_00000;
wire [fgallag_WDTH-1:0]          fgallag_00116_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00116_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00116_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00116_00001;
wire [fgallag_WDTH-1:0]          fgallag_00116_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00116_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00116_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00116_00002;
wire [fgallag_WDTH-1:0]          fgallag_00117_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00117_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00117_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00117_00000;
wire [fgallag_WDTH-1:0]          fgallag_00117_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00117_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00117_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00117_00001;
wire [fgallag_WDTH-1:0]          fgallag_00117_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00117_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00117_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00117_00002;
wire [fgallag_WDTH-1:0]          fgallag_00118_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00118_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00118_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00118_00000;
wire [fgallag_WDTH-1:0]          fgallag_00118_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00118_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00118_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00118_00001;
wire [fgallag_WDTH-1:0]          fgallag_00118_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00118_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00118_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00118_00002;
wire [fgallag_WDTH-1:0]          fgallag_00119_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00119_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00119_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00119_00000;
wire [fgallag_WDTH-1:0]          fgallag_00119_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00119_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00119_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00119_00001;
wire [fgallag_WDTH-1:0]          fgallag_00119_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00119_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00119_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00119_00002;
wire [fgallag_WDTH-1:0]          fgallag_00120_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00120_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00120_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00120_00000;
wire [fgallag_WDTH-1:0]          fgallag_00120_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00120_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00120_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00120_00001;
wire [fgallag_WDTH-1:0]          fgallag_00120_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00120_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00120_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00120_00002;
wire [fgallag_WDTH-1:0]          fgallag_00120_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00120_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00120_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00120_00003;
wire [fgallag_WDTH-1:0]          fgallag_00120_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00120_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00120_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00120_00004;
wire [fgallag_WDTH-1:0]          fgallag_00121_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00121_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00121_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00121_00000;
wire [fgallag_WDTH-1:0]          fgallag_00121_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00121_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00121_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00121_00001;
wire [fgallag_WDTH-1:0]          fgallag_00121_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00121_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00121_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00121_00002;
wire [fgallag_WDTH-1:0]          fgallag_00121_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00121_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00121_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00121_00003;
wire [fgallag_WDTH-1:0]          fgallag_00121_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00121_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00121_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00121_00004;
wire [fgallag_WDTH-1:0]          fgallag_00122_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00122_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00122_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00122_00000;
wire [fgallag_WDTH-1:0]          fgallag_00122_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00122_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00122_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00122_00001;
wire [fgallag_WDTH-1:0]          fgallag_00122_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00122_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00122_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00122_00002;
wire [fgallag_WDTH-1:0]          fgallag_00122_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00122_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00122_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00122_00003;
wire [fgallag_WDTH-1:0]          fgallag_00122_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00122_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00122_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00122_00004;
wire [fgallag_WDTH-1:0]          fgallag_00123_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00123_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00123_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00123_00000;
wire [fgallag_WDTH-1:0]          fgallag_00123_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00123_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00123_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00123_00001;
wire [fgallag_WDTH-1:0]          fgallag_00123_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00123_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00123_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00123_00002;
wire [fgallag_WDTH-1:0]          fgallag_00123_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00123_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00123_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00123_00003;
wire [fgallag_WDTH-1:0]          fgallag_00123_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00123_00004;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00123_00004;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00123_00004;
wire [fgallag_WDTH-1:0]          fgallag_00124_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00124_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00124_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00124_00000;
wire [fgallag_WDTH-1:0]          fgallag_00124_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00124_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00124_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00124_00001;
wire [fgallag_WDTH-1:0]          fgallag_00124_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00124_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00124_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00124_00002;
wire [fgallag_WDTH-1:0]          fgallag_00125_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00125_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00125_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00125_00000;
wire [fgallag_WDTH-1:0]          fgallag_00125_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00125_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00125_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00125_00001;
wire [fgallag_WDTH-1:0]          fgallag_00125_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00125_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00125_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00125_00002;
wire [fgallag_WDTH-1:0]          fgallag_00126_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00126_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00126_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00126_00000;
wire [fgallag_WDTH-1:0]          fgallag_00126_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00126_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00126_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00126_00001;
wire [fgallag_WDTH-1:0]          fgallag_00126_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00126_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00126_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00126_00002;
wire [fgallag_WDTH-1:0]          fgallag_00127_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00127_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00127_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00127_00000;
wire [fgallag_WDTH-1:0]          fgallag_00127_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00127_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00127_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00127_00001;
wire [fgallag_WDTH-1:0]          fgallag_00127_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00127_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00127_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00127_00002;
wire [fgallag_WDTH-1:0]          fgallag_00128_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00128_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00128_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00128_00000;
wire [fgallag_WDTH-1:0]          fgallag_00128_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00128_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00128_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00128_00001;
wire [fgallag_WDTH-1:0]          fgallag_00128_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00128_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00128_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00128_00002;
wire [fgallag_WDTH-1:0]          fgallag_00128_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00128_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00128_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00128_00003;
wire [fgallag_WDTH-1:0]          fgallag_00129_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00129_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00129_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00129_00000;
wire [fgallag_WDTH-1:0]          fgallag_00129_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00129_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00129_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00129_00001;
wire [fgallag_WDTH-1:0]          fgallag_00129_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00129_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00129_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00129_00002;
wire [fgallag_WDTH-1:0]          fgallag_00129_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00129_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00129_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00129_00003;
wire [fgallag_WDTH-1:0]          fgallag_00130_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00130_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00130_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00130_00000;
wire [fgallag_WDTH-1:0]          fgallag_00130_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00130_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00130_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00130_00001;
wire [fgallag_WDTH-1:0]          fgallag_00130_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00130_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00130_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00130_00002;
wire [fgallag_WDTH-1:0]          fgallag_00130_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00130_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00130_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00130_00003;
wire [fgallag_WDTH-1:0]          fgallag_00131_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00131_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00131_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00131_00000;
wire [fgallag_WDTH-1:0]          fgallag_00131_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00131_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00131_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00131_00001;
wire [fgallag_WDTH-1:0]          fgallag_00131_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00131_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00131_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00131_00002;
wire [fgallag_WDTH-1:0]          fgallag_00131_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00131_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00131_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00131_00003;
wire [fgallag_WDTH-1:0]          fgallag_00132_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00132_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00132_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00132_00000;
wire [fgallag_WDTH-1:0]          fgallag_00132_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00132_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00132_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00132_00001;
wire [fgallag_WDTH-1:0]          fgallag_00132_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00132_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00132_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00132_00002;
wire [fgallag_WDTH-1:0]          fgallag_00132_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00132_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00132_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00132_00003;
wire [fgallag_WDTH-1:0]          fgallag_00133_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00133_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00133_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00133_00000;
wire [fgallag_WDTH-1:0]          fgallag_00133_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00133_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00133_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00133_00001;
wire [fgallag_WDTH-1:0]          fgallag_00133_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00133_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00133_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00133_00002;
wire [fgallag_WDTH-1:0]          fgallag_00133_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00133_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00133_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00133_00003;
wire [fgallag_WDTH-1:0]          fgallag_00134_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00134_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00134_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00134_00000;
wire [fgallag_WDTH-1:0]          fgallag_00134_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00134_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00134_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00134_00001;
wire [fgallag_WDTH-1:0]          fgallag_00134_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00134_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00134_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00134_00002;
wire [fgallag_WDTH-1:0]          fgallag_00134_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00134_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00134_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00134_00003;
wire [fgallag_WDTH-1:0]          fgallag_00135_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00135_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00135_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00135_00000;
wire [fgallag_WDTH-1:0]          fgallag_00135_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00135_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00135_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00135_00001;
wire [fgallag_WDTH-1:0]          fgallag_00135_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00135_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00135_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00135_00002;
wire [fgallag_WDTH-1:0]          fgallag_00135_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00135_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00135_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00135_00003;
wire [fgallag_WDTH-1:0]          fgallag_00136_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00136_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00136_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00136_00000;
wire [fgallag_WDTH-1:0]          fgallag_00136_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00136_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00136_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00136_00001;
wire [fgallag_WDTH-1:0]          fgallag_00136_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00136_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00136_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00136_00002;
wire [fgallag_WDTH-1:0]          fgallag_00136_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00136_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00136_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00136_00003;
wire [fgallag_WDTH-1:0]          fgallag_00137_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00137_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00137_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00137_00000;
wire [fgallag_WDTH-1:0]          fgallag_00137_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00137_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00137_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00137_00001;
wire [fgallag_WDTH-1:0]          fgallag_00137_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00137_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00137_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00137_00002;
wire [fgallag_WDTH-1:0]          fgallag_00137_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00137_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00137_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00137_00003;
wire [fgallag_WDTH-1:0]          fgallag_00138_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00138_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00138_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00138_00000;
wire [fgallag_WDTH-1:0]          fgallag_00138_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00138_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00138_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00138_00001;
wire [fgallag_WDTH-1:0]          fgallag_00138_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00138_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00138_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00138_00002;
wire [fgallag_WDTH-1:0]          fgallag_00138_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00138_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00138_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00138_00003;
wire [fgallag_WDTH-1:0]          fgallag_00139_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00139_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00139_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00139_00000;
wire [fgallag_WDTH-1:0]          fgallag_00139_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00139_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00139_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00139_00001;
wire [fgallag_WDTH-1:0]          fgallag_00139_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00139_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00139_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00139_00002;
wire [fgallag_WDTH-1:0]          fgallag_00139_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00139_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00139_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00139_00003;
wire [fgallag_WDTH-1:0]          fgallag_00140_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00140_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00140_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00140_00000;
wire [fgallag_WDTH-1:0]          fgallag_00140_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00140_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00140_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00140_00001;
wire [fgallag_WDTH-1:0]          fgallag_00140_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00140_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00140_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00140_00002;
wire [fgallag_WDTH-1:0]          fgallag_00140_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00140_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00140_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00140_00003;
wire [fgallag_WDTH-1:0]          fgallag_00141_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00141_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00141_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00141_00000;
wire [fgallag_WDTH-1:0]          fgallag_00141_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00141_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00141_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00141_00001;
wire [fgallag_WDTH-1:0]          fgallag_00141_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00141_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00141_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00141_00002;
wire [fgallag_WDTH-1:0]          fgallag_00141_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00141_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00141_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00141_00003;
wire [fgallag_WDTH-1:0]          fgallag_00142_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00142_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00142_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00142_00000;
wire [fgallag_WDTH-1:0]          fgallag_00142_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00142_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00142_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00142_00001;
wire [fgallag_WDTH-1:0]          fgallag_00142_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00142_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00142_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00142_00002;
wire [fgallag_WDTH-1:0]          fgallag_00142_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00142_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00142_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00142_00003;
wire [fgallag_WDTH-1:0]          fgallag_00143_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00143_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00143_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00143_00000;
wire [fgallag_WDTH-1:0]          fgallag_00143_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00143_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00143_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00143_00001;
wire [fgallag_WDTH-1:0]          fgallag_00143_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00143_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00143_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00143_00002;
wire [fgallag_WDTH-1:0]          fgallag_00143_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00143_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00143_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00143_00003;
wire [fgallag_WDTH-1:0]          fgallag_00144_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00144_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00144_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00144_00000;
wire [fgallag_WDTH-1:0]          fgallag_00144_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00144_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00144_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00144_00001;
wire [fgallag_WDTH-1:0]          fgallag_00144_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00144_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00144_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00144_00002;
wire [fgallag_WDTH-1:0]          fgallag_00144_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00144_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00144_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00144_00003;
wire [fgallag_WDTH-1:0]          fgallag_00145_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00145_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00145_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00145_00000;
wire [fgallag_WDTH-1:0]          fgallag_00145_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00145_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00145_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00145_00001;
wire [fgallag_WDTH-1:0]          fgallag_00145_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00145_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00145_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00145_00002;
wire [fgallag_WDTH-1:0]          fgallag_00145_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00145_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00145_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00145_00003;
wire [fgallag_WDTH-1:0]          fgallag_00146_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00146_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00146_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00146_00000;
wire [fgallag_WDTH-1:0]          fgallag_00146_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00146_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00146_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00146_00001;
wire [fgallag_WDTH-1:0]          fgallag_00146_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00146_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00146_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00146_00002;
wire [fgallag_WDTH-1:0]          fgallag_00146_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00146_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00146_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00146_00003;
wire [fgallag_WDTH-1:0]          fgallag_00147_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00147_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00147_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00147_00000;
wire [fgallag_WDTH-1:0]          fgallag_00147_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00147_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00147_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00147_00001;
wire [fgallag_WDTH-1:0]          fgallag_00147_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00147_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00147_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00147_00002;
wire [fgallag_WDTH-1:0]          fgallag_00147_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00147_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00147_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00147_00003;
wire [fgallag_WDTH-1:0]          fgallag_00148_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00148_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00148_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00148_00000;
wire [fgallag_WDTH-1:0]          fgallag_00148_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00148_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00148_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00148_00001;
wire [fgallag_WDTH-1:0]          fgallag_00148_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00148_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00148_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00148_00002;
wire [fgallag_WDTH-1:0]          fgallag_00149_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00149_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00149_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00149_00000;
wire [fgallag_WDTH-1:0]          fgallag_00149_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00149_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00149_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00149_00001;
wire [fgallag_WDTH-1:0]          fgallag_00149_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00149_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00149_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00149_00002;
wire [fgallag_WDTH-1:0]          fgallag_00150_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00150_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00150_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00150_00000;
wire [fgallag_WDTH-1:0]          fgallag_00150_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00150_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00150_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00150_00001;
wire [fgallag_WDTH-1:0]          fgallag_00150_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00150_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00150_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00150_00002;
wire [fgallag_WDTH-1:0]          fgallag_00151_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00151_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00151_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00151_00000;
wire [fgallag_WDTH-1:0]          fgallag_00151_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00151_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00151_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00151_00001;
wire [fgallag_WDTH-1:0]          fgallag_00151_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00151_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00151_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00151_00002;
wire [fgallag_WDTH-1:0]          fgallag_00152_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00152_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00152_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00152_00000;
wire [fgallag_WDTH-1:0]          fgallag_00152_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00152_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00152_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00152_00001;
wire [fgallag_WDTH-1:0]          fgallag_00152_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00152_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00152_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00152_00002;
wire [fgallag_WDTH-1:0]          fgallag_00152_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00152_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00152_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00152_00003;
wire [fgallag_WDTH-1:0]          fgallag_00153_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00153_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00153_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00153_00000;
wire [fgallag_WDTH-1:0]          fgallag_00153_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00153_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00153_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00153_00001;
wire [fgallag_WDTH-1:0]          fgallag_00153_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00153_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00153_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00153_00002;
wire [fgallag_WDTH-1:0]          fgallag_00153_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00153_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00153_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00153_00003;
wire [fgallag_WDTH-1:0]          fgallag_00154_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00154_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00154_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00154_00000;
wire [fgallag_WDTH-1:0]          fgallag_00154_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00154_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00154_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00154_00001;
wire [fgallag_WDTH-1:0]          fgallag_00154_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00154_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00154_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00154_00002;
wire [fgallag_WDTH-1:0]          fgallag_00154_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00154_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00154_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00154_00003;
wire [fgallag_WDTH-1:0]          fgallag_00155_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00155_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00155_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00155_00000;
wire [fgallag_WDTH-1:0]          fgallag_00155_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00155_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00155_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00155_00001;
wire [fgallag_WDTH-1:0]          fgallag_00155_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00155_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00155_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00155_00002;
wire [fgallag_WDTH-1:0]          fgallag_00155_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00155_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00155_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00155_00003;
wire [fgallag_WDTH-1:0]          fgallag_00156_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00156_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00156_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00156_00000;
wire [fgallag_WDTH-1:0]          fgallag_00156_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00156_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00156_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00156_00001;
wire [fgallag_WDTH-1:0]          fgallag_00156_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00156_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00156_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00156_00002;
wire [fgallag_WDTH-1:0]          fgallag_00156_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00156_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00156_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00156_00003;
wire [fgallag_WDTH-1:0]          fgallag_00157_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00157_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00157_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00157_00000;
wire [fgallag_WDTH-1:0]          fgallag_00157_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00157_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00157_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00157_00001;
wire [fgallag_WDTH-1:0]          fgallag_00157_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00157_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00157_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00157_00002;
wire [fgallag_WDTH-1:0]          fgallag_00157_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00157_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00157_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00157_00003;
wire [fgallag_WDTH-1:0]          fgallag_00158_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00158_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00158_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00158_00000;
wire [fgallag_WDTH-1:0]          fgallag_00158_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00158_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00158_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00158_00001;
wire [fgallag_WDTH-1:0]          fgallag_00158_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00158_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00158_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00158_00002;
wire [fgallag_WDTH-1:0]          fgallag_00158_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00158_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00158_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00158_00003;
wire [fgallag_WDTH-1:0]          fgallag_00159_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00159_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00159_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00159_00000;
wire [fgallag_WDTH-1:0]          fgallag_00159_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00159_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00159_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00159_00001;
wire [fgallag_WDTH-1:0]          fgallag_00159_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00159_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00159_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00159_00002;
wire [fgallag_WDTH-1:0]          fgallag_00159_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00159_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00159_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00159_00003;
wire [fgallag_WDTH-1:0]          fgallag_00160_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00160_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00160_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00160_00000;
wire [fgallag_WDTH-1:0]          fgallag_00160_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00160_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00160_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00160_00001;
wire [fgallag_WDTH-1:0]          fgallag_00160_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00160_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00160_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00160_00002;
wire [fgallag_WDTH-1:0]          fgallag_00160_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00160_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00160_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00160_00003;
wire [fgallag_WDTH-1:0]          fgallag_00161_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00161_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00161_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00161_00000;
wire [fgallag_WDTH-1:0]          fgallag_00161_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00161_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00161_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00161_00001;
wire [fgallag_WDTH-1:0]          fgallag_00161_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00161_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00161_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00161_00002;
wire [fgallag_WDTH-1:0]          fgallag_00161_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00161_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00161_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00161_00003;
wire [fgallag_WDTH-1:0]          fgallag_00162_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00162_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00162_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00162_00000;
wire [fgallag_WDTH-1:0]          fgallag_00162_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00162_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00162_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00162_00001;
wire [fgallag_WDTH-1:0]          fgallag_00162_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00162_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00162_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00162_00002;
wire [fgallag_WDTH-1:0]          fgallag_00162_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00162_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00162_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00162_00003;
wire [fgallag_WDTH-1:0]          fgallag_00163_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00163_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00163_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00163_00000;
wire [fgallag_WDTH-1:0]          fgallag_00163_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00163_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00163_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00163_00001;
wire [fgallag_WDTH-1:0]          fgallag_00163_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00163_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00163_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00163_00002;
wire [fgallag_WDTH-1:0]          fgallag_00163_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00163_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00163_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00163_00003;
wire [fgallag_WDTH-1:0]          fgallag_00164_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00164_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00164_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00164_00000;
wire [fgallag_WDTH-1:0]          fgallag_00164_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00164_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00164_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00164_00001;
wire [fgallag_WDTH-1:0]          fgallag_00164_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00164_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00164_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00164_00002;
wire [fgallag_WDTH-1:0]          fgallag_00164_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00164_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00164_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00164_00003;
wire [fgallag_WDTH-1:0]          fgallag_00165_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00165_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00165_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00165_00000;
wire [fgallag_WDTH-1:0]          fgallag_00165_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00165_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00165_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00165_00001;
wire [fgallag_WDTH-1:0]          fgallag_00165_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00165_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00165_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00165_00002;
wire [fgallag_WDTH-1:0]          fgallag_00165_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00165_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00165_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00165_00003;
wire [fgallag_WDTH-1:0]          fgallag_00166_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00166_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00166_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00166_00000;
wire [fgallag_WDTH-1:0]          fgallag_00166_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00166_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00166_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00166_00001;
wire [fgallag_WDTH-1:0]          fgallag_00166_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00166_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00166_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00166_00002;
wire [fgallag_WDTH-1:0]          fgallag_00166_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00166_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00166_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00166_00003;
wire [fgallag_WDTH-1:0]          fgallag_00167_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00167_00000;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00167_00000;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00167_00000;
wire [fgallag_WDTH-1:0]          fgallag_00167_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00167_00001;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00167_00001;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00167_00001;
wire [fgallag_WDTH-1:0]          fgallag_00167_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00167_00002;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00167_00002;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00167_00002;
wire [fgallag_WDTH-1:0]          fgallag_00167_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_full_00167_00003;
wire [MAX_SUM_WDTH_L-1:0]        fgallag_final_00167_00003;
reg  [MAX_SUM_WDTH_L-1:0]        tout_00167_00003;



reg                              I92cb615e2c439914e72ce001256518e4;
wire [MAX_SUM_WDTH_L-1:0]        Iea07d1adf9016a29cffd61d183e268d0;
reg                              Iad799775eb657f8973e6dfcf70a9875c;
wire [MAX_SUM_WDTH_L-1:0]        If92db65b39a83e1c699e4cc6d7f9e57b;
reg                              Ifb064c69c7110c014593149ae69c75fb;
wire [MAX_SUM_WDTH_L-1:0]        I8f2986bc015fcc64ac5e5395ac6dd851;
reg                              I7f7b30f2acbb8e31f50b58096b738254;
wire [MAX_SUM_WDTH_L-1:0]        I355725a804e0df68b4acf96ca98f2448;
reg                              Iefe4099ff7e457f6b9fefc83e176c1a0;
wire [MAX_SUM_WDTH_L-1:0]        I78212ae965ab2dcb2eed0b060d6b253f;
reg                              Icddb43f9b760a4597a0bb637fb405616;
wire [MAX_SUM_WDTH_L-1:0]        I0b56aa7a1b7549c91dddd3a06ecbaacf;
reg                              Ic76e72b434b47c10ebac3fac4ea50bde;
wire [MAX_SUM_WDTH_L-1:0]        I71412803cc5229025487255aec62ec4f;
reg                              I9eb87e62d23bc87d7cd82c0f329f247f;
wire [MAX_SUM_WDTH_L-1:0]        I32fcb28a27356bc6f403528836ea4c1f;
reg                              I2eac5b39c6f485c9ae0bd341f894633d;
wire [MAX_SUM_WDTH_L-1:0]        Iad354d876cb9fc72fc0143e6f7da9357;
reg                              I76992221b1edff5684c482df7ac4693d;
wire [MAX_SUM_WDTH_L-1:0]        If6e745bb85abba7282dae1f6f701225e;
reg                              Iada5bc4a51dc1bf57bb9cca11326bdff;
wire [MAX_SUM_WDTH_L-1:0]        I93bb43c1b89d4c70a57bdc019d64fd22;
reg                              I364ed3f83c49626bc3b939e53524d9c7;
wire [MAX_SUM_WDTH_L-1:0]        I7a2e554d07bbea291f2cfc18694fca3a;
reg                              Ic2b000c3b2ca3beff2d427caab04701a;
wire [MAX_SUM_WDTH_L-1:0]        I3e59b2419c7dd1553b792d536208514e;
reg                              I8e873fb2321eea82bb590a92411e2e2c;
wire [MAX_SUM_WDTH_L-1:0]        I46894c6526983bf1ce4b503159131b41;
reg                              If4cb744ee52b6ae793431cd038069b57;
wire [MAX_SUM_WDTH_L-1:0]        I6404d0df952b5bf8292c753e4c6f35d8;
reg                              I7741e239c16828889d488cc87647c154;
wire [MAX_SUM_WDTH_L-1:0]        I8522c402e654d007abffcb0e904af5e6;
reg                              I7979161aa1e2262ebea862004c387697;
wire [MAX_SUM_WDTH_L-1:0]        I5ed85845c39337c37791f16e718069b4;
reg                              Ic62fc602da3d16fe13d03a49a21269d0;
wire [MAX_SUM_WDTH_L-1:0]        I89013d61c1ea8da8b1c6071cc21c316f;
reg                              I94009bb7239be96243902ab0f0abea7e;
wire [MAX_SUM_WDTH_L-1:0]        I4102100fa5f1dd299af0190862efcc42;
reg                              Iae7b72abf4d3c536330a229e3836b441;
wire [MAX_SUM_WDTH_L-1:0]        I4939f69abb1eac56d5021e06406a93b5;
reg                              Ie5d9cc18b2dd300132470f206452ff17;
wire [MAX_SUM_WDTH_L-1:0]        Iadbd245bf842aebb456417579a3e6296;
reg                              I7c791c854d0bc28e8dd787545f8fbda0;
wire [MAX_SUM_WDTH_L-1:0]        Ifc8ece44a4e68c3117eda9e65f3084d2;
reg                              I5b177dd5c14ad082516b47f550875682;
wire [MAX_SUM_WDTH_L-1:0]        I91679dfab57a372eddc7f9b94a231edb;
reg                              I55e4ad2d71a29ad63b4999d64ac0dc4f;
wire [MAX_SUM_WDTH_L-1:0]        I2213c1a2b831f421707a261f5a58b1b1;
reg                              I59c5da6338f431a626c86a065a355c35;
wire [MAX_SUM_WDTH_L-1:0]        Ic53b875b2ddcba11406eb2ca39354757;
reg                              Ia098bbeda8b755ece6b88eac83d03e55;
wire [MAX_SUM_WDTH_L-1:0]        I634484f00590216c0f74f975c9c83400;
reg                              Ie7470dd75b54d14038de19e4d3043ba9;
wire [MAX_SUM_WDTH_L-1:0]        Ib3b1db2d8b669988c887ed780e439b26;
reg                              Ie95662d4faf6b5a4cd5ecfa41697b983;
wire [MAX_SUM_WDTH_L-1:0]        I735db8b0ee0ec98e4cce0030b11508da;
reg                              Ia1b617e3d141263b51e58c5ef0bd7a89;
wire [MAX_SUM_WDTH_L-1:0]        If1607e907e626902ee26d15020a64c21;
reg                              If9a5d830e3ade0fd96b98f5949f165f0;
wire [MAX_SUM_WDTH_L-1:0]        I081b38dbb37d4c14a6a9fd3fefa13daa;
reg                              Id3de87169c440f95d406693ef77cacd6;
wire [MAX_SUM_WDTH_L-1:0]        Ibac5e7b6d4bf5cd6926358318f0c418f;
reg                              I3751f191f5009322acb7c9be4f8d7129;
wire [MAX_SUM_WDTH_L-1:0]        Iadfc60386481092ae85cc148a2c40abb;
reg                              Ic1927bb3335f6a28c0816eba12d3975e;
wire [MAX_SUM_WDTH_L-1:0]        Ie0ee5445c56a5f9b41640b57422206de;
reg                              Ia659126b51468cfef48c97a135a71500;
wire [MAX_SUM_WDTH_L-1:0]        Ie5f8620371236cb11c9e88c16b509ee8;
reg                              I3c3c22bf63e55a81ae91b1dd1ef615a0;
wire [MAX_SUM_WDTH_L-1:0]        I8d7c1fe2e33bbd45379b0325a3c5e989;
reg                              Ia62832d325f86160285c4d1a790a32cb;
wire [MAX_SUM_WDTH_L-1:0]        I4fbdc4ee57a3be42b62d9bd43078d6ef;
reg                              I83c7d177eec2dad0a924557cdc91ba77;
wire [MAX_SUM_WDTH_L-1:0]        I5510b88bfd65811b3200adf4ef975b48;
reg                              I7050adb9d06f767549b7f35c4679e391;
wire [MAX_SUM_WDTH_L-1:0]        Ib57ef2f577cca54713c16717cbbd1ce9;
reg                              I04aacd95d9e44657f616e01c9053f0fb;
wire [MAX_SUM_WDTH_L-1:0]        I15943aa74e9fbbaebdc0d54eb6a3bffa;
reg                              I2ff317d57f59747c4524ef4278d51092;
wire [MAX_SUM_WDTH_L-1:0]        I6ac24c46319a787daa5c545de8c6eeea;
reg                              I8bd2a9d90074500698b302cb8db7f03a;
wire [MAX_SUM_WDTH_L-1:0]        I52403a0454e5fa002e79eaab7ea497bd;
reg                              I3b8cdfb1440732ce98cd1676e05a2af1;
wire [MAX_SUM_WDTH_L-1:0]        I634f0ce28934600a1a31ab0d8e59b4a9;
reg                              I671de3d408b5b783541663c7f1e3a6fa;
wire [MAX_SUM_WDTH_L-1:0]        I7103aa739616a39c03e675ea0efb0335;
reg                              I446857735e680cae93a24dccb59b1924;
wire [MAX_SUM_WDTH_L-1:0]        I0296d01fd3f9a269a617efd4beea9b8b;
reg                              I77b05a8aa92c66a235195a66dc13c0cc;
wire [MAX_SUM_WDTH_L-1:0]        I065a81ba25962785215583e7ece27661;
reg                              Ie92110d19f4886cdfcfacd0920c06a4e;
wire [MAX_SUM_WDTH_L-1:0]        I631a3300cb6685f47da7781940ec5d27;
reg                              I36ba87b69b5b9dd919319230f697dfad;
wire [MAX_SUM_WDTH_L-1:0]        I8bbe1a2ace8f51aa22cca5d9fc66f136;
reg                              Id20e72ac258d1d1b6cdca1e6c9e3596d;
wire [MAX_SUM_WDTH_L-1:0]        I38c3e3e136acb79c8a0ff850bcc55f16;
reg                              Ifc34f5d6b7a7d0533439794958959856;
wire [MAX_SUM_WDTH_L-1:0]        I35b2c7e9cdc53a98913e1c16a3a47b37;
reg                              I849ee5d34760be03d4285185136aa52e;
wire [MAX_SUM_WDTH_L-1:0]        Ib1a2b31d49ae476e2f1fb9acba2d5af0;
reg                              Ia3559d98eb372b7307f30ad1f7c4c7cd;
wire [MAX_SUM_WDTH_L-1:0]        Ic72f41f9bbf470aee3c9b9b8787b31c3;
reg                              I7332e088bbff69db19c62685e033d26a;
wire [MAX_SUM_WDTH_L-1:0]        I3ea4c33a9419820ed54460eb64134dff;
reg                              I44daa5992b00e7af19adbee70bf01f2b;
wire [MAX_SUM_WDTH_L-1:0]        Ia0d940e16c8cbd4f7544f5a5cd7d83b2;
reg                              Ie517386cb5832e406fefc5e85eb2e7d1;
wire [MAX_SUM_WDTH_L-1:0]        I4a8abfa0896ce414d9b98093ef84455f;
reg                              I9b096ce09467c10f448496fda13987d2;
wire [MAX_SUM_WDTH_L-1:0]        I680be647bf2a62e0ee9b5d379dc87b4f;
reg                              If1c0a3726041f70e508d68cbf6e40e04;
wire [MAX_SUM_WDTH_L-1:0]        If4d75f83299a21802b6fbe136913489f;
reg                              Iaf36ce8598a29573979c683a5e2cf9fd;
wire [MAX_SUM_WDTH_L-1:0]        Ibddfda6413e3dd2f483c3174ea836b6a;
reg                              Ice82cfe55a5f226746e59e5c8beb46be;
wire [MAX_SUM_WDTH_L-1:0]        I33bddb0adcc2af7b12a83bf843036385;
reg                              Iea1297491d1dfe98f395d8c73808a893;
wire [MAX_SUM_WDTH_L-1:0]        I529f92b82248efe2cf64f7da0ec8283c;
reg                              If43dd31198c8a0da6fabd194cf13bb70;
wire [MAX_SUM_WDTH_L-1:0]        I2f34af0036985cd94ade9cc905bec065;
reg                              Ibeb8c72b90b50c6897224ca1a792fa56;
wire [MAX_SUM_WDTH_L-1:0]        Ia1a0d8d7dfd6e877f15cce773f85f5b7;
reg                              I8e87530a131b5a73cad6df68b9e4967f;
wire [MAX_SUM_WDTH_L-1:0]        I5dd29fd1a73df5662d2b636e7285bad9;
reg                              Idf8d15c7bd7705b9aafbda09c3a5b46c;
wire [MAX_SUM_WDTH_L-1:0]        Ide530e6f4622c8a7b101b6dce9650e42;
reg                              I2aea17846a53e2eb2968581ee2c48226;
wire [MAX_SUM_WDTH_L-1:0]        Ibaf00a6780325882067a79f0c4d693d2;
reg                              I169d8f2bb5fde5b202b4239b7a7f1ed5;
wire [MAX_SUM_WDTH_L-1:0]        I16e3559c63ebfed83d6698fc9a9cd93a;
reg                              I40a223380fb4414a3f26a08cb90025ec;
wire [MAX_SUM_WDTH_L-1:0]        I9747a02384abb1c2dd1f52b3a5a999cc;
reg                              Ie117f6ec475f5d6444998af151ce4e69;
wire [MAX_SUM_WDTH_L-1:0]        Iceb7a1d4c23806b8f5824016779ad129;
reg                              If7f3174da35dd39af7f4792aaa649bf1;
wire [MAX_SUM_WDTH_L-1:0]        I40ef50004a60ae58aedc49eb5e6797c9;
reg                              I719a892ad54e63b217c7271741b29cc5;
wire [MAX_SUM_WDTH_L-1:0]        I753f92da60980736440aba814a156f1e;
reg                              I4acf6d84471cd237f65c9b2391b7a20c;
wire [MAX_SUM_WDTH_L-1:0]        I4ac79b67a8904b95f7912d24af420585;
reg                              I7a387a1f887c32e9d0f8e89912a8618c;
wire [MAX_SUM_WDTH_L-1:0]        Iad44c932cfa5c249c5e59f8c706173a8;
reg                              Ib862ac63c230ccde7fae0e62f9d047fe;
wire [MAX_SUM_WDTH_L-1:0]        I10f14b6433498e3b9e9bf021b60115e8;
reg                              I8f1a8a22637d37c3692e808d5eb3d543;
wire [MAX_SUM_WDTH_L-1:0]        I96008f47b9f134c9c4274cfcfb28e550;
reg                              I6f420c64640dfb0c001f57df7e3b4504;
wire [MAX_SUM_WDTH_L-1:0]        Id0344146d1a53d418add6d2b185377dd;
reg                              I3600031716c2b4e21c9f577d34e033dc;
wire [MAX_SUM_WDTH_L-1:0]        I1eede74f12d37331b399eb7136bc621f;
reg                              I002820a37fa7c6c504c487df4368e2cf;
wire [MAX_SUM_WDTH_L-1:0]        I3e4754acc31d99bc71525789bdee0c1a;
reg                              I8a4c1f23212ff846400651b100add502;
wire [MAX_SUM_WDTH_L-1:0]        I11c1fc94a3bd6dffa17e1571cc6ae97c;
reg                              Ice1ce5b4c30841dd92268559ebadafcf;
wire [MAX_SUM_WDTH_L-1:0]        I5395ee57418c31e11cf847f0f514ec19;
reg                              I3eeeb1949945032d6c1759875426b733;
wire [MAX_SUM_WDTH_L-1:0]        Iff125392fa39afebae1637a19c4e23ec;
reg                              I384d5377ee6b8f7eb2db23a2e444ddbc;
wire [MAX_SUM_WDTH_L-1:0]        Ia6308e16fae5428f4ab6560f5b21479a;
reg                              I30d615203b697787ead37394953925cc;
wire [MAX_SUM_WDTH_L-1:0]        I5ea02b5349cd4d99ccbcb6b26f0cfdd7;
reg                              Ib16548d471f0a4f4625852ea04335dcc;
wire [MAX_SUM_WDTH_L-1:0]        I21de4f6194dec9e3c401934db92c25e7;
reg                              I0987c561670b7b2b6683303c1be39561;
wire [MAX_SUM_WDTH_L-1:0]        I57d0920119f8901bd4dea2d5f8fb5d90;
reg                              I2bdf4736022e5da7294a0e851006a124;
wire [MAX_SUM_WDTH_L-1:0]        I89537301987d6da0dbe6cff3caab3ff4;
reg                              Ic6fd9592d2ffcb8f4ca83c6f0bd19975;
wire [MAX_SUM_WDTH_L-1:0]        Iaf0bbbe791bb71d0f557dc71caa5fb87;
reg                              I14bf11ad80890227e47fda26ae1b9c24;
wire [MAX_SUM_WDTH_L-1:0]        Ic7ff9cde71054c1ee9eef81eabdd7061;
reg                              I8ca17b6cf35e1b1f8f601604575d3f27;
wire [MAX_SUM_WDTH_L-1:0]        I88c10c47ae424fbdcb852fbf1e94127c;
reg                              I275cd09649a750edb8ae8313e4e1e279;
wire [MAX_SUM_WDTH_L-1:0]        Icd2e75e47cab1d539ba9ff1b6e1d7155;
reg                              I7d6a6026eb3c4d06e682523424f9628f;
wire [MAX_SUM_WDTH_L-1:0]        I37e6bc7aff363ed0ed1f84b23c5f3e34;
reg                              Ia0c192e590d8c914555b434ce5a634a8;
wire [MAX_SUM_WDTH_L-1:0]        I733605337bf6972630c089d32fd7f98f;
reg                              Ic98c8641d2022080297c54ff2539e75d;
wire [MAX_SUM_WDTH_L-1:0]        Idcb1d8bbdeaed6768c2a418c3048e6ee;
reg                              I87f34821cd0b58f8855b25c75f2dd32d;
wire [MAX_SUM_WDTH_L-1:0]        Ia89da2f1890524ad3519ab403dd0686c;
reg                              I87211ac14d832ad3205d47fb83cf256a;
wire [MAX_SUM_WDTH_L-1:0]        Ie33a780b0221084898c9fc5b237b244a;
reg                              Ib81431cfb3b281555fa7e5b4582a2524;
wire [MAX_SUM_WDTH_L-1:0]        Iabbd1668e0014df518ede5216232834c;
reg                              I835b902949c2c4c09b757d4d35574a76;
wire [MAX_SUM_WDTH_L-1:0]        Ibd89458312687610aa166a9538968851;
reg                              I8510240df7dc41f85ad58a39868a1fd7;
wire [MAX_SUM_WDTH_L-1:0]        Icbaf92a8e9875bcb19a1d074779a9ea5;
reg                              I1b6abc8fbab3849b285e9f88a4fe867b;
wire [MAX_SUM_WDTH_L-1:0]        I80f3c8559da8e97bc5397bb8b621a0bd;
reg                              Ied638fee34f8baed4154b0b72e43a21e;
wire [MAX_SUM_WDTH_L-1:0]        I7a0eada108891aba06cecab5071232c9;
reg                              I14fa7aebb608d4a3d67176ba27d34d9a;
wire [MAX_SUM_WDTH_L-1:0]        Ie21a2c9b22e7bf8425fb5c0f33e5f4f7;
reg                              Iad90879acba3fc2101829549264960f3;
wire [MAX_SUM_WDTH_L-1:0]        Iaa5b2807e5cc2403c5787eeb3d10ca6b;
reg                              Ife0952b85f14a960007b67646b0cd969;
wire [MAX_SUM_WDTH_L-1:0]        I6da2b3a481ee71b85f3087b36b399288;
reg                              If876ca6a14ffb4323503ed46666bc25f;
wire [MAX_SUM_WDTH_L-1:0]        I11094e852295755925c3c61f1df81643;
reg                              If2dfcbf493b761fb5d7c622e739b23f3;
wire [MAX_SUM_WDTH_L-1:0]        I9c633aa620cca127b0ff8cf882178e76;
reg                              I2c8f4a147b363d9c5ef0e080d9a9ed40;
wire [MAX_SUM_WDTH_L-1:0]        I694d471fd353eb54aae08a2afa7b645a;
reg                              I485f9d1104a965d5d035feef912a2ca8;
wire [MAX_SUM_WDTH_L-1:0]        I816704585ad393f685731104ad3ec64f;
reg                              I10fca5f2cbf5e2bc3433c0dda579a051;
wire [MAX_SUM_WDTH_L-1:0]        I85d95015a9ce27a18ccbf73bbbcdbd70;
reg                              If8572800d5d80cc92dd917b60447b63b;
wire [MAX_SUM_WDTH_L-1:0]        I992e7c551b4aa818606c3465d33eb798;
reg                              I24645082ef16129eed1c574f5fc601ca;
wire [MAX_SUM_WDTH_L-1:0]        I2ead0e9941e2280309ab53535b1e1ac1;
reg                              I207a0f6184a0b3be71766a8b47ea5535;
wire [MAX_SUM_WDTH_L-1:0]        I56873feb8418005b5661c7382f2dbeec;
reg                              I5cac08dabbb6de3b01c821d4db93a8e3;
wire [MAX_SUM_WDTH_L-1:0]        Ib6ea4a822da2ea32e0abf6cf8a33d295;
reg                              Ibe6b8c57d7ff47b6fdad5fadf1f6b841;
wire [MAX_SUM_WDTH_L-1:0]        Id1659ccdeaea3e59eb2d3f65a65ebd05;
reg                              I477326720157df2503149125a43ee987;
wire [MAX_SUM_WDTH_L-1:0]        Ic2171967791a0329f3e39fc19d0a6bc8;
reg                              I2c741a5fed7d88e9bdd6b7459feac649;
wire [MAX_SUM_WDTH_L-1:0]        I7d5041a6796c00188f74936d283defe6;
reg                              I17a6511072c7fb4846be5844decf17d6;
wire [MAX_SUM_WDTH_L-1:0]        Iba7608ee0a01af103e022bcaf564bf6b;
reg                              I5ebc3047985651f4b9a957d502a97e95;
wire [MAX_SUM_WDTH_L-1:0]        Iedbe9d0e48bd36064f59faea51afddb9;
reg                              Ifa09fc1b009d073d5a9973b430c63469;
wire [MAX_SUM_WDTH_L-1:0]        Ic3871325d57b310c95ca02fcaca529eb;
reg                              Ie6212a29c7c6b035cfff4c869f945b68;
wire [MAX_SUM_WDTH_L-1:0]        I42f9b1f8ef24ad56c10086852678b456;
reg                              If343015b4815b01dae88bbb6f2017b3d;
wire [MAX_SUM_WDTH_L-1:0]        I3ed5d0fca86f35b3d4b4a89c6147d0cd;
reg                              Ia0116a3cebf94318ed5b287960957ad6;
wire [MAX_SUM_WDTH_L-1:0]        Ib0126fb335e32793c400a97c5a4a337c;
reg                              Id75c23e80cdf25d883806ed20d4ae783;
wire [MAX_SUM_WDTH_L-1:0]        I20590d8fb97ec0b2164ffe17826136a7;
reg                              I1b43f29e0ddb72467befd6f3a9c1c829;
wire [MAX_SUM_WDTH_L-1:0]        I3c128efc9f80c9b8334bf7b61de71b43;
reg                              I3fd0fa3b774d30a267d61e9427d09f3f;
wire [MAX_SUM_WDTH_L-1:0]        Ic7147944f8835e26b9838fdbdc18ca41;
reg                              I2eb08ebaa07a1004638cdd61a7209b7d;
wire [MAX_SUM_WDTH_L-1:0]        I698b1dbc9d8664d1c86c7a763d97b3b7;
reg                              I258c45897919cec5c6acaddee7f3a41b;
wire [MAX_SUM_WDTH_L-1:0]        I508bbade361787127e1a2e8687ec884c;
reg                              Ib42d37576e3aff3d205f1f8822cc58b5;
wire [MAX_SUM_WDTH_L-1:0]        I2afeb2a7b199c0c6738938f156ae4274;
reg                              I1c2ee281cd47a8414851c5e1c758ea65;
wire [MAX_SUM_WDTH_L-1:0]        I86255756ddd1f88b74e070b19f8c3bfa;
reg                              Ie644d131c4f2c603e8e64c5581fdf822;
wire [MAX_SUM_WDTH_L-1:0]        I7d4924388dc5373ad7936dca76797473;
reg                              I9b76f0121a3f7e887e7121db50024ab4;
wire [MAX_SUM_WDTH_L-1:0]        Ie317e5ea2ca4ba2060d0f491290af96f;
reg                              I9eaf4e9ebe07717503ff69b51f0e1905;
wire [MAX_SUM_WDTH_L-1:0]        I56ea52c50a188ec47e48740839a031c9;
reg                              Icb0841ecf142687c3aa23e68f01c927c;
wire [MAX_SUM_WDTH_L-1:0]        Id9b9a8fe43992ec0793845715dd2226c;
reg                              Ie8c0fac00a9de74870e59cbf9e87a39b;
wire [MAX_SUM_WDTH_L-1:0]        I93b69bfb228db4b569a6772179d603be;
reg                              Iae5d6faac1f5685cb1d400ee2b1d85e0;
wire [MAX_SUM_WDTH_L-1:0]        I71afab29cdb962e1f1ca21b61dfb50c6;
reg                              Ib62b02ddf0f57bee49838d19783ef6c3;
wire [MAX_SUM_WDTH_L-1:0]        I9905e2686b350e8a6e7f790563a91294;
reg                              Ibd59d0e5a062f149bd0e91ba76985a13;
wire [MAX_SUM_WDTH_L-1:0]        I524e78ae6a4204e17ba4532dba047d4b;
reg                              I876fdba97e755b74532f7ab191fbac14;
wire [MAX_SUM_WDTH_L-1:0]        I71228fe4188ab1d9796081184a422094;
reg                              I8edf1a08ef943f06ee28771c6e140e28;
wire [MAX_SUM_WDTH_L-1:0]        Ie19b39200436b0bfca13502ad36c21b9;
reg                              I7e12ad8a8ef857e02f4563b2f3a7f0ca;
wire [MAX_SUM_WDTH_L-1:0]        If6657f90c84ca5e2ba08ec705f34be03;
reg                              I17b3a9df6752da6cc987e902e6bbad48;
wire [MAX_SUM_WDTH_L-1:0]        I60ec7459bbe99fce295406bee1f2af46;
reg                              I487496233a32f657171b3789590d0522;
wire [MAX_SUM_WDTH_L-1:0]        I29ab844f80c105d247c5c15faa35863c;
reg                              Ie34534dfd435b3d1cf35e82ca71e83ba;
wire [MAX_SUM_WDTH_L-1:0]        I856fa68463aa5ef1ae53442699d38b33;
reg                              I0e8679271ba733bb87c44b6b9f0b6ed2;
wire [MAX_SUM_WDTH_L-1:0]        Ic3d00a27f15f8983a120395082854d6b;
reg                              Ic14760b65c6fe150c3c48e64389a41d8;
wire [MAX_SUM_WDTH_L-1:0]        I6b1d01c3cb8fb51e43cdb788b89816be;
reg                              Ied6c684cdd280b41ffab93a026d27282;
wire [MAX_SUM_WDTH_L-1:0]        Ib74a56900c1f8b159ad381f61acee801;
reg                              Id0f4dbb72da33748d8baf723c5a32567;
wire [MAX_SUM_WDTH_L-1:0]        Ia5eba52d169755c507b9e0094e467fab;
reg                              Ib0bb71b1f8829347b3a9a7543f9dd964;
wire [MAX_SUM_WDTH_L-1:0]        I0899e8fec1a7209cd94757c0b2f87c9a;
reg                              I47cbb92d2284aef7b9e56e88f0ba6f7e;
wire [MAX_SUM_WDTH_L-1:0]        I08ece7cd684e593e02321612b7a88cee;
reg                              Ic69094123b75ae36e3e54f179a9f2cb5;
wire [MAX_SUM_WDTH_L-1:0]        I691c84d81c60a462e28e2b2bae3ea845;
reg                              I07abbbd75d91018ac53f53e64cffafb9;
wire [MAX_SUM_WDTH_L-1:0]        I58dc9cce6384160c0a85c6efb3319cdb;
reg                              Ib02268d5048c7c8e83118070e927453f;
wire [MAX_SUM_WDTH_L-1:0]        I56bf74b5890ec67090f499afdc0a9c88;
reg                              Idc2a9c6dd8d2aa912548c918c8a488f4;
wire [MAX_SUM_WDTH_L-1:0]        Ibaf2f1f8bda2f6b932dc30f8369c0e1f;
reg                              I5ad7eb9d3ce7c712515254f892d1670d;
wire [MAX_SUM_WDTH_L-1:0]        Id9364a29fd79b52d0442e18dc0227854;
reg                              Ife25829fb3c5023b7d69bbaadf9cf77e;
wire [MAX_SUM_WDTH_L-1:0]        Ica3a41ace27f7d94377981079952f4f7;
reg                              I8b2a79aa4ac88e6b4ca8188a7852022e;
wire [MAX_SUM_WDTH_L-1:0]        Ib57795a63d642a73456324bab41384b6;
reg                              I081e2595b18f306a74d070203447ecf6;
wire [MAX_SUM_WDTH_L-1:0]        Iabf572c97b48c6a7dcc19e56676e3a82;
reg                              I68b152a599887c0039dd9d45c528c219;
wire [MAX_SUM_WDTH_L-1:0]        Iefd370d0df1a93639af482f78a1e8706;
reg                              Id051f1d5454802e0eb37e22248efe8ca;
wire [MAX_SUM_WDTH_L-1:0]        I995d2809ffaf0ecda6a004d01cb9c8c4;
reg                              Ic4c6f707f461cebbc4c93f2ba664ae7b;
wire [MAX_SUM_WDTH_L-1:0]        I4e8ebc46bc068c3f9889d970db131112;
reg                              Ia538dadbd6ae3711740595a18c89b65d;
wire [MAX_SUM_WDTH_L-1:0]        I7b561638da1b4a45ff59be81243e4471;
reg                              Ie7d9730b191781c78391141d95d4f8bd;
wire [MAX_SUM_WDTH_L-1:0]        If0a3b88a66a816b25f17ced5d0e8f775;
reg                              I12f2f886517647044cc251861721bbb9;
wire [MAX_SUM_WDTH_L-1:0]        I0374ada4fe50717f2158468b7ad205d4;
reg                              I615053b36a1851a06125e2ed5ec7f880;
wire [MAX_SUM_WDTH_L-1:0]        I357137b41bb91e0659b1ac6ead9b5c12;
reg                              Ifbc6aa14cd448bbe416897a3671ba857;
wire [MAX_SUM_WDTH_L-1:0]        I5d70bc64cf7b3d3ef4180e082e533237;
reg                              Ie596289582a73e37f78f4ca4cab21e3c;
wire [MAX_SUM_WDTH_L-1:0]        I7d9ad929660cd212387d893266b681da;
reg                              Ifad8c7bacf72583f91be27fbe5b7a1e1;
wire [MAX_SUM_WDTH_L-1:0]        I34be4b353cf75603301372840c2f91c2;
reg                              Ie74c72742807ae4243748fd27d80d626;
wire [MAX_SUM_WDTH_L-1:0]        I14834fc8e6489775359bcecf5a37ff4d;
reg                              Ie7a68c2b368a295f95571bc4a109b9f1;
wire [MAX_SUM_WDTH_L-1:0]        I633a74e4dfa841c9fd13dbb6564c8493;
reg                              Id88a7edf897eea1b4a137141789a04f5;
wire [MAX_SUM_WDTH_L-1:0]        I157bd468200e63385583b9045758d81e;
reg                              Ib13436ad16a37d656d6b1ee95b9aee20;
wire [MAX_SUM_WDTH_L-1:0]        I918c46173eebc5b2a95e041cfd91d958;
reg                              Idc07dc30c0a957e474546ac7a60df38f;
wire [MAX_SUM_WDTH_L-1:0]        I4f8792c18bd07b23e82bbc44b4ca947f;
reg                              I595665d8128bb87ab62741d7ac520a4b;
wire [MAX_SUM_WDTH_L-1:0]        I8d0a1ae4c47edf1f2b99d1175aaa7197;
reg                              I256050251d23250854ff337bef28e460;
wire [MAX_SUM_WDTH_L-1:0]        I734e601f5f9d568a44a48834559e04db;
reg                              I82f0e5a32d1bcd761a74f1f9ce8c88ba;
wire [MAX_SUM_WDTH_L-1:0]        Ie421da1dc5aaea57c50d0c7d9c5a2717;
reg                              I98febac90cccb5fc1f3d966b6e38c4d3;
wire [MAX_SUM_WDTH_L-1:0]        Ief5cbddfbfb98fce4812a676849b9a98;
reg                              Ib534288c2cf976b6ec85db743bc2a823;
wire [MAX_SUM_WDTH_L-1:0]        Id113cab2dd1949d32e3c1c15273185c8;
reg                              If988b82b86db1f4ff6d3695f7b0197e4;
wire [MAX_SUM_WDTH_L-1:0]        Icfe1a689e33b2b9aa9dba692d6d610b9;
reg                              I6ef260ef75e47b011a46ba2080ac3684;
wire [MAX_SUM_WDTH_L-1:0]        Ia4b671f3360f3ce55db0dc0e4d78ddbe;
reg                              Ifc1da524e7670772834d521a6fc4c96f;
wire [MAX_SUM_WDTH_L-1:0]        I60cbd4369e7ba9b6532f279e5c59084c;
reg                              I852d5295a32984af00c95f6d9389555e;
wire [MAX_SUM_WDTH_L-1:0]        Ifb6c65a00d9a2c31d8b1119b949828d8;
reg                              I3c0a621dbef864fd1f566bc2e47f32c6;
wire [MAX_SUM_WDTH_L-1:0]        I4a777f0dd62b19dd340ad31517c4e789;
reg                              Ic04828ba2db8239b093043c27476d345;
wire [MAX_SUM_WDTH_L-1:0]        Ib75747cb32130d44b338ed8c8af8ca11;
reg                              I319012bc6fe93d78de57bcace0caaef5;
wire [MAX_SUM_WDTH_L-1:0]        Ic7e35cf8d5cd230b94c40714f16e2418;
reg                              Ibb35bace971548c9fc98d773d1aff712;
wire [MAX_SUM_WDTH_L-1:0]        Ic51bb9184dfd103703cd0c6ad6edff4b;
reg                              I90023493600924a76d2192080cf6194e;
wire [MAX_SUM_WDTH_L-1:0]        I103f1449c78c47396d6a54dc1c810934;
reg                              Ia9f5ce4603af279bbd9b486b67016482;
wire [MAX_SUM_WDTH_L-1:0]        I56b3a97dc3037f0bb2eed93a9482c813;
reg                              I05721e06a1acdcc0571907c7d853f18c;
wire [MAX_SUM_WDTH_L-1:0]        I51e98035b35a35fdc52f5bab8f19c152;
reg                              Ibfcfd3151af0d82bfce293ada44059b3;
wire [MAX_SUM_WDTH_L-1:0]        Ia6a7f9beaceb08d81012f0e72171252f;
reg                              I9539fcc40d26b13015a864718b116d5b;
wire [MAX_SUM_WDTH_L-1:0]        I21b062856ced09cb9131c01b5e166f32;
reg                              I5490039998187a1a2efc3549e3dee7d6;
wire [MAX_SUM_WDTH_L-1:0]        I4f1221ce7880729fe584b42ef3afe6b2;
reg                              I2b97a79c90f6578c8b2f321f8d598cc8;
wire [MAX_SUM_WDTH_L-1:0]        Ie7f3f1d6cee7f02ae1b17740ed54c049;
reg                              I0c616f736879c28a5222de3d6f49a587;
wire [MAX_SUM_WDTH_L-1:0]        Ib196f5bcf9152703dc32c5101076600a;
reg                              I5590d801fd7fb496019d4c31b7c6d898;
wire [MAX_SUM_WDTH_L-1:0]        Ide9ef5a16d8fe32353c2c2a30e8ee3b0;
reg                              I27e1d2e0e980216b27b90ea48c061025;
wire [MAX_SUM_WDTH_L-1:0]        Iee6f2484a381bd42e441ff072ec582e4;
reg                              I474f6bd977f4197742d0bddb3bece684;
wire [MAX_SUM_WDTH_L-1:0]        I53121a39de0bcba91a4d0438be2ae958;
reg                              Iaa1e981134f5a5c02983c49562683bc5;
wire [MAX_SUM_WDTH_L-1:0]        Iff7950f24f0a6b0073942c37fff49d37;
reg                              Ib051eb1091a85f85a1e50007f1b27cab;
wire [MAX_SUM_WDTH_L-1:0]        Ide86f019e9573706c25bd8b4552396a8;
reg                              I6b5645cdde4b35a16fe3e91d90caaa4e;
wire [MAX_SUM_WDTH_L-1:0]        I2370042234b0e93bb66e44b97fca3e43;
reg                              I8850ab26807dcd55fefadf6310729ca7;
wire [MAX_SUM_WDTH_L-1:0]        If9efe7a1c359ec03014a52870ac13aec;
reg                              Ic5cb81c821716a8aabf8cc2283ff73ba;
wire [MAX_SUM_WDTH_L-1:0]        I6a6eb62960b616043415406ebfc21346;
reg                              I9a6923c6368526a53ef70e16471386ef;
wire [MAX_SUM_WDTH_L-1:0]        I06c7728ef64be8311f48d10d766d0c44;
reg                              I620b8ecdcaccc1ec80ebcf9fa6af0017;
wire [MAX_SUM_WDTH_L-1:0]        I9fe11f6c8147391aa4a5afd1a4e4f731;
reg                              I141cda06bae0c5666e3bc61c6fe5ad66;
wire [MAX_SUM_WDTH_L-1:0]        Id50edc56fce48130247fdbc42eeff9ea;
reg                              Ia9c273b32d0701c7f185ab2de9e57829;
wire [MAX_SUM_WDTH_L-1:0]        If3e5161254eb9056914c46263b865c10;
reg                              Ic3fb524ab434e80b3289c9241b65d224;
wire [MAX_SUM_WDTH_L-1:0]        I58703e8b6d04f8c69ac38f5fcfdc4efc;
reg                              I23c8b64e433af0bd00cef44e38df99f8;
wire [MAX_SUM_WDTH_L-1:0]        Ie1f41720e296ced1b74cb325b666d88f;
reg                              If6a5dc79c0f6ce348956286737a369d8;
wire [MAX_SUM_WDTH_L-1:0]        I5d5701435c96f1078e741921b56e3c65;
reg                              I34e6e9d2153e4a70ee36ab85e72d5318;
wire [MAX_SUM_WDTH_L-1:0]        Id96e744d9b10dcddd1ae0115ea57a76a;
reg                              Ifdabf743a8cb46b7053000ff48ea0c60;
wire [MAX_SUM_WDTH_L-1:0]        I0c0060fe260afa3cdc72f35ffb6938ff;
reg                              I22f5bb821a2571d1764978fd76c8f1d0;
wire [MAX_SUM_WDTH_L-1:0]        Iaec1f186cb4a65da21d41e637fc628f7;
reg                              I1b695aa715615662eff7065c742b0859;
wire [MAX_SUM_WDTH_L-1:0]        I9c15a6a5c0db11ede80ff6d04c9a56d8;
reg                              Iec91b3ca3b54010755d57f8b8ea4a544;
wire [MAX_SUM_WDTH_L-1:0]        I8922487573e02d684a3d71448c3828f5;
reg                              I06ad520cb02e46d34c45f207d42a9243;
wire [MAX_SUM_WDTH_L-1:0]        I47f17afcd5871fc3ac378316fd3d7ae9;
reg                              I9d18ff3465afd8cae63abba68487542e;
wire [MAX_SUM_WDTH_L-1:0]        Ia9642d79bb50567348083b4435c7d66d;
reg                              I914dedc1d5e5e21c9b8d07ec0ecc01f9;
wire [MAX_SUM_WDTH_L-1:0]        I2b2bd845428c49346ef8e94e95b618f8;
reg                              I3375fff5ee0d4b4b12c5a70fbdee59fe;
wire [MAX_SUM_WDTH_L-1:0]        Ib730fdb59198f23d1e590f6d6039e96a;
reg                              Ia8e304ca12c82e41cb8e4de7be199394;
wire [MAX_SUM_WDTH_L-1:0]        I644e83f0a7d432fba38ffb2d99088eca;
reg                              I3566f2779e860008b1a5d305366a07c9;
wire [MAX_SUM_WDTH_L-1:0]        I97f2b15ce0a74e68d5a4438111adcb0a;
reg                              Ie68b31360c12a83c6095254b6f14603c;
wire [MAX_SUM_WDTH_L-1:0]        I84c88b631bed5311cb6e99e58941149e;
reg                              I42ae0c42360c977b35429ce290516a6f;
wire [MAX_SUM_WDTH_L-1:0]        I45c5e6710240685bf54b73b0d7a64271;
reg                              Ibe01835305315fab50269c72ef849b61;
wire [MAX_SUM_WDTH_L-1:0]        I5827bc87b5db1801b7db16e1e61515db;
reg                              Id806a2df1c4519bbbe811791cb4072f9;
wire [MAX_SUM_WDTH_L-1:0]        I1c85c8f73ef80a6808c6aec0c8eca8ab;
reg                              Ifb70a30f8bade95f402e71f95fe6644b;
wire [MAX_SUM_WDTH_L-1:0]        Id13c99b7f7500c8195b54627efbc4232;
reg                              I592a495aecc800236c3470ff8e6adbb5;
wire [MAX_SUM_WDTH_L-1:0]        I4636821315d702a677dc93113872e647;
reg                              I1c8024aa9d81704d2dcf63e34853f8cf;
wire [MAX_SUM_WDTH_L-1:0]        I9c981b0614a29386ca5e8ebc06a17f15;
reg                              Ief03713f5cf37200373a20d42c7fc9eb;
wire [MAX_SUM_WDTH_L-1:0]        I4df3d4dac24877b14e6d361bafc1a800;
reg                              Ic3cb34aae74c5f1a870b3635f8a40764;
wire [MAX_SUM_WDTH_L-1:0]        I913d818403024510c55b65b56a38dd89;
reg                              Ifa3df8b249467cc1e827c69925ef415f;
wire [MAX_SUM_WDTH_L-1:0]        I57015930f5b09a6c6b030ed01dad2177;
reg                              Icf3ad912aaeaa0c5cd1ab0edb898d6e8;
wire [MAX_SUM_WDTH_L-1:0]        Ib54d55a70605119e37e9898b940ff636;
reg                              Ib774f380e3d7cfd1f5f064e93d8134b4;
wire [MAX_SUM_WDTH_L-1:0]        If7e146da4f3bd255b8457fd6902005f6;
reg                              Ic07c650e6e49892a41cfaf3a37471426;
wire [MAX_SUM_WDTH_L-1:0]        Ied00d87af99ae55144fdde41ebfc1357;
reg                              Ib1073489d63ea33d7f3892f4ff875358;
wire [MAX_SUM_WDTH_L-1:0]        I7774313f1ae5a2de98855aad572b3676;
reg                              I174b6c36f2af82f8047cc76543a3b4ee;
wire [MAX_SUM_WDTH_L-1:0]        I679baea452c3c6d04c53baa88edd8eb3;
reg                              I953b975a89adcc88039284970e9b3404;
wire [MAX_SUM_WDTH_L-1:0]        If4132b39ddb92aa02d8d0346fb0e6691;
reg                              If2b40d249c531e10cc22d1335f350441;
wire [MAX_SUM_WDTH_L-1:0]        Iba70e737d52e6812a67c159520e5192f;
reg                              I44ccc3ae897109dd51f9afeef93daca4;
wire [MAX_SUM_WDTH_L-1:0]        Ib9ceb8315f0cd848f861bab677c2c694;
reg                              Ie9236599cea94cfb603c6b977fdbb44a;
wire [MAX_SUM_WDTH_L-1:0]        I7846bc2cc11e08d05f7c853c4920d555;
reg                              I25f1ee9cee4d04bd8fec1fe601d016d7;
wire [MAX_SUM_WDTH_L-1:0]        I0865623d3350645e63fa6e6c9b78ac57;
reg                              I5ec1e530b9007a75a778af4d82ab427b;
wire [MAX_SUM_WDTH_L-1:0]        I0262b30a4efa9f1cfb11d1c3940de9e7;
reg                              I8a9e516aa824260998d10db758642bb0;
wire [MAX_SUM_WDTH_L-1:0]        I7a2e79d42779ad235bca6ce3757cf588;
reg                              I70dd1350d65155ee7b562f4c79024a3d;
wire [MAX_SUM_WDTH_L-1:0]        I09e9a3cd4c12d204f760758e873a177b;
reg                              Ic9146d8b3dd0c612073b70b8a8791e8c;
wire [MAX_SUM_WDTH_L-1:0]        I30b0b1d54912c1a41a02a25ab238bb54;
reg                              I857d3155df0b6dd704514b039c66fa97;
wire [MAX_SUM_WDTH_L-1:0]        I49fb0909ddf66fc0073e6400f1a07844;
reg                              Idc1b8aa2f81a7fbd87e4f5821d14bf01;
wire [MAX_SUM_WDTH_L-1:0]        I9938397dc94002481984f5b560fadc58;
reg                              I68b585571699a57bc6ba5e8955467119;
wire [MAX_SUM_WDTH_L-1:0]        I4378d139db4b710e3587aa72df22b70d;
reg                              Ib70e99c3acc76286a6811bcacc9284de;
wire [MAX_SUM_WDTH_L-1:0]        Ifa43d74fa91b7b9884969f575ef9ca8e;
reg                              Iee17ece482d04964d3c21a092ec955a4;
wire [MAX_SUM_WDTH_L-1:0]        I7c19a79f441ecbb73685db5a505e7479;
reg                              I5a247475beb737d470f03507e55f5b24;
wire [MAX_SUM_WDTH_L-1:0]        If2af8106efc1f7dd02c074af68278b3d;
reg                              I13b0c9578f7b6b3b7e6704d7b44079c4;
wire [MAX_SUM_WDTH_L-1:0]        I89a3f8d5f760d1a650f85814cbfdc017;
reg                              I41eff06fe1dea8be4613945de596d3ca;
wire [MAX_SUM_WDTH_L-1:0]        Ifae345c79662c3df3dff0fe68ad68746;
reg                              I08f22261d5713c0636d77c7938f592d6;
wire [MAX_SUM_WDTH_L-1:0]        I88a61cf72347d695489909d0819332ab;
reg                              I1c7e41b9cb1bdb6f649c88c0ed3f4100;
wire [MAX_SUM_WDTH_L-1:0]        I9aaa036a6158d11c235bdc8406d79f4c;
reg                              Idd59a5357d4c835379ed180ac0924bf1;
wire [MAX_SUM_WDTH_L-1:0]        Ie8df350430970b5f1229cda772440f85;
reg                              Ibe7e5c2cb9c50eca34a3859d13e83a92;
wire [MAX_SUM_WDTH_L-1:0]        I7d77ac9b64b2e8cae21c6e36947e3ca2;
reg                              Ibf5c141c5cc0a6a20c05b52bf8282476;
wire [MAX_SUM_WDTH_L-1:0]        Ic1faed76fca5a9ceb7db26c2f43623d9;
reg                              I0038305f94aaefe2cd1a243580d95932;
wire [MAX_SUM_WDTH_L-1:0]        I3ca2b9b77ed8d78a10aff42a07a53b07;
reg                              I5364deb983adc2ae505ed2b8c57f876d;
wire [MAX_SUM_WDTH_L-1:0]        I1f00849ea055a7893df386aed162a7b6;
reg                              Ifdb5589982db805a0416e1c01276249a;
wire [MAX_SUM_WDTH_L-1:0]        Iaf8a19fde3de660c3fa925593bebbe0c;
reg                              I8bb5522183b65583fda83067990b3e94;
wire [MAX_SUM_WDTH_L-1:0]        Icd1da43a4d95230e79dbd35a7ae41066;
reg                              I1e77fe6aeaba852aba34ed37dd53add6;
wire [MAX_SUM_WDTH_L-1:0]        Ice9079fb6e08d629f8c0c9ce332c8f11;
reg                              I9171019227f35760d02d0c8ce786f4d3;
wire [MAX_SUM_WDTH_L-1:0]        I15fafe2baba4d2f28037023a81ce0a81;
reg                              I6e92a48aaab94074a555efa9bd1e7243;
wire [MAX_SUM_WDTH_L-1:0]        If4d5b48882e9e628cf51ad2ac2f38c22;
reg                              I3bc094d67805664859fdcb66f1360e64;
wire [MAX_SUM_WDTH_L-1:0]        Id0eef1adba01447c14a6f005782dd9a2;
reg                              I2518ccf385b3b677d95983bc550282e8;
wire [MAX_SUM_WDTH_L-1:0]        I1d1a7c5928982c278d068ebd262254da;
reg                              I7547c56b32513ad45d775b4502596d9d;
wire [MAX_SUM_WDTH_L-1:0]        I6354a0e638340378124e4df7f3d145b8;
reg                              I013d84bfd582acc7accf07ec522961fa;
wire [MAX_SUM_WDTH_L-1:0]        I0236c912c6d684bf4862b725be9d5951;
reg                              I0ec27b590ee6dcdd9c1086105e3b6c23;
wire [MAX_SUM_WDTH_L-1:0]        I6f3be51d69b2b64a04e55b8946d5dd56;
reg                              I4cdc955fa9afc75c2c977de4ec540e1e;
wire [MAX_SUM_WDTH_L-1:0]        Icde3e6dbcf985682041f30903ad95572;
reg                              Ieefbb5d6f4ac1e586832c5c0f513c5a2;
wire [MAX_SUM_WDTH_L-1:0]        I46ee30b46020d91707689f3468f00e26;
reg                              Ic828cdd5dfde844df4c150921af2a443;
wire [MAX_SUM_WDTH_L-1:0]        I2605f078c1a9006c93855a9a2b0cf6b9;
reg                              Idf1ecab26889c4adcb835fda6b1cb368;
wire [MAX_SUM_WDTH_L-1:0]        I4d226dd2f0bfcdbea6a2e6a6613c1b64;
reg                              I00d3f14b20e1ea7d726533386e0eba27;
wire [MAX_SUM_WDTH_L-1:0]        I5c942076b173cf527e1be2ddb8560e84;
reg                              I7f720a18542528f0c9bfb14f699ff4da;
wire [MAX_SUM_WDTH_L-1:0]        Ic95191bccb18e26c10e56be395ca6b1a;
reg                              Ia98a6f01e4eb5bc74d50d350e79be426;
wire [MAX_SUM_WDTH_L-1:0]        Ia284f974dd8a526f31eb81ed71a06e94;
reg                              I182b43872d50de6f7afb700f178b160e;
wire [MAX_SUM_WDTH_L-1:0]        Icc93450a007cee4c0a42717ed7600528;
reg                              Ic9b72b2a91d951cf08cf54ed215ecaa8;
wire [MAX_SUM_WDTH_L-1:0]        I9ec9f389d0489908d497487e44c6edcd;
reg                              I93084ccf5b5e4efaee968b497bb2a775;
wire [MAX_SUM_WDTH_L-1:0]        If8a527cc7f06a9963a80a880d225d34c;
reg                              Id38852415486e6989b89a0d85ad6771b;
wire [MAX_SUM_WDTH_L-1:0]        I39ff4663007dbc89b403f3b08a69bb6c;
reg                              I17cf58ef5326978c62c03c56090a299f;
wire [MAX_SUM_WDTH_L-1:0]        I9590eb28a81c730b83b92ef7653e71a1;
reg                              Ie41ca18c7d11a47e274f9c33f75393ec;
wire [MAX_SUM_WDTH_L-1:0]        I2ba1acca919bddcc22a41a28d43a4e3e;
reg                              I7b80b4902fe98c10dd72c9eb082346e5;
wire [MAX_SUM_WDTH_L-1:0]        I62d8efd4227cb3dc88aa08b6585fafc8;
reg                              I20ffba20af04b99954bf719589e90d1a;
wire [MAX_SUM_WDTH_L-1:0]        I749e987266a20840bb8a4b1a2a2fc5b0;
reg                              If8fe5af7e5c3c97b5a713f6bcf919f1f;
wire [MAX_SUM_WDTH_L-1:0]        I7607af5d98e8070e3d15cee23cdf877e;
reg                              Idc5fb0f3a04ab32948e249e088a11b11;
wire [MAX_SUM_WDTH_L-1:0]        I2e11a697d7f17ac30302eadb500de72d;
reg                              Ia9f1e580e8f441394d719d52a7bad688;
wire [MAX_SUM_WDTH_L-1:0]        Ia0886ce792e062e22d0c224158cdfb7d;
reg                              I02849282dd1bd663fd39baccf41762f9;
wire [MAX_SUM_WDTH_L-1:0]        I6b3cd79aa87235ff174c0299b855dd3d;
reg                              Ie4cda4648f6ceb76b8fb74f290ab6439;
wire [MAX_SUM_WDTH_L-1:0]        Ie4ae993ddb776bdffec843db0def2f5c;
reg                              I24135210c23b2422a42c90ee25594191;
wire [MAX_SUM_WDTH_L-1:0]        I3ed2da9b53daac0852a06ad1acfad21b;
reg                              Ib08897f9216599042f7b97b137e07fe1;
wire [MAX_SUM_WDTH_L-1:0]        Idefa29d4d4e2a6e9147f84893520096f;
reg                              I51e14ece9ab6607f83e6ba27f3f046a9;
wire [MAX_SUM_WDTH_L-1:0]        Id1fbbe0594dae272856566522633bb3d;
reg                              I7a626ec321bf963a5401892a7e3891c7;
wire [MAX_SUM_WDTH_L-1:0]        I8070a3b7d8b1a7ae90c1a2d27aed09aa;
reg                              If76f04fe0baf171d7df2c0cd849aea2b;
wire [MAX_SUM_WDTH_L-1:0]        Ie88285ce2b9c71de02ebd62e8f44ca72;
reg                              Ia9c8cc5e3becf3d48feedec8fa2c93a4;
wire [MAX_SUM_WDTH_L-1:0]        Ica1997c6c569c1d1f45224fbaa4e6b59;
reg                              If3b77c41fabcdb283f2c6fdacaa5e9a4;
wire [MAX_SUM_WDTH_L-1:0]        Iaf08bcaaeb15bb0c971432f7f8b16d0a;
reg                              Ie5373b01a92f2ff85be8077cfef2175a;
wire [MAX_SUM_WDTH_L-1:0]        Idcb37cfc357cc088c775409fb9225b51;
reg                              I5109afc4dc91780e05704ea5e1399e3e;
wire [MAX_SUM_WDTH_L-1:0]        Ic419255414995e7168afb97b051fa64f;
reg                              I3e0b41bee4c76eb5f3340ad23bfa01ad;
wire [MAX_SUM_WDTH_L-1:0]        Iee6da3120d73373627b25ab7c0dedd28;
reg                              Ic0732810fd355d59a3168be896a0f9ac;
wire [MAX_SUM_WDTH_L-1:0]        I56fc99a22960232b305d6e683c66fcc7;
reg                              I220e32641265b46527ca61111f7ebf1b;
wire [MAX_SUM_WDTH_L-1:0]        I0a9a09b0ab43d2a0f1d1d01e13f0333c;
reg                              Ice59d2af73d0b0f2ae91a2ef0c2b7f04;
wire [MAX_SUM_WDTH_L-1:0]        Ibc73d07e0c97a6fcae791e04106cb082;
reg                              Ic308610ea8bb62ecb6094192e02dbdba;
wire [MAX_SUM_WDTH_L-1:0]        I224bbdf94ac86c5c376d1db4f4d4e060;
reg                              I33ee415d85e2bcd8f975d34b880f6ea7;
wire [MAX_SUM_WDTH_L-1:0]        I43f2b69c6b427de3095c44d4166b77cd;
reg                              Ie61f299252b8fecfd3e8634b64df5a90;
wire [MAX_SUM_WDTH_L-1:0]        I1e50c90010a3df1a8ce1cff811cc7a0c;
reg                              Icc67656ad2dd3fffae4e5abe02f8fff9;
wire [MAX_SUM_WDTH_L-1:0]        Ie1817cbf3a80dae435a5571dfbd2f5ad;
reg                              I0c47ccef4b55410286248884a7249703;
wire [MAX_SUM_WDTH_L-1:0]        I0052d562fb3182890c8828e52d437b11;
reg                              I94e4041b482064334fd0ed92b91bde89;
wire [MAX_SUM_WDTH_L-1:0]        I1eedecb1d8ff505c75be7787199afada;
reg                              I39d3bce4060032a81e6b6a1c1805cfe8;
wire [MAX_SUM_WDTH_L-1:0]        I7ef544597a185b1de63b4ffc4a1d44c2;
reg                              Ifb422c30663eb4824caa72326b238df6;
wire [MAX_SUM_WDTH_L-1:0]        Iadeedf3870f0b1eae98d0f7dbbeff04a;
reg                              I41ab6fb6ec6ef7ffff70e50f25f217b6;
wire [MAX_SUM_WDTH_L-1:0]        I70ae07db9b44d530be220f06401d3d3d;
reg                              I3ce10718a2211184999663c3c2493cc1;
wire [MAX_SUM_WDTH_L-1:0]        I7992ea31927b4f0e268462a3b0f18c5d;
reg                              I877e8d94236c3d8b0a31858a98fba5d6;
wire [MAX_SUM_WDTH_L-1:0]        Iadf927d18644a232ad1f1eba7db82934;
reg                              Iff2f1716cbd73b406d8f07c22dc79fc8;
wire [MAX_SUM_WDTH_L-1:0]        I2a9c673cdd7ded79e09ada38c0f47e6f;
reg                              Ibc48fabc172f27ebce18d0a9b5120dc5;
wire [MAX_SUM_WDTH_L-1:0]        Ia86740e870d8063f0266b68ad6d7481d;
reg                              Ie562ebb336e476a81f20a652d4cb20f1;
wire [MAX_SUM_WDTH_L-1:0]        I6627bcdbaa8afb115123777abd45435b;
reg                              Ib5ee5a6ffc45ed1fece0822dc4619b57;
wire [MAX_SUM_WDTH_L-1:0]        I96fe3eb633eff6958ac575b997460bb9;
reg                              I86ba73ee348f80e2f9891d2ebc8a02ed;
wire [MAX_SUM_WDTH_L-1:0]        Iefdcb71f2903b11f5cb0b8857f7a1727;
reg                              I1e96d5af3d0e3fdce39530dfd0131a7d;
wire [MAX_SUM_WDTH_L-1:0]        I2eb90278aaa54b9c8212b3b4af7c3617;
reg                              I38352b363fa37f6f822fbc1a39100968;
wire [MAX_SUM_WDTH_L-1:0]        I43493f70f0336453d77caf7f27503daa;
reg                              I4ba41864bb1d2130c6971e0b2903027a;
wire [MAX_SUM_WDTH_L-1:0]        I26a7fe395eb583258c1ac58aaaa3234a;
reg                              Ib68deeb7bec4ca3585d1a4dcbf8793f1;
wire [MAX_SUM_WDTH_L-1:0]        I21668ff77cf75570cae97f575cbcf644;
reg                              Ida3d808d100e0bba290f96ed9e744e65;
wire [MAX_SUM_WDTH_L-1:0]        Ie48be9e6b6fd63baa104d0a6a4561a1a;
reg                              I4d4901ff372f6820ca9c8c29cefa664a;
wire [MAX_SUM_WDTH_L-1:0]        I05370777439b01811fe7f750d2f724f4;
reg                              Ib99e1b93fb7fbda260d93eea3d24c3e9;
wire [MAX_SUM_WDTH_L-1:0]        Icdcd83341f6b5c404f91ec7e97d0550c;
reg                              I019e399a1cef87745e025a7d74e94db0;
wire [MAX_SUM_WDTH_L-1:0]        Ibba4e82d1510ddc16eb4ef64893cec02;
reg                              Ia8974083bfd064f2c27dcd421490fcfd;
wire [MAX_SUM_WDTH_L-1:0]        Ifb00ae47340bc99669c71da34cccc59e;
reg                              I8fd5787ebf758919e7cb75d7419441e8;
wire [MAX_SUM_WDTH_L-1:0]        I75a4cf2948bebc58e12bb039ed273ff2;
reg                              Id14074d5230885c38b89b09b130ecf68;
wire [MAX_SUM_WDTH_L-1:0]        I5a9fdec7d7ff99fe33ad6cd8afd9e059;
reg                              I86fefad34d3c864dd0e725133f303b4f;
wire [MAX_SUM_WDTH_L-1:0]        I47b1695a74e4d27389b97543415dcc67;
reg                              I1ca188bcdebbf41d84f7a5220bd1d195;
wire [MAX_SUM_WDTH_L-1:0]        Ieb38fa62119a5a77c060d6634e051298;
reg                              Ifc640243288c9b37b7eb9e00351b23f0;
wire [MAX_SUM_WDTH_L-1:0]        I3459d98131faef5a5040a03847890b55;
reg                              I3d149293f106ae8680c7f4702daa0bd6;
wire [MAX_SUM_WDTH_L-1:0]        Ie9b9221b2122087cd5f309570b6d31ca;
reg                              Ie232799bd6c4ec99e24c78f3ad798265;
wire [MAX_SUM_WDTH_L-1:0]        Id4451722e8e2393d627dcd0175dc9903;
reg                              Ifebcf64858d5e2d07ad7894d6182eb11;
wire [MAX_SUM_WDTH_L-1:0]        Ic10356f9069e3651b9c045c906e63512;
reg                              Ibab55499323660588ec82ebd07ab0572;
wire [MAX_SUM_WDTH_L-1:0]        Ic3a431f39c678b7175ed30fde1fa6424;
reg                              I89af7644c48a80d7d22f50b008d35841;
wire [MAX_SUM_WDTH_L-1:0]        Ib01cfd833a63500e03333f263805db3d;
reg                              I0152dc6e6a7acd72a2144623e63998ef;
wire [MAX_SUM_WDTH_L-1:0]        I0b7b4c0a8503c751229edfe0237cc903;
reg                              I951dedd7af44c3865a8f36888432d0c9;
wire [MAX_SUM_WDTH_L-1:0]        Iace01234164c8a9f7c98eeb83268745b;
reg                              I8188dd7cb03854c6f709de06ff785d91;
wire [MAX_SUM_WDTH_L-1:0]        Iace8b3b3a4c16763132b5aaa6b24212d;
reg                              I3b30b4ab00a49e10a75587aa324d6132;
wire [MAX_SUM_WDTH_L-1:0]        I80a89644e278e96b1cd1c4b7f764dc34;
reg                              Ie50aca688b3433fad7565998cb900155;
wire [MAX_SUM_WDTH_L-1:0]        Ia92d2276a8a23521ad1b88df7c27bc2e;
reg                              I3342fe0c5d3ee5021892d53eb45bde21;
wire [MAX_SUM_WDTH_L-1:0]        I39bbec42c442d1e8c818f46ad9c096a8;
reg                              I5134b762ac428bed07ce102d8927a418;
wire [MAX_SUM_WDTH_L-1:0]        I88f1b5c12759a5efb2d2ded8483c9ed2;
reg                              Ic14f948884da19a272a4760ffaab9ea9;
wire [MAX_SUM_WDTH_L-1:0]        Iaf4ae293c576af16f5f43a8b86c1aa3d;
reg                              I46e1047bca2b38e62b4de80d1d2249de;
wire [MAX_SUM_WDTH_L-1:0]        I68b575fcbc5321d4d26a22bcdbb506f6;
reg                              I866b30a63b3b5fb708934a1cbb0e1d9a;
wire [MAX_SUM_WDTH_L-1:0]        Idf600b93ee1018ecf969ed7944b6bc7b;
reg                              Iaddc1f2e822fd2fe9d9046d759a82cb4;
wire [MAX_SUM_WDTH_L-1:0]        I1cd93172cf5996bc870063aa642188a2;
reg                              If9285bf7611bcc5ea6432215c349e021;
wire [MAX_SUM_WDTH_L-1:0]        I4af080cb4e5cc525db95e5f401019e8c;
reg                              Id277f5f05551eeb5dec1701056330da1;
wire [MAX_SUM_WDTH_L-1:0]        I6fc8044eb226a14ff1a786ddc96d2414;
reg                              I9963d0b24763ed8038b1f3922b8f9548;
wire [MAX_SUM_WDTH_L-1:0]        I27fd0073dbcdee599fbe85cf48806efc;
reg                              Ia98de3691917dfb63bebdc3f8655c8be;
wire [MAX_SUM_WDTH_L-1:0]        Iaee6d725a8b2653eeac6d5acb91f8f36;
reg                              I0bce960fcc58938e6a1e01b912eabbf2;
wire [MAX_SUM_WDTH_L-1:0]        I4afdeba4fc2a12a6cbe3567a519367fc;
reg                              Ice5f7168aeb940d48093cc9df7cba36b;
wire [MAX_SUM_WDTH_L-1:0]        Ib42816335dd8475dcc78662c4c0786c1;
reg                              I859d795a7d141eb777c1f3c038203794;
wire [MAX_SUM_WDTH_L-1:0]        I343c9efe71164c01e9c7d599e032864a;
reg                              I0dccb8eaad52ce4d780696a8485420f1;
wire [MAX_SUM_WDTH_L-1:0]        I108c269ceec4adcff9afeda01101b838;
reg                              I6d4fc81ced37c159303c243af04d345e;
wire [MAX_SUM_WDTH_L-1:0]        I761983331fb6e3c6c437b3f1660f0b6b;
reg                              Iefdb8bd28839af9413a3906cbfe715e6;
wire [MAX_SUM_WDTH_L-1:0]        I70d32affde22f9dcb2d77430fca39069;
reg                              I0615acb0f7cf79b5f6ae8e91cb525dc9;
wire [MAX_SUM_WDTH_L-1:0]        Ic08e85346f61da036a15345a13ac12f0;
reg                              Ieed4c810a5bb69de112522dcf00b16ed;
wire [MAX_SUM_WDTH_L-1:0]        If5dfdadb3868ed5a495007362f7db648;
reg                              If533578cacb685a95afbb8e1c05d3c07;
wire [MAX_SUM_WDTH_L-1:0]        Ia1ee5579358b564de06c08ca418a9bf4;
reg                              Ia858ff5551286beffd4cf82f876d30ac;
wire [MAX_SUM_WDTH_L-1:0]        I9bb81dda8102b829441be46460eb8900;
reg                              I4c66570630a650fa7b9bec543f685487;
wire [MAX_SUM_WDTH_L-1:0]        I8eef6ca0a61a21882ea28b3d63735228;
reg                              If10f33385e236eaba56cbab8c2883399;
wire [MAX_SUM_WDTH_L-1:0]        I438522d92cce6f7010246424746ca255;
reg                              I7cb58e4c486e683faa4acad4756815d5;
wire [MAX_SUM_WDTH_L-1:0]        I92496f68b44a94565af28a2c28d6fbae;
reg                              I452e51cca9acec44e36e4efd21b43034;
wire [MAX_SUM_WDTH_L-1:0]        I66528f43f614f0edb715564eba3c77c1;
reg                              Ice0234f25de4ab1f03a3cb01a2d61dbf;
wire [MAX_SUM_WDTH_L-1:0]        I8cab9fba615b94fd4bb6934325be8ab8;
reg                              I12a18a1f8d4416e9bc8abee6ac3dacfc;
wire [MAX_SUM_WDTH_L-1:0]        I92d9fec22d36b1baac8bd78abfc1bbd5;
reg                              Id17ada8dae3f9810d1892d34f2288859;
wire [MAX_SUM_WDTH_L-1:0]        I4eadce87f47df6d8f0e4acd057de5a09;
reg                              Ia2c5fe53cb5b318fa63d09881609655f;
wire [MAX_SUM_WDTH_L-1:0]        I73203143fe37933c16fff873c1abf512;
reg                              I579c7926e7b78f4ffc606adc10522f53;
wire [MAX_SUM_WDTH_L-1:0]        Ibed2a63af723a7abf96dacf1951e5266;
reg                              Iffa06a336949f56f4e5a88a06d8b7e60;
wire [MAX_SUM_WDTH_L-1:0]        Id667c80003b5541de9f84d3b8709c828;
reg                              Iaf82668eb49248709540f2f529f1b3e4;
wire [MAX_SUM_WDTH_L-1:0]        I02cbb4255db2b21ea32140f9e9ddb36b;
reg                              I90b3708abdf742370f06cc513ee307e1;
wire [MAX_SUM_WDTH_L-1:0]        I65354f2069de0c25bbe7cd50fbe892aa;
reg                              Ia17906696bd0e095d7a5297da2e049ea;
wire [MAX_SUM_WDTH_L-1:0]        Ic279867ebf3055980f3d813d5dc8dec6;
reg                              I180d4f3b23b518271d7cb8189fbeadc5;
wire [MAX_SUM_WDTH_L-1:0]        I5c05da8a222ad5effb9815cbf3ec25f3;
reg                              Id79636d195efff260c430978f0bcee9c;
wire [MAX_SUM_WDTH_L-1:0]        Ib8bf21f32c0e8b9cfa42a53807bfe3a3;
reg                              Idbf4ad11ab2a27044193448c8739fec6;
wire [MAX_SUM_WDTH_L-1:0]        I7208256bb198bfce1be71390b01bc028;
reg                              I3051f561a5e1131ebf167cb6ccb5adf4;
wire [MAX_SUM_WDTH_L-1:0]        I49f2a06ceb3a59773c65b19f54ff362b;
reg                              I9322a2a61900943075bbc23c72a3f65d;
wire [MAX_SUM_WDTH_L-1:0]        I86e495dc894d2aace15c1aff89798bf7;
reg                              Iedc463e359dd3003d9f7e50f3e858e93;
wire [MAX_SUM_WDTH_L-1:0]        I0d53bb5344cabe5fa5ce3ecf7122a260;
reg                              Ie7cfdd25541414ff3f8d6e5d7677fbe5;
wire [MAX_SUM_WDTH_L-1:0]        Ib2f5f5fc77ea8b529f2471c54388f2d1;
reg                              I1e93f0470d2818249f1c28ef2a399a0e;
wire [MAX_SUM_WDTH_L-1:0]        Idcada1bfb3c0d1f2a09aab58a2071a57;
reg                              I5d6e576b0fa7e3219aaf9ccc345085b8;
wire [MAX_SUM_WDTH_L-1:0]        I814b62120953991f9da055f118967e05;
reg                              Id962beade26396738ba0e97f67d5e261;
wire [MAX_SUM_WDTH_L-1:0]        I123a212546a8ac394051425db4924812;
reg                              Id0ab747d92288f23cef793567b2363d1;
wire [MAX_SUM_WDTH_L-1:0]        Ie95f1a7e0effcec0aa423dc803056a13;
reg                              Ie536879e6fa9be65376d7f00e0fc40d0;
wire [MAX_SUM_WDTH_L-1:0]        I106deaff50b8480eac31ddbae2ec7c61;
reg                              Ibf312ae4f51fbc44b43848f9df62a45f;
wire [MAX_SUM_WDTH_L-1:0]        I68528be9951f5b8805411711cd11ea59;
reg                              Icfc03646b36b971b9fa57d04a26dbfc4;
wire [MAX_SUM_WDTH_L-1:0]        I0f034a8f077b0ab231727b6298e366d8;
reg                              I4f134c0669b5a6a8c7e03be7eee30c6c;
wire [MAX_SUM_WDTH_L-1:0]        If9c12f8662333fb54a45cfa1bc5da487;
reg                              I6c765e677f42fe600b848698c8a78349;
wire [MAX_SUM_WDTH_L-1:0]        Ie1681d905517daafcc7584725cd6014c;
reg                              I284b23051c85300c2a1e3afe8f25e99e;
wire [MAX_SUM_WDTH_L-1:0]        I2ff3edcdb6158f1e3c9a555aeefc0850;
reg                              I9b560d9baf8a7422b0dd84720e924ced;
wire [MAX_SUM_WDTH_L-1:0]        I43b380be6df7df0d354223d0a0d6d6b6;
reg                              I457ae11ad90c8478751eb4b42764e158;
wire [MAX_SUM_WDTH_L-1:0]        I23eb1dc4d1c992f804dd04a2d823c778;
reg                              I2b7822d5d77aaed61eee87570564df76;
wire [MAX_SUM_WDTH_L-1:0]        I7f90f96c0260560ad5e6dc7448b2670a;
reg                              Ibdad0ab78e4404c852e60a2b04c3a5f6;
wire [MAX_SUM_WDTH_L-1:0]        I07b417cdcc99eaea3413f563e26ddc73;
reg                              Ic4efba3932e598784f5b9ad6ad04772d;
wire [MAX_SUM_WDTH_L-1:0]        I2f3ab9654e515a54e22e73d6c130ccc3;
reg                              Ia03836a4e93d2f36513227d1dfaea0fa;
wire [MAX_SUM_WDTH_L-1:0]        Iebdc41368d57498a04fa73e30b10a966;
reg                              I138fb0c48f2d27e3315e237d9e61d653;
wire [MAX_SUM_WDTH_L-1:0]        I5b4305bef5b4350c1d7ae143667afddd;
reg                              Id0b1c46fa4caa63a4c63a44ba3c5ef8a;
wire [MAX_SUM_WDTH_L-1:0]        I2795d21d343b83a69146314a2407cfa2;
reg                              I3566033cf5c9a06977c9182925750707;
wire [MAX_SUM_WDTH_L-1:0]        Ic6386d7d8813731d612e24b715740275;
reg                              I02812a8a833bb69eb168a1004b6fafdf;
wire [MAX_SUM_WDTH_L-1:0]        I4c366a57920ff090a98a2cb8b9caa00b;
reg                              Ie886c5effc85f1fe0b6411db4a2cde77;
wire [MAX_SUM_WDTH_L-1:0]        I14cf5d43fc9864820a8a25efcc5c6d86;
reg                              Ibab1d13cd6a4f7b0c79c9f845339e53f;
wire [MAX_SUM_WDTH_L-1:0]        I33b99994abbb5ecf8eed4de39033e4f8;
reg                              I7b813d83b13bb7bc13940cf5714c06ba;
wire [MAX_SUM_WDTH_L-1:0]        I7c3291f0250d13ca94802b0b071a95c6;
reg                              I09031235f61238b0e32ff52641aab70e;
wire [MAX_SUM_WDTH_L-1:0]        I2c926fd9d306e9ae13364e07c4b0395b;
reg                              I5402fd208dc7ca81dfd2920a9cfa2715;
wire [MAX_SUM_WDTH_L-1:0]        Ib23edc35fa5bbfe0415fcf0861a22d9b;
reg                              Ia01c82761aeb124cd92fb15ee367ee8b;
wire [MAX_SUM_WDTH_L-1:0]        I3e0e682047f7cc36142e668828cbff1e;
reg                              Ib1a40247057324b0bd810c844bf11f51;
wire [MAX_SUM_WDTH_L-1:0]        I99fb9030e8361e57818c07511479a9b8;
reg                              Ied8bd4b6fd0e4fbcced6d20eb7435f55;
wire [MAX_SUM_WDTH_L-1:0]        Ic87c3d7762a18772972552162e1d1a8c;
reg                              I4ee312036de8c08300c358edcff1e1e9;
wire [MAX_SUM_WDTH_L-1:0]        I7e393e6c1d1bc44daaab120d55f5dd59;
reg                              I477a920e2326828bf026b0a6b6a18e2b;
wire [MAX_SUM_WDTH_L-1:0]        I448f126fd3932d5065abbe7bb2d92c56;
reg                              Ic11a6b77b84c44180eb99220a0c4c9f6;
wire [MAX_SUM_WDTH_L-1:0]        Ifc8c6df8904b97674f2970ebc95b523c;
reg                              If0970d9f7b053fce3ced3521b4885588;
wire [MAX_SUM_WDTH_L-1:0]        Icd0622a90782b9c451950e7ab0399567;
reg                              Ic7ebdc317c978eb275eca41d5b9106a5;
wire [MAX_SUM_WDTH_L-1:0]        I6493b3c087d4685a6b3f98c73dc2ff49;
reg                              Ibe3d3e6bc58efc2e9d9eb1f96cdfe424;
wire [MAX_SUM_WDTH_L-1:0]        I20c2057240417146df144b518b43d052;
reg                              I1dd4671765f8826c2fe20c592c5e32c8;
wire [MAX_SUM_WDTH_L-1:0]        Ied029d0bdea3bf134744c99426fa72dc;
reg                              I6cde57127c5bd2732e71ecb7738fad6d;
wire [MAX_SUM_WDTH_L-1:0]        Icb82c9ff4cb58159a1c3115c6fdd5f8c;
reg                              If6ce2fa9f0b8bc74442ed8262b5089cf;
wire [MAX_SUM_WDTH_L-1:0]        Ia3450e134e4086c35acbdee1e6042396;
reg                              Ib0001d7298ad1f3b1c7603173a70d8b5;
wire [MAX_SUM_WDTH_L-1:0]        I5a0f27df5158309f32f0df31e8ae3ae3;
reg                              I05e739fc87e962848f265e2c73338cac;
wire [MAX_SUM_WDTH_L-1:0]        I17d9e19854cef197fd3267618617efc3;
reg                              Iaaaf373f7e6f55214915b93da9bd71d3;
wire [MAX_SUM_WDTH_L-1:0]        I2993acb61f1abe529f8a60c94a438550;
reg                              I47b0847946b0e00961233ac0101fa2a7;
wire [MAX_SUM_WDTH_L-1:0]        Ic8be2c94235fb40f78da33179ce4873a;
reg                              I2f23d4cdb6f5f827513aa60266936e4f;
wire [MAX_SUM_WDTH_L-1:0]        Ib3367565e4456da15e7c2315dccdb5e4;
reg                              Ia67f9b902a21de0414eb8dda52171991;
wire [MAX_SUM_WDTH_L-1:0]        I15a1671def323cd294591564ae6ef8b1;
reg                              I87b10521099179c18652c86d5887c908;
wire [MAX_SUM_WDTH_L-1:0]        Ic512effb493a06ece58a2af155135004;
reg                              I84057a3b319ab3d6a2ed8f2310f970fc;
wire [MAX_SUM_WDTH_L-1:0]        I2c72248cbe49ec0a0febac2437b8a6dc;
reg                              I67d57e38df8cb35ca686ac2eb44e233e;
wire [MAX_SUM_WDTH_L-1:0]        I964e17c41a134c080e9c43412a514f3f;
reg                              I23955b54e486f0f0d21a2809a9472b86;
wire [MAX_SUM_WDTH_L-1:0]        I94f1724740defe5bb7e40041d0e266a0;
reg                              I1e11f0088959aa40b4ad1a047b59caf4;
wire [MAX_SUM_WDTH_L-1:0]        Ic19486b6ab0373b9c0ad8f7597782d8f;
reg                              I68c35d63dc95baff41b4dc27a86d2342;
wire [MAX_SUM_WDTH_L-1:0]        I31243de90dc2a1656ca9d5e03bdd78da;
reg                              I837183265ee22d080e81fea468ab0887;
wire [MAX_SUM_WDTH_L-1:0]        I242a30bdc8699d8ff550b25dd53d6c59;
reg                              I413b1c1985a6c9c6f202e85ff901e3a8;
wire [MAX_SUM_WDTH_L-1:0]        I9d15f76bb68b214057566cba4b511214;
reg                              Ic32c6734132776c290155a80025fe366;
wire [MAX_SUM_WDTH_L-1:0]        I9cc16a00912e7dfc05fb505a9db23cd8;
reg                              I624958486d181501c7a8ec2642cb503c;
wire [MAX_SUM_WDTH_L-1:0]        Iacf9640cbf486411d6ceb8fe1a2fd5c9;
reg                              I04864c28351edb33b61a103add6fb875;
wire [MAX_SUM_WDTH_L-1:0]        I9015033ab0caf3fa41dae4de43f24a82;
reg                              Ida3dd5e990ce3c237e9628a9a090901e;
wire [MAX_SUM_WDTH_L-1:0]        Ia630e59cbce82a570ae3890a6c0221e5;
reg                              Id182a776b03f48fb139c28194ae7ab6b;
wire [MAX_SUM_WDTH_L-1:0]        I4904ab14b19fa1b6befc218bc7be3842;
reg                              I0c5539373b3868d0664a92157b4b4226;
wire [MAX_SUM_WDTH_L-1:0]        I282d2eb4e74e034694e33273b9cb19d5;
reg                              Ic0191941cb968bbd7644c21767423d2e;
wire [MAX_SUM_WDTH_L-1:0]        I3f33901c407a87e10d86c13c83dd52eb;
reg                              I163cf58b9a308e0439a8dc7c1526e6b5;
wire [MAX_SUM_WDTH_L-1:0]        I43f41bf07836cee48069e9890c1de2a0;
reg                              Ie08ad9bd71329858c1742c8f571a1c36;
wire [MAX_SUM_WDTH_L-1:0]        Id88480a0a350bb5fcf01ed5fff0bbd4c;
reg                              I3c10d579f80bd0106506ad047d75f188;
wire [MAX_SUM_WDTH_L-1:0]        I1d9b9ff357667a362f0442f19986f451;
reg                              Ieca2767ac27170058499d83016447aa7;
wire [MAX_SUM_WDTH_L-1:0]        Ice73589836da9028def6efb24a04dbbd;
reg                              Ib9c194ec16f435a9357cb344cf25bdcc;
wire [MAX_SUM_WDTH_L-1:0]        Idb72c046c5996fbbd80b706666ffbd92;
reg                              Ic920452d5997a8477724fa78c86c0fba;
wire [MAX_SUM_WDTH_L-1:0]        Ie5757e7b1647ab7d43cdbcf98cbb77fc;
reg                              I6eea5fde8e2517554ad6ba25018572dc;
wire [MAX_SUM_WDTH_L-1:0]        I6072331f838d82329a07a4ffa340c7b6;
reg                              I9ad2f6fd2d7f68011fc926ec9abd5c34;
wire [MAX_SUM_WDTH_L-1:0]        Idf6875955525d80dc660ce956f4a84e7;
reg                              Ied33f18cbb778d5ba744d249f91c950b;
wire [MAX_SUM_WDTH_L-1:0]        Ia96955d9c0a8a587e0afab37c8415d8c;
reg                              Ibabf61085ca7af8dfc7927b3656a76f7;
wire [MAX_SUM_WDTH_L-1:0]        Ifec374bce7f5507438f550df22d61a01;
reg                              Iddc5b5b4501f9f13bcaf22081e5a70f4;
wire [MAX_SUM_WDTH_L-1:0]        Ief67e897e57b96e2ec200e82bbc7caeb;
reg                              I67f87fbb746dd937fffc534c596f36c4;
wire [MAX_SUM_WDTH_L-1:0]        Ide604e9bbe35cb55892a4602e18b2527;
reg                              I45bdd0cfe107da0d57cad1333bf95e3b;
wire [MAX_SUM_WDTH_L-1:0]        I262f2390e77ec486ccd3a6ed05816e2d;
reg                              I4d54dd2ee2f32909098d3cc2b6689220;
wire [MAX_SUM_WDTH_L-1:0]        I280e20c20c0b4f26278b3de9b2ff84e4;
reg                              I7bfb4c5d9e22d1bd8811844d9c74dff8;
wire [MAX_SUM_WDTH_L-1:0]        Ib3a0307176d424a4733720416d71069d;
reg                              Ib9d58222da98f29fa302b4896594fe26;
wire [MAX_SUM_WDTH_L-1:0]        I76060709de3ea188748849f043c59ac0;
reg                              Iea3e35ece9fdb3aff3b9ff5369e9a7e0;
wire [MAX_SUM_WDTH_L-1:0]        I8be20605d26d218911e80a883a90d085;
reg                              Ic44eab478be232721e7a43d14beca32f;
wire [MAX_SUM_WDTH_L-1:0]        Ieafa9d74d4a61d28ac4a913db460bf33;
reg                              Ifab075b1437495268b6a3be4cb022e71;
wire [MAX_SUM_WDTH_L-1:0]        I6fd1b4395af175eff85b3bfeef4c329b;
reg                              I2919272e9ae3996a3e1d602ff72ba86d;
wire [MAX_SUM_WDTH_L-1:0]        I39e6d3fb468aa40ea73535e81556ea65;
reg                              Ib6fbe376477afa58bfcc17a8564f78b2;
wire [MAX_SUM_WDTH_L-1:0]        Iae449b74e50e0907feae9e60f2329426;
reg                              I659322a9fd0d5eac514437b02e0491b3;
wire [MAX_SUM_WDTH_L-1:0]        Iebf769a6bdaf214c1006c55c608d4eda;
reg                              Ic68f500938d80460ffdb33a0adc48298;
wire [MAX_SUM_WDTH_L-1:0]        Ia030c08757123aae947f86ab8bfb6d94;
reg                              If5ae6fbf843fdeee17945bc5ce81aec8;
wire [MAX_SUM_WDTH_L-1:0]        I8c35c5b343b552c22000e194c517ca12;
reg                              I94460b6ce7b776bcc5eca149eab80c26;
wire [MAX_SUM_WDTH_L-1:0]        Ibf80bb564263ea85bd886a8617f09bb2;
reg                              I3347717ba9556e69de30ce7533d4f5a4;
wire [MAX_SUM_WDTH_L-1:0]        Ib8dfd9b8badef282ca00a4f793c3c868;
reg                              I2db290170ddae8dc52ce07edaf48b365;
wire [MAX_SUM_WDTH_L-1:0]        I596ad7e132f272cb196b74faa8c75aa4;
reg                              Idd775d9fe6fa8dbdbfb07d4071b9caa5;
wire [MAX_SUM_WDTH_L-1:0]        Idc629414f6d0236ce0714cfaae23f065;
reg                              I6cbc06919b9c695d99621db6f8d768cb;
wire [MAX_SUM_WDTH_L-1:0]        I157fdf8775206858c08682db3039b084;
reg                              I5b8a1e1a6b904b0f6822c224ee0486e3;
wire [MAX_SUM_WDTH_L-1:0]        Iacbb4daf5ce5c7eb1a2afe30d0cb5382;
reg                              I3f5053e519a928640ae49cf4e5b39d1e;
wire [MAX_SUM_WDTH_L-1:0]        I4e08021c0235fafb60200aab97827a8f;
reg                              I7c965c047d862c973d09a81abe03a845;
wire [MAX_SUM_WDTH_L-1:0]        I730634ea15ac94d241f3ad2d6393a227;
reg                              I9b8023f4dced915cd52c91bc9d4ed78f;
wire [MAX_SUM_WDTH_L-1:0]        Iee367c535d9c39f872d2ec043e7e7b33;
reg                              Idc6b6357741c9887a9db1037ccc2d922;
wire [MAX_SUM_WDTH_L-1:0]        I68bb1f26f878862f288c1f57049cf58b;
reg                              Ibe97860165dc5d9a076ebd935385ae51;
wire [MAX_SUM_WDTH_L-1:0]        Ia9b5d9ede006c56a6d83905529c77b7b;
reg                              I777ee54ff20d0544af18ad8a870d6915;
wire [MAX_SUM_WDTH_L-1:0]        I1487170cb1f3370ad45efc801cefc8ab;
reg                              Id18c5a1d4eaa73a94e699e5f9e3c3d35;
wire [MAX_SUM_WDTH_L-1:0]        Id88568dd34fbee42c9cb8cc15ac5c31d;
reg                              I72939e49bf2d9c6a84e404419fc644a1;
wire [MAX_SUM_WDTH_L-1:0]        Ia30539545e66c4cfc16828140149180a;
reg                              I57b7b48f13436b19a8d6a47e014eb41f;
wire [MAX_SUM_WDTH_L-1:0]        Icbfbb37bad6344005dd233b3605a784f;
reg                              Ia3ef2f70c5abaa852586a33c505aee0d;
wire [MAX_SUM_WDTH_L-1:0]        I91a6408a11fab36a8ba3dbd3f895a803;
reg                              I6d423a7d17e05a3c597ec6ef6c5a7cba;
wire [MAX_SUM_WDTH_L-1:0]        I47b878f27c30f79a37e97e022307e9e9;
reg                              I48e3309c61918c3991852b45d9c72ea5;
wire [MAX_SUM_WDTH_L-1:0]        Ie76b0739aec66f8860870e66e87a6445;
reg                              I472352e7027b9df2fa957d9fd68443ff;
wire [MAX_SUM_WDTH_L-1:0]        I50383e3d7c172eedfa00aa50a9faac4c;
reg                              Idbbf2ce4a30787c5f07c3b908a73da75;
wire [MAX_SUM_WDTH_L-1:0]        Ifeaa99e03bda8ded058f98387de3d49d;
reg                              Ibc9a860879ccc58c815b9f6caa23320a;
wire [MAX_SUM_WDTH_L-1:0]        I4255ac1af4367c321567c4e46b06ab25;
reg                              Ia71cf07b645c58cffe33be1a9a960eb2;
wire [MAX_SUM_WDTH_L-1:0]        Ia445bdc7def7d8c1eec31ab892c25c41;
reg                              I0ceb14ac0187d804f9692e0c55b8e941;
wire [MAX_SUM_WDTH_L-1:0]        Ic3b4752136ac08e343933ccc3a4ec47c;
reg                              Ief18a19d451f05f6051e3cc8de16d73c;
wire [MAX_SUM_WDTH_L-1:0]        Ica6707efd6d44ba6bbb87c0593a3d828;
reg                              I30be0b18e4415ca50f2d8149efaaafe6;
wire [MAX_SUM_WDTH_L-1:0]        I739267bcc50c54b8a685cb3c6afc5cc1;
reg                              I7ec15b73b2811b44e1e50c74a9f921e9;
wire [MAX_SUM_WDTH_L-1:0]        I9160d11439c5140c0109b5190eb82e6b;
reg                              I0fd2f706e374a4eb57ee26ab50201e15;
wire [MAX_SUM_WDTH_L-1:0]        I6ff7b86cd7f63f9243646f1be10b2577;
reg                              I44f170d02bae7fe044456e125a98451d;
wire [MAX_SUM_WDTH_L-1:0]        I165653ab165cfafe2b74cd441331f9e1;
reg                              I30c0fcd89e0cc7c5fa348df7b4fa2ccf;
wire [MAX_SUM_WDTH_L-1:0]        I08a8cd6965c23af6650568b654831b20;
reg                              I13a98f98c54b2e412cd88c96f016c41b;
wire [MAX_SUM_WDTH_L-1:0]        I9b6a674dbcbfcf65f1ae0deb8fc3566d;
reg                              I9890f7fc708c7b8cf460849b4a30025b;
wire [MAX_SUM_WDTH_L-1:0]        Ie3a336de822ac7baf8486b1618ef1126;
reg                              I5e69e930a318dcb0594a823b3129d650;
wire [MAX_SUM_WDTH_L-1:0]        I5fc3c26d6c5aa893dfd5caa0f677233a;
reg                              I403303228c0df825f67436f4a7e64061;
wire [MAX_SUM_WDTH_L-1:0]        Ie22b94121b58f17af14c75bfb27f96dd;
reg                              I946246be5b4745508b7d4b578f83aaa2;
wire [MAX_SUM_WDTH_L-1:0]        I0d9f8c99194d9d6e187b4ad02fcce8b4;
reg                              I95f0acd4f955058041c035789c3a4d99;
wire [MAX_SUM_WDTH_L-1:0]        I71e101962e766a4d1484b3235359a4b5;
reg                              I4082b3564c1949a19ed35bd5a88e1ef4;
wire [MAX_SUM_WDTH_L-1:0]        If2539da6722562bbf31786fd0036666a;
reg                              Ia7606050c683ecefc510ba92ac539a9c;
wire [MAX_SUM_WDTH_L-1:0]        I22c8ccd4a9018ad1c129aa058bf579d8;
reg                              I5446c1c323774715371c73bd1be66697;
wire [MAX_SUM_WDTH_L-1:0]        I83330fef69470d2f5def8e6d7d9c50d2;
reg                              I3a8e9e7d2cd6751e8500a5567cef5acc;
wire [MAX_SUM_WDTH_L-1:0]        I0539d598bbe3d50940329a282c801328;
reg                              I621b20d29d3a9a9f41065bc3c3bbd2d8;
wire [MAX_SUM_WDTH_L-1:0]        I202f88fdc946494d55fc8831c2e8a34c;
reg                              I263aad78110a1136eb7012c6983b2a8d;
wire [MAX_SUM_WDTH_L-1:0]        I3ee10f6a7785a236db317515fdd23a2d;
reg                              If4308ed204e33952c9931f8fe257aca4;
wire [MAX_SUM_WDTH_L-1:0]        I453fdf4fbb5af5bd28a20d7643da9eb2;
reg                              Iddcfab4a7022e0f12fd20cb34e9b9d02;
wire [MAX_SUM_WDTH_L-1:0]        Ic4a6c02880a9aead7353332708e3f388;
reg                              I759409e242eaeb144a53e630a8cfd514;
wire [MAX_SUM_WDTH_L-1:0]        I7fb3b66cb48521f8715f66bf5642cdb2;
reg                              I5f96a68d20e3ebc71dad4b43305baa20;
wire [MAX_SUM_WDTH_L-1:0]        I2fd872df07f50688486c0d602cfc5549;
reg                              I5d92fdff96b9cd64f3af2b28b13e9956;
wire [MAX_SUM_WDTH_L-1:0]        Iccefa45795486757515d95e5908b306a;
reg                              Iab2f643f81921ed8464e1bbd9fa8c68e;
wire [MAX_SUM_WDTH_L-1:0]        Ib1357cb20f471f1670ac2448f964f8eb;
reg                              I17d7f36fdade16dbcf621fe302bd7e57;
wire [MAX_SUM_WDTH_L-1:0]        Iab953a8974a1eb619dc0f074c003b5f9;
reg                              I23afd747ecece714e32fbb896b5c022a;
wire [MAX_SUM_WDTH_L-1:0]        I6e37582849c2c98fd15ad92d22c222da;
reg                              I388528eaf83566cc56b23485a9c05962;
wire [MAX_SUM_WDTH_L-1:0]        If004de0cac6e5f7701a1fce48c6936d5;
reg                              Iea424dd9d8916c4951b8746408b8a521;
wire [MAX_SUM_WDTH_L-1:0]        Ic1efa395cc1fd2c5a1d1559fb169a5a0;
reg                              I73bbf90b625d56f663ad10f9d21d8e76;
wire [MAX_SUM_WDTH_L-1:0]        I8e96c69e7d872be23229353808c34953;
reg                              I41796b587316c600bf583edc62649bd8;
wire [MAX_SUM_WDTH_L-1:0]        Ib6aded6c73a8cc3cb964b0ae895b859e;
reg                              I7009c18515dd43d8dd2e5d1ee6779641;
wire [MAX_SUM_WDTH_L-1:0]        I939368b76d98b43826c68c7f468a5632;
reg                              I797c9cb725f88c07be28f017871d17f8;
wire [MAX_SUM_WDTH_L-1:0]        I544f6263f16cd5e0b7cf28c511a8f6e3;
reg                              I06b48093d4c9b0327c3efc6fa4ca7daf;
wire [MAX_SUM_WDTH_L-1:0]        I484545c4d2c869d79eb17f51e11070a3;
reg                              I04c734eb876aa722e84d6b9edd297978;
wire [MAX_SUM_WDTH_L-1:0]        I39289e6385a9bc378a9b8dd440249a7f;
reg                              Ifb89e7ad8ef661959d82b7c22f187243;
wire [MAX_SUM_WDTH_L-1:0]        Ie9cce5746a83479a567bbaeac6dbf497;
reg                              Id1dce2b9eafc35fa71df33ada4aac539;
wire [MAX_SUM_WDTH_L-1:0]        Ic044d7419cc43736d278c2df33b4a3cc;
reg                              Ied19cb51636bfb029ba8a2c390f97105;
wire [MAX_SUM_WDTH_L-1:0]        I6714551e8885ef5e4490673fe1b2dad1;
reg                              Ie46b71f55aef4d00168202431d47dce0;
wire [MAX_SUM_WDTH_L-1:0]        Ie9ab3c88ac62369e3d92d110165a94a8;
reg                              I8c0c1a0a35f4f7a688f516c567242d39;
wire [MAX_SUM_WDTH_L-1:0]        If38feb4f76f761dce6145731ad235d7f;
reg                              I53222c82827cab7c770e057ae91bc10e;
wire [MAX_SUM_WDTH_L-1:0]        I6359856a1843d8c8b65dc478bccb3acd;
reg                              I8015717cd36aabbf2cf4aa3a5c234690;
wire [MAX_SUM_WDTH_L-1:0]        If6f3d91c3c7a43622b9a522492cd83d3;
reg                              Ic0c13c9a929c8c46e8702cef74de8955;
wire [MAX_SUM_WDTH_L-1:0]        Id023a6298e65da1f4da3831f5136afc2;
reg                              I71d7f72d83b7410de31e09ea96adb95c;
wire [MAX_SUM_WDTH_L-1:0]        I6b24690f394792edb0d82b3b9e110851;
reg                              I1db4ea6916125702e7fb09d0f742e60a;
wire [MAX_SUM_WDTH_L-1:0]        I5b55c285f7e3e78447fee68532ab9f7f;
reg                              Idc445d3f5b3b62562b0ac83e5f17e92a;
wire [MAX_SUM_WDTH_L-1:0]        I32701d9e4b96853c53f0ab651a6a4ba2;
reg                              Iee6e52d75c093a24eb4e5e0b45feb256;
wire [MAX_SUM_WDTH_L-1:0]        I82f266e5792cdb6e7ebd264e246161f5;
reg                              Id48fe0672aa98f987162931527e9f9bc;
wire [MAX_SUM_WDTH_L-1:0]        Ibfacfe5b83819afe7fbd4bffa2d6d4e2;
reg                              Idce46f6d03376bea1ba361e8c59f8bd1;
wire [MAX_SUM_WDTH_L-1:0]        Ib8e68a77ad8b9e7cf415bee17645c3f9;
reg                              Ie79ce8adeef2c3c24a3386f054d0cf5b;
wire [MAX_SUM_WDTH_L-1:0]        I644ee0055a55f54ab3544bb532e39c61;
reg                              I0d41bef808860bde56d48792764612d5;
wire [MAX_SUM_WDTH_L-1:0]        Ic5467e42aa377c6ffd8f70673808774f;
reg                              Ib6ae81df8db1dae269437861ee11ec0d;
wire [MAX_SUM_WDTH_L-1:0]        Ic57eb4a034247a4c952d8224ea9f2bac;
reg                              I33ddee677715877c11a1df45cbfb01ac;
wire [MAX_SUM_WDTH_L-1:0]        Ia642db613c0ec1ca4e69afde7a14a839;
reg                              I433dd5092cf1851cd196feade3cfa6d8;
wire [MAX_SUM_WDTH_L-1:0]        I432aa7cb844286c442356954f8814260;
reg                              I71d3a999d88e591e102398409b3adebf;
wire [MAX_SUM_WDTH_L-1:0]        If520c1cd27f9d4bc52d0d029f693b660;
reg                              Iebecd2d19f9174d87deedc1a273e7baa;
wire [MAX_SUM_WDTH_L-1:0]        Ie87075ac979410cc11099a356966b8a2;
reg                              I168afc1863f909dbcb6a9230db9f3e00;
wire [MAX_SUM_WDTH_L-1:0]        I6fab46b1766878b26b53f352fee98223;
reg                              I1c4b29e48d0effac4839037ae5688334;
wire [MAX_SUM_WDTH_L-1:0]        Ieaf14683f40374c4531326d228cb43c3;
reg                              I431fc2e9533012c8571d8158d4777dea;
wire [MAX_SUM_WDTH_L-1:0]        I5149125aaaad943d891df6a3c2be93a0;
reg                              Ief72606c77113ae37845e4aa4a2ae5e7;
wire [MAX_SUM_WDTH_L-1:0]        I770dff588ee1f52f58bea1921cb23383;
reg                              I641539560711ff1824bd90baa0f21f96;
wire [MAX_SUM_WDTH_L-1:0]        I8f0a90e761111a613d2488285534a500;
reg                              I3ac0799861144b599995318bdade2114;
wire [MAX_SUM_WDTH_L-1:0]        I765a8825e42180a6c63f7b33703bb483;
reg                              Ie83fa8157a7cce44c2e25f46ce897dbb;
wire [MAX_SUM_WDTH_L-1:0]        I512cc8f6519aa08aee18225b56d47c9f;
reg                              I8be4711146486fea913843e497065b50;
wire [MAX_SUM_WDTH_L-1:0]        If08370fd0e8af818c6db20f43e74034d;
reg                              I65171c9ee8449407484e5c82d13c6751;
wire [MAX_SUM_WDTH_L-1:0]        I0ff382edfc8051459657ffa3899f5f73;
reg                              I7353ebf3a1cde89d2bb3fa667f7f5485;
wire [MAX_SUM_WDTH_L-1:0]        I9d2864024148337277523ef7fa2e1600;
reg                              I669d34b955d2991ebbb31c149ad1b6f8;
wire [MAX_SUM_WDTH_L-1:0]        I1c85a2d1df6749a194072eb731506bfe;
reg                              Iabb01dc9980b4879a7356712b51df0d6;
wire [MAX_SUM_WDTH_L-1:0]        I3e3ce8b4ead150a6eae2e5c701c7b598;
reg                              I373841aa2bcbad8232d54ac9035a3ef9;
wire [MAX_SUM_WDTH_L-1:0]        I45bc13ae0e0554a79c62cd9c6aa8f2a5;
reg                              Ib6124faff821158c6a2c9a9c454ab68c;
wire [MAX_SUM_WDTH_L-1:0]        I92678f5b52c9c55556ff7f17f0f607b7;
reg                              I6f7a45fe64ffeda9ed120be3a4519aea;
wire [MAX_SUM_WDTH_L-1:0]        Ib4bdc9069d0c08655f5e87f705943eda;
reg                              Id1dafb7e45b860d506e0c2c91b28142e;
wire [MAX_SUM_WDTH_L-1:0]        Idbf9094c94c931f16fba468b9dd59a25;
reg                              I5f1609647f1e71cef4ba2d605c6c8445;
wire [MAX_SUM_WDTH_L-1:0]        I1c3c4ce44610e04c5eef2fcbc2ea5114;
reg                              If17c0096ce34b88007247bf4c429d5c4;
wire [MAX_SUM_WDTH_L-1:0]        Ie84be0ae8311d906eff08f7f5b214943;
reg                              Ifc2963762403a00c4f3662b2863c991e;
wire [MAX_SUM_WDTH_L-1:0]        Ic90b98708faa8c8b75d4bd9a52c292f7;
reg                              I5fdd8e1550feaecd81b82069fe73ed7e;
wire [MAX_SUM_WDTH_L-1:0]        I8eba6f14f42701d22859fbea94bd1871;
reg                              I85654bd3a07b4329aba17d8b27777f4e;
wire [MAX_SUM_WDTH_L-1:0]        I6d83efa9f988328f487e9232bf2633a2;
reg                              Ibf2a253afde05c905d0b2404c5a808a0;
wire [MAX_SUM_WDTH_L-1:0]        Ic23e01562c8a753fd70c343297be288a;
reg                              I3ade5535a79ce83857481ac771cd8618;
wire [MAX_SUM_WDTH_L-1:0]        I5669856f88f5e2c98f64df696db76414;
reg                              I221524a69e18854f029cad30e8f94e8a;
wire [MAX_SUM_WDTH_L-1:0]        Ic3a608b850709286ea0ad2f67425d9ac;
reg                              Ied764ee7730ad129b6f62837ef50774a;
wire [MAX_SUM_WDTH_L-1:0]        I5267fa34449e6eebe891017fc32d0749;
reg                              Ic98f33c6a4613534bcc9b6bc4b4f2d17;
wire [MAX_SUM_WDTH_L-1:0]        I599d01cfe6e54d8e45d64446c446818d;
reg                              I92eb6f60c14ee9eecb01718b01ea980f;
wire [MAX_SUM_WDTH_L-1:0]        I8f94dbafaac589ac9f14b56d4556ff96;
reg                              I97e82e5f6775d1e31537b891597223bd;
wire [MAX_SUM_WDTH_L-1:0]        I754563caea429d3d0e22df5d193b84eb;
reg                              Iba1c0ebd9cefeb0dd7f690bdbbbfec58;
wire [MAX_SUM_WDTH_L-1:0]        If7f373506cac70f8ba1222db135c27e8;
reg                              I235c3a9fd3e8ea1cee762c10bc8e2c53;
wire [MAX_SUM_WDTH_L-1:0]        I69f563e7b7ad483893ac9c4684349769;
reg                              Idd474d80b50992537d6f527faf279800;
wire [MAX_SUM_WDTH_L-1:0]        Ia0a02781c674fe5d769206448d475245;
reg                              I88a89b2d938552458dab9bc34728959b;
wire [MAX_SUM_WDTH_L-1:0]        I1b7a401bc11741e6f011fb9895b5c797;
reg                              Ib105151d91678f81978495ff94b1e651;
wire [MAX_SUM_WDTH_L-1:0]        Ieb528d666fdb708279184bb59eac25d9;
reg                              I4edd64d1f1da865b1eb886e22726a033;
wire [MAX_SUM_WDTH_L-1:0]        Ic3ff7ce12c836bf0693252b9a7a7cfe8;
reg                              Ia7c9c24f8e993526e76c6915e56908c4;
wire [MAX_SUM_WDTH_L-1:0]        I19bba6a58ad3ef959b33701f82761984;
reg                              Ib0dadebad37d9ea9d01350054872863c;
wire [MAX_SUM_WDTH_L-1:0]        I8acc93b34974c1e708b0e1591f7b2d3d;
reg                              I76fd9005abd511c3c5bf6c77de8bf2f3;
wire [MAX_SUM_WDTH_L-1:0]        Ib60d4ac0fcadcdfce5a14fb92f58423f;
reg                              Ic124975d36a292816146a2fe61ab3ab9;
wire [MAX_SUM_WDTH_L-1:0]        I039f05d5be891a37e04556f1eae674d2;
reg                              I70a4926e9e6a05fa9ee51a26988862fe;
wire [MAX_SUM_WDTH_L-1:0]        Id0f75e19b94541ed5c5c352d13390d2d;
reg                              Idc5e98f6958786ccf95d39b922b42ea9;
wire [MAX_SUM_WDTH_L-1:0]        Ife1190f76c2e251704c2960c23330a48;
reg                              I8879df010bbdf6e5fc9370e2fb3289b4;
wire [MAX_SUM_WDTH_L-1:0]        Id3e0c98bff2636e216b4d3a0ffd51054;
reg                              I94a9de743d5bedbea3876de954f479bd;
wire [MAX_SUM_WDTH_L-1:0]        If4d3b31b87c0f723241d35ce7e854eba;
reg                              I17c9d8f658dd6b2916b645d103f4702a;
wire [MAX_SUM_WDTH_L-1:0]        I72369dedfe36cb22269033cc305b730c;
reg                              I384e50fa8daa639124f083dda56fac00;
wire [MAX_SUM_WDTH_L-1:0]        Iec71fe7fcebccf1ae0d10a5d187fcc44;
reg                              Ie165d0729542c81ca89f45d15e0afd3d;
wire [MAX_SUM_WDTH_L-1:0]        Ie11da10808c4ca84f399535df6261307;
reg                              Ie8e29053f122a9247b0dec291c6ef4f3;
wire [MAX_SUM_WDTH_L-1:0]        I280fa9d114e227cd649bf0e55e845651;
reg                              I453dd7d7c0a2f003f0b67e909630d641;
wire [MAX_SUM_WDTH_L-1:0]        I94c4e11670b4233fa072517a8f19c901;
reg                              I5707d30ca29842b6a96cfaeb44ac6668;
wire [MAX_SUM_WDTH_L-1:0]        I4dca2dd40a7127ce44f83b430a34c738;
reg                              I3fbd40faa4c3b78b547b8348c466fd1f;
wire [MAX_SUM_WDTH_L-1:0]        I1a24e98165afa62bd14986911a36fb6e;
reg                              I9a403c511fe2d44472ab319a9477199c;
wire [MAX_SUM_WDTH_L-1:0]        Ife1164cad7cda4aa9a08d94dfe86add6;
reg                              I9db50007841762c9a10f6b7e9d40f858;
wire [MAX_SUM_WDTH_L-1:0]        I8d8d95ff26f33f69a182b32ccde23905;
reg                              I89c5af1a6176cefa1f77ee69996473cb;
wire [MAX_SUM_WDTH_L-1:0]        I2508854bcbab37bd09c9465c377c06aa;
reg                              I5ede62333e0f7ddc5446b653ba9a2382;
wire [MAX_SUM_WDTH_L-1:0]        I140078292f7209eccacd53a8bab18016;
reg                              I69d82ab774d52c219509e993e7cc4deb;
wire [MAX_SUM_WDTH_L-1:0]        I141fb1cbe09f9abe282cffd4de815d25;
reg                              I0eaa22f5eca8f33dd254fe241017a098;
wire [MAX_SUM_WDTH_L-1:0]        If79d1d378f7c6fd29fc3335ec5f5c51d;
reg                              I570c036d0237c53bb069c52d621e539e;
wire [MAX_SUM_WDTH_L-1:0]        I4a41999cea9357a85c73a0af509eeac9;
reg                              I9d7614d286377329eb3999213889b707;
wire [MAX_SUM_WDTH_L-1:0]        I8e517c401d62dbb10dcc96ab536f6afb;
reg                              I3eab1582cc42db0ac7739386cce2a712;
wire [MAX_SUM_WDTH_L-1:0]        I8ad3627f171eadcc960a688ac0afcbc0;
reg                              Ie4827dc0983c1a63053c08de6e36d375;
wire [MAX_SUM_WDTH_L-1:0]        I85c4d3d6c8408c6f38741257ed177ca6;
reg                              I2eed3d32a27d51036e17c4a21382b4c1;
wire [MAX_SUM_WDTH_L-1:0]        Id66c47fd69c175a4393e975a269cf053;
reg                              Ie039ab562e9cf90289047b5425186123;
wire [MAX_SUM_WDTH_L-1:0]        I37dca40506d61bdeab1255ed4892ca20;
reg                              Iefbdf686d9452a62cb99cf023a4d9fe7;
wire [MAX_SUM_WDTH_L-1:0]        I340c98b886123c541a1b8d9fc8a6d48c;
reg                              Idc5dd6caa4ed17a63746d30d381a944e;
wire [MAX_SUM_WDTH_L-1:0]        I2dc64c3b06588542b027f997437bee63;
reg                              I17086dc5193aa55e5c6f56ecd365cc00;
wire [MAX_SUM_WDTH_L-1:0]        Id92a37c091100e9df08e24498ecb4022;
reg                              Ib2fe0f68044c11f879e512a200f8099e;
wire [MAX_SUM_WDTH_L-1:0]        I74a4b9365391fd20c34588002ad40547;
reg                              I768720af835b02a8dab376ef23d17a15;
wire [MAX_SUM_WDTH_L-1:0]        I461195b7ae78743e09ee50486ad6ebe5;
reg                              I1d98943b01a6a2d8c4db18b98dd62f5c;
wire [MAX_SUM_WDTH_L-1:0]        I356d747600182675699a2d2634d4c5ce;
reg                              Id3b089fb6edd5bcfdbca142fddd5ff89;
wire [MAX_SUM_WDTH_L-1:0]        I87d6a5d30c3e4202cf51f33c7a770c51;
reg                              I5196382b75d16892d550f17893de15ec;
wire [MAX_SUM_WDTH_L-1:0]        I960768a84aec9d5b8bc7c1c523024a25;
reg                              I6387919f2426c283e2d70e471cda54a6;
wire [MAX_SUM_WDTH_L-1:0]        I09b5273bb15d48a7fd78559930fa6d1c;
reg                              I3b84dad6d0dd8730312b3e20c6d5a2a8;
wire [MAX_SUM_WDTH_L-1:0]        I5814a85c45fd0f7be21ed325235fe4b7;
reg                              I2a4bbedf880a9a7b4e1bf946f9f96c0e;
wire [MAX_SUM_WDTH_L-1:0]        Ib06b60cf9933dd8952206c5f3ccced8e;
reg                              I49d35ec6369de10afb15be8e0cf135c3;
wire [MAX_SUM_WDTH_L-1:0]        I67347c413b5efd8ff9e0d5bc7ab2a047;
reg                              Ic3ba4531855366e9a060cec1c7694844;
wire [MAX_SUM_WDTH_L-1:0]        I72b1bb104bf2843f161448baf7aab44b;
reg                              I4dbabfd592b74aef93b819163130ef5e;
wire [MAX_SUM_WDTH_L-1:0]        Ib23d889edb5a6d9f27de977d3b1a2616;
reg                              I9ece87047aec25abc02a5eea72f0e647;
wire [MAX_SUM_WDTH_L-1:0]        Ifaff9dd032cf96487be819c59b03000a;
reg                              I3ed6426fbdba8aaf1c948cca7442b3a6;
wire [MAX_SUM_WDTH_L-1:0]        I028ce03be0618b816e0ecdf43d4cd6e6;
reg                              I24075f37c6bbd90c83370de1a2e58af2;
wire [MAX_SUM_WDTH_L-1:0]        I6ae2523095237282533e0b5f1c26b488;
reg                              I3175159add7b814df637c2db8feb43f6;
wire [MAX_SUM_WDTH_L-1:0]        I5aba6218461e8d571be03a3ef041ebaa;
reg                              I0a569f6536789efb7ad2377c11842830;
wire [MAX_SUM_WDTH_L-1:0]        I6ca8a1fa2c72b1c61d11dc7d1ba5f37b;
reg                              Iae6ed7748692f2edf1aa9d73380075f0;
wire [MAX_SUM_WDTH_L-1:0]        I3ec5819176ad4b0895a9118d90ab22b5;
reg                              Ib4ae1cedd09d72c235765a6cd7e91366;
wire [MAX_SUM_WDTH_L-1:0]        I49b64469d298012dbb131d879bff38d6;
reg                              Ie2d946edaddd3c87f328e861f3e72c0a;
wire [MAX_SUM_WDTH_L-1:0]        I95361d5f524ccb9feb42811af5c482e2;
reg                              Id6b508145cd21ba088ab8fda34577c35;
wire [MAX_SUM_WDTH_L-1:0]        I9c4b34b5fb1d59c132bcaeb6258675df;
reg                              Ifa6e3541f5e12bf9677ffc51d0392749;
wire [MAX_SUM_WDTH_L-1:0]        I613d4b1e3b9e812b785c9cf14fefdfe6;
reg                              I21e72a7e5870151c3247d15121e5fb4f;
wire [MAX_SUM_WDTH_L-1:0]        I848ed394bd4f0b199d11c0ff458394a7;
reg                              Iba283e99a57d0a3b78ad2e309c316b65;
wire [MAX_SUM_WDTH_L-1:0]        Ie65a0634454381e24bb3223a333e3ad0;
reg                              Ifba3e46933049cb093d2c1809f3a8a3e;
wire [MAX_SUM_WDTH_L-1:0]        Iad166146f7df5e8068fc6efe4d3e4141;
reg                              I4af3e2bf2ebc913ac902b48da672c5b6;
wire [MAX_SUM_WDTH_L-1:0]        I63e45abd4d27219bddcef06108b72021;
reg                              Ifbadefd3a7ab50719a703400ddd742c6;
wire [MAX_SUM_WDTH_L-1:0]        Id1bacd13718f7c29c26b63c239d04dd8;
reg                              If2042aede3390bd208a281f0380c95a4;
wire [MAX_SUM_WDTH_L-1:0]        Ia3104c69fb4f7abfb5efa3874169a7ad;
reg                              I19b73c5c93a71e90f620572f23f0e6d2;
wire [MAX_SUM_WDTH_L-1:0]        Ie1b7257c99831ec5864f65958ecf14fb;
reg                              I4b99891bed4f5c149cd4a5b4f1dde0f0;
wire [MAX_SUM_WDTH_L-1:0]        I4accbad1b451ed2b622e15ef9ae16d13;
reg                              I3472ee8c06644490252e606b62bf9bd5;
wire [MAX_SUM_WDTH_L-1:0]        I5ce8b2f633011e89356243a1a71edeb6;
reg                              Idb1efe99b5d7fd567a7f82cfd52f7eb8;
wire [MAX_SUM_WDTH_L-1:0]        I3e5139f24e3d082eb31b0e61ea9fa1aa;
reg                              I24f82a3f2c0e8df486fe495dd95cf8bc;
wire [MAX_SUM_WDTH_L-1:0]        I61cc8a0f49e393721a62a776e4793deb;
reg                              I83ecf12f3b38fc14c3b75e47b71ecc09;
wire [MAX_SUM_WDTH_L-1:0]        Ie631e40caade823a196370fc3358f042;
reg                              I74cbc0ec3bb682e0f927890eef8d7a58;
wire [MAX_SUM_WDTH_L-1:0]        I4c971e714427664c59c6371e14781bae;
reg                              I989dda9add29306d7b3c0f376822763a;
wire [MAX_SUM_WDTH_L-1:0]        I36ca732e811d67cd742d24fd4cae887b;
reg                              Ibc929201e2eeb3e61cc8f0acbade497a;
wire [MAX_SUM_WDTH_L-1:0]        I354fdd241d5d07f0d8380fe8924e0a8c;
reg                              Ib0dfbbbca2d3d264065f73b4241caed5;
wire [MAX_SUM_WDTH_L-1:0]        Id38b705f5d2863a020a475ffffc8afd6;
reg                              I339786aa60d4c71d12c65db27ac420fe;
wire [MAX_SUM_WDTH_L-1:0]        Id6e5d67e7bb7c4b999459374ea80459a;
reg                              I3ade020bbdf8f954821f737439513043;
wire [MAX_SUM_WDTH_L-1:0]        I05341013abd4206eb66fcddfd63bfe26;
reg                              Ia50526cd3a3174bebc5a7a0889fda661;
wire [MAX_SUM_WDTH_L-1:0]        I15da71a21f5842cb65b543d9bc3e267b;
reg                              Ie9f37dba0791359bc426a73639ce33ad;
wire [MAX_SUM_WDTH_L-1:0]        Iccf255fb3422c558465e45226068a16d;
reg                              I9518532a8617fc8290eb6a5e981dea94;
wire [MAX_SUM_WDTH_L-1:0]        I1c2674b2e6b269ed539827412c5199a5;
reg                              If66524125bfde5aa48ac70c4e448b38f;
wire [MAX_SUM_WDTH_L-1:0]        I6a3f405bb4a0c4448d9b9d3dd95d036c;
reg                              Ic3ec6375998b05a3e48f6c5fe7b3910b;
wire [MAX_SUM_WDTH_L-1:0]        Ib528bb7a64cce4f694081d151fa6fa86;
reg                              I0ac421af6e311b6005c3e02e93ff94ce;
wire [MAX_SUM_WDTH_L-1:0]        Iaa40bd3abf668a21e0f87c7bda7b3f69;
reg                              Ib9db80f43718305a8a8774d8d80c86c9;
wire [MAX_SUM_WDTH_L-1:0]        I919d36a7f6ad42c4bbc23222beb73106;
reg                              I3b775b06b5d78fcd7373c966a62f44ad;
wire [MAX_SUM_WDTH_L-1:0]        I648d2a279dd1f587b1e45eeb35f2fa90;
reg                              If2372a5956f21f97eeb9c76281b6675e;
wire [MAX_SUM_WDTH_L-1:0]        I194a64bef92ecf6714141eaa5d41c9d4;
reg                              I7b32c2b108e24750e2a24785668af3ea;
wire [MAX_SUM_WDTH_L-1:0]        Id332e7f482524adeac7f7cdafcf5ca46;
reg                              I8ec99197a7d823f5745d382c10161430;
wire [MAX_SUM_WDTH_L-1:0]        I226383d68f89db716cfd8d08b837865a;
reg                              Ib895fec0b3756932b85962c1d129a03e;
wire [MAX_SUM_WDTH_L-1:0]        I2bdf5d319ba9089a4da34b108f5c5ae5;
reg                              I76aab345d13c6678fe37a4a7133cfd7d;
wire [MAX_SUM_WDTH_L-1:0]        Ia91800792941ec7cc60415c3f844e4ed;
reg                              Ib4f368fa3d3ec11d9ffb2ae9a2ae6310;
wire [MAX_SUM_WDTH_L-1:0]        Id7c507d96098ee7a955af8a48ee5d72a;
reg                              Idd0f3cfc5599481c954a2bfe69f044e5;
wire [MAX_SUM_WDTH_L-1:0]        Ie15e4c1bcdb0e18085d4b320ac6a925c;
reg                              Ie624c4dad5036a25ca314b94cf3c4b95;
wire [MAX_SUM_WDTH_L-1:0]        I5485d9edcafc6202f6e5f0969979802f;
reg                              Ibf4b3caa5655cfb6663f9b7e2383bbbf;
wire [MAX_SUM_WDTH_L-1:0]        I7fe364f9f537cbef782e7007848a1c10;
reg                              I049d1c09c15def12ba7bae95fc1c3d55;
wire [MAX_SUM_WDTH_L-1:0]        I52dcf5bace9cadcf8a895aaa6a8c1da8;
reg                              Ide06ba186ddb179b489ba6e3e209e3e8;
wire [MAX_SUM_WDTH_L-1:0]        I13a9eec6175e695ab8bc4516cf57d6ec;
reg                              I1b78785ebe2e7f77a3125a6334c4dc54;
wire [MAX_SUM_WDTH_L-1:0]        Iee73a7c685a4cee03f33d3ef379b1c8a;
reg                              Ie79c93f1703121713fb9401617f349a8;
wire [MAX_SUM_WDTH_L-1:0]        I740dc91716e3906ad078e2c7cc3c925a;
reg                              Icf25f076eec2bf81c899c66f6cfbebc0;
wire [MAX_SUM_WDTH_L-1:0]        I514d2dc697e9b39ba027c418a6df6cb9;
reg                              Ic5c837a0556d1cb66edbf0294d08283a;
wire [MAX_SUM_WDTH_L-1:0]        I782726e317a2aada9e755bcbc4b0d3fa;
reg                              I51ff4bda38746682e3cd4c68118c3216;
wire [MAX_SUM_WDTH_L-1:0]        I11eb26cf0f0b3a334e8f7317bf8d9eb0;
reg                              I1c074a53e6c0f2467bcdd7c952f51670;
wire [MAX_SUM_WDTH_L-1:0]        I26cb63ba20245b2c332b09e25c4409aa;
reg                              I37c49c5a2af240496f5a5706b0d42ea6;
wire [MAX_SUM_WDTH_L-1:0]        Idd7691d31f8d0c09ee988116d574ec59;
reg                              Ia94c439131e1df5c95fc8ad3cfdba473;
wire [MAX_SUM_WDTH_L-1:0]        Iecc02842a2d2b9b9e8187f2d39e62e05;
reg                              I723a6fee3b2496f23c48b3584f8bf9ce;
wire [MAX_SUM_WDTH_L-1:0]        I5551342f1751fc64f32744a46b9649be;
reg                              I648b62fa0bc2185c1756ee531e8e34de;
wire [MAX_SUM_WDTH_L-1:0]        Iff7c29299f005c1cd5a16b64601e727e;
reg                              Ife631f9a3c4c64a3d92aa9586ae75f3c;
wire [MAX_SUM_WDTH_L-1:0]        I17a5446e942bcc1dc2c96930e0a87a70;
reg                              Iaac1d82f0846fce1bd88ebf8e60300ac;
wire [MAX_SUM_WDTH_L-1:0]        I719b67f84e07e90dfd29a8cd5d94cf39;
reg                              I48cd09f035f668536cd288a23010b07b;
wire [MAX_SUM_WDTH_L-1:0]        I2c835dfb3596b8bf057a7cc21122c81f;
reg                              I119b2e5c2fea5338244c4019884af26f;
wire [MAX_SUM_WDTH_L-1:0]        Ib71b3d357c98dcdfae5c777ca3082275;
reg                              I2bd34b2fd12f12bc301fd0d5d69c0fb6;
wire [MAX_SUM_WDTH_L-1:0]        I086bf19f620c8a8f6888e775cb1ed7f4;
reg                              Ib715b1e0061b84ce614a30d961a83e7e;
wire [MAX_SUM_WDTH_L-1:0]        I802c554d5b04af6b949677819a4966ed;
reg                              Ief8c2838abac83370fd7ec25c06d509b;
wire [MAX_SUM_WDTH_L-1:0]        Iceefb06cb3715e1b41e6f7d89420e5ba;
reg                              I561d79eb079915c0b1732cbddb119c2d;
wire [MAX_SUM_WDTH_L-1:0]        I56948bc48c0220893d68004615a6ebaa;
reg                              I8bb75bf828d5ef337fa6a965808e4638;
wire [MAX_SUM_WDTH_L-1:0]        Iec1368f034655d61354ab5b5e94d7d89;
reg                              I11ba339c8250d07b497c88a39a6df1ac;
wire [MAX_SUM_WDTH_L-1:0]        I1e43c0aeeb8a2461d208eba24967af30;
reg                              I173aa69cf52114e223ac1410d90b4bfe;
wire [MAX_SUM_WDTH_L-1:0]        Ia6eb85b127cf9c1a437611556296b967;
reg                              Ia4e89e99acb95f4183474b94798ca35d;
wire [MAX_SUM_WDTH_L-1:0]        Ieba89aa901e61218074af53a2484a74b;
reg                              If4c36727ab1c29bf78f72e8acfc00d7c;
wire [MAX_SUM_WDTH_L-1:0]        I8b3b875c6c07bd97ba598a5139156fa4;
reg                              I6426943b4ab66f17c2b7b399ccc7a6a9;
wire [MAX_SUM_WDTH_L-1:0]        I7b33ddad346077928620344542b9481e;
reg                              Iddcffa815489773b3688fd68dba18bd8;
wire [MAX_SUM_WDTH_L-1:0]        I11d967a5c5d14c88b5587d4cfed1d05f;
reg                              Id00642563679fa9a6696f8e7bbdf6576;
wire [MAX_SUM_WDTH_L-1:0]        I27458d76b3ac6520fb379405c6b2956f;
reg                              Ifda1c55899cd3506853cc82b450b3936;
wire [MAX_SUM_WDTH_L-1:0]        I2525111a2fb5f10d64bbd16e148653b8;
reg                              Ib5d1a7cdbcba0b654c12063d4f1768e1;
wire [MAX_SUM_WDTH_L-1:0]        I7b7cbcd1c6d2a2eeaaff474536a69eed;
reg                              I5e8ed024e2f2548bb375a2ecf1918a5f;
wire [MAX_SUM_WDTH_L-1:0]        Id2a7f0781d18dccc7c4e0b383b7cddfa;
reg                              Id25deba967318f049de8163e67262f4b;
wire [MAX_SUM_WDTH_L-1:0]        If8bc141d98ebe1be7fa81cde5c65868e;
reg                              I925f6b549a25cdc8f85152eb21ea3b58;
wire [MAX_SUM_WDTH_L-1:0]        I8645e1326c66f5efef4b9c923599d1a3;
reg                              I9b49e1acb81ef5b088b808d2e4ce9954;
wire [MAX_SUM_WDTH_L-1:0]        I0426ef66185128dd1ef4dbb68dcda585;
reg                              I6386a4dd26e7c36165dc265b3a2c93cf;
wire [MAX_SUM_WDTH_L-1:0]        Iddd954df5bae9b4240e0512f746669a9;
reg                              Ia20709f08cfff3a51d4af1e81d640400;
wire [MAX_SUM_WDTH_L-1:0]        I29e940970d87e8e09b26ab1b0b8f2286;
reg                              I1ff042bdb52aac5d69791e96e2f9706c;
wire [MAX_SUM_WDTH_L-1:0]        I488f6d9676aa85a55d030bf12e8997a7;
reg                              Iaa2cbf59f6f61198b4fcf5a741cd5bc8;
wire [MAX_SUM_WDTH_L-1:0]        I99d761b75ade1fb2e8afbb1a77752609;
reg                              I01c94743a11042e75638ba6618356203;
wire [MAX_SUM_WDTH_L-1:0]        Iac4e3d20178049f9c59abf374752dccc;
reg                              I0a0340a0e52145f3597accfe4a4e8624;
wire [MAX_SUM_WDTH_L-1:0]        I618d33f26badabfa578908903a613bce;
reg                              I3bb4d24caaa0882a75125e466070f0b1;
wire [MAX_SUM_WDTH_L-1:0]        I822d7973afe090b2764335f1b72dfd0e;
reg                              I44ead0ab5ccc53226fccc03024643771;
wire [MAX_SUM_WDTH_L-1:0]        I12c1035353e553b3b6a13bb174ce6020;
reg                              Iaded125f7fd5c833e7206dd7071069be;
wire [MAX_SUM_WDTH_L-1:0]        Ia6d61947d36fc128c689808c82db80f6;
reg                              I373be7c3f9511a2906584e33e5048abf;
wire [MAX_SUM_WDTH_L-1:0]        Ie9b042f686381739b9ff219041f1e0ce;
reg                              Ie0b5f51835ebdb508a596eeebf0e4847;
wire [MAX_SUM_WDTH_L-1:0]        I0c4268c01aed70ce4fc71531bf4bb862;
reg                              Iddb75e0197b9a76b36a59ac2a7ccdf3a;
wire [MAX_SUM_WDTH_L-1:0]        Ia34e42f8de91fa4861b0c6cac5dcfc29;
reg                              I08c03198b9599b2f4590e3022e398f7c;
wire [MAX_SUM_WDTH_L-1:0]        Ib7c5850b4f7cc77be2048d114a2128d9;
reg                              Ia4f3cff223e24815ee1d86bf41756f06;
wire [MAX_SUM_WDTH_L-1:0]        I32bb50faa2b246b2d3b462a79be597c5;
reg                              I56592e1452c4b559af19465b30230ec0;
wire [MAX_SUM_WDTH_L-1:0]        Idc6d40a49f05c5422758cee50f787eb1;
reg                              I213ce488e5345fa405a9c5df297d6f74;
wire [MAX_SUM_WDTH_L-1:0]        Ide1d7dc22a4b271ef764df14ac22366a;
reg                              Iefac1e428116a797c2c0803410ac5601;
wire [MAX_SUM_WDTH_L-1:0]        I7ace6778ac86b3e05939a3fcc716136f;
reg                              I8b419d5827e5b1af9649d602401c189a;
wire [MAX_SUM_WDTH_L-1:0]        I044e01e8d2df46e03f00a0af2beb0bf5;
reg                              Ie989550c9101de382056dd60d5da0e01;
wire [MAX_SUM_WDTH_L-1:0]        I45a7ddcda2662e36b7617dfe64514346;
reg                              I259010e323e1e8dcd9dd719091131f6c;
wire [MAX_SUM_WDTH_L-1:0]        Idada779a1ac7b844867571d77054b657;
reg                              I389ac86954fd70464c9550e3fed4ed33;
wire [MAX_SUM_WDTH_L-1:0]        Ieeba01b18a244ab8c0ac263c138fabcc;
reg                              I77371f0e55b4684d1af196ed52d3d997;
wire [MAX_SUM_WDTH_L-1:0]        Ie4c9797a955778694dd8615219cb51e7;
reg                              I5a21996f5724a2a49fcf8e928c01b062;
wire [MAX_SUM_WDTH_L-1:0]        I28a5ed4c239e64c76bb6e566b50cfd23;
reg                              Id46108963921efa50aff64d4dd7d1701;
wire [MAX_SUM_WDTH_L-1:0]        I79a705ee1e414fe4a5fb14e9b3ce9597;
reg                              I8da50e5093acefb6f809aed64564a53e;
wire [MAX_SUM_WDTH_L-1:0]        I04f90a907f10a7fa1ae3591b48094d5c;
reg                              I03b0694777d0160a83cbc82ac1397736;
wire [MAX_SUM_WDTH_L-1:0]        I31d25b1b49e65216e90b39aa27acd6be;
reg                              I85c2bffb93569d9fe1b1bcb10b98bcac;
wire [MAX_SUM_WDTH_L-1:0]        I1f6540c5f037d861dee2c0091cba01ec;
reg                              Id00274c88b93867a80606343add1cdab;
wire [MAX_SUM_WDTH_L-1:0]        I9632bb500b7faaaaeb649d74c21cbe8c;
reg                              I61e829cbf7d6c0ef8ddc11677981e2cf;
wire [MAX_SUM_WDTH_L-1:0]        Idd0217a35c3adc8abc7bb581a5df7a2d;
reg                              I9e8ae2aed048068b01b3bd46f30baae8;
wire [MAX_SUM_WDTH_L-1:0]        Ic05b46168884322644db4e331d37d759;
reg                              I7dab71adbe62687846fc027d2789451d;
wire [MAX_SUM_WDTH_L-1:0]        I53c88dc237bb2cd02d50fd7f0a168a48;
reg                              If1295608bd218ed60922a0b95bf1d098;
wire [MAX_SUM_WDTH_L-1:0]        I7450d4ab3ef0227e93a02bfd620d047b;
reg                              Idf04e08c120ed116af14a62659675b44;
wire [MAX_SUM_WDTH_L-1:0]        I2b16e5b4e279bb29c3c675b72083e5fe;
reg                              Ieb7614ad1b1bfed3e2b0089a72fe214a;
wire [MAX_SUM_WDTH_L-1:0]        I70c92e8ada46476d15ef4b3c620d2601;
reg                              I589062eca318b25dfe5735da455b6fe1;
wire [MAX_SUM_WDTH_L-1:0]        Ib193b07804d6d5f111b06bda487bfa5f;
reg                              If3db87afb3ea184c9e4020c5e45cb161;
wire [MAX_SUM_WDTH_L-1:0]        I885433b0ab16c6d87abe45af13c9e529;
reg                              Ia14bc1fcd5bbdcb60b8e68298f7d716a;
wire [MAX_SUM_WDTH_L-1:0]        I198c055930cb89d0390c336eda8fed4f;
reg                              I268b60cb371b3d46dc3f8b0009f541b1;
wire [MAX_SUM_WDTH_L-1:0]        I688a2c72e69b217d2673e8da75146a83;
reg                              If2cd93b57cd1c2b91ee7a73a97dd19f2;
wire [MAX_SUM_WDTH_L-1:0]        I3b6fde4ed14cd68af1468ae1d4cc1a22;
reg                              Id81305359a07db527e49fda05cd2784f;
wire [MAX_SUM_WDTH_L-1:0]        I5d3df1e7563630311f56143ee6d97a8e;
reg                              Id8292eca087c1a17dc8b5a572a76f21f;
wire [MAX_SUM_WDTH_L-1:0]        I90a7ea789d3bf7f9126c786474a56da0;
reg                              Iddb19725b093506e5e521d8d68dcb8e1;
wire [MAX_SUM_WDTH_L-1:0]        I5029424c9d9fe923eeb858b1e62cd758;
reg                              I0b573d3a86a3111451da661e46384876;
wire [MAX_SUM_WDTH_L-1:0]        I1e805c70d50c2765b4a03ad2982dc421;
reg                              I0ff479e61d1a0cede88ebffb073c60be;
wire [MAX_SUM_WDTH_L-1:0]        Iba58175a7fd5c5da650222193caff0b3;
reg                              Icd6f8f5df6b4ca4c81855e974db76526;
wire [MAX_SUM_WDTH_L-1:0]        I7401a0501ba69c5559fbf00c77e58dc5;
reg                              I7ce064a756dad56d37684d5d7d168047;
wire [MAX_SUM_WDTH_L-1:0]        Idd9f7ea657ea9cdcb45a7e4b573b9d50;
reg                              Ied2ea62cfb21602645babc36e27b8218;
wire [MAX_SUM_WDTH_L-1:0]        I53f275395dd6be17961a5edc3e8da7f2;
reg                              I79b85da6e5ce0b02ebd1619115c98e24;
wire [MAX_SUM_WDTH_L-1:0]        Icab010d78cd66b02e089c74f04bf4e75;
reg                              I8e1ddd7e4185c28caa71d30bc28138f3;
wire [MAX_SUM_WDTH_L-1:0]        I376a48b7e0195a5aacc76a0ad8bd14b2;
reg                              Iab0bff1633e2f3ea0bfbc291f3ab5d29;
wire [MAX_SUM_WDTH_L-1:0]        I241622b0367dde514f96ece55c8c3964;
reg                              I5f0751fceaa008feba5c6867ced453dc;
wire [MAX_SUM_WDTH_L-1:0]        If94a1abfb972f63629d07e64dc23863c;
reg                              I9f6751c15237c20b0cf2175575195ea7;
wire [MAX_SUM_WDTH_L-1:0]        I07b9b1f4fa01b16cc69356057d3b6154;
reg                              I6ea50be10bc990a1206cdc9e28e0c4c2;
wire [MAX_SUM_WDTH_L-1:0]        I2288a6ad3b748b716249f4adc42d52c4;
reg                              I43c2fab87f70ea883321ab82de85f133;
wire [MAX_SUM_WDTH_L-1:0]        I022df337bcc05ac5648b8ae2e42f3a76;
reg                              I1af02ed6cf00d4cb0704b5e44c83bfa3;
wire [MAX_SUM_WDTH_L-1:0]        I60d9a7f95fb8623753002ecaf9a4efcc;
reg                              Ib71611afdd0381cc1884f5ddbbae1acc;
wire [MAX_SUM_WDTH_L-1:0]        I23a74ea5e7174d95e6d16a5e85ac236b;
reg                              I38fc49afce0298846ae8ed63ae715e81;
wire [MAX_SUM_WDTH_L-1:0]        Ie697d28d757df82b3901564bda43251c;
reg                              Iddc3e44d83e8253e5129b6cbf5082df7;
wire [MAX_SUM_WDTH_L-1:0]        I8572aedc94f7243ce5eacb332c81eae2;
reg                              I975a87bdda30c5b6be8d2f0e4b107450;
wire [MAX_SUM_WDTH_L-1:0]        I6734123aaf6320da75638b212812732f;
reg                              I582bd96afa764ded148202f738b7a1df;
wire [MAX_SUM_WDTH_L-1:0]        I7f6dc6f0f403c58f9aaaa70c2383a666;
reg                              I6fb88d97bc9ed37a06b729020a1df140;
wire [MAX_SUM_WDTH_L-1:0]        I66391978843c39b6acbdb4847a01050a;
reg                              I1500943c4a550e78fc169437b0a663b7;
wire [MAX_SUM_WDTH_L-1:0]        I4f756e4125c8af5c412944b273e01cb0;
reg                              I0b83f4ef8ba9badb27e81b32765ec5b6;
wire [MAX_SUM_WDTH_L-1:0]        Id2c9f7ac95de07148c54803f69347f56;
reg                              I2c420acf428e44cdd9ca9998e276f258;
wire [MAX_SUM_WDTH_L-1:0]        I5061e13a179d27e1ba5f89ce8ee0fd4a;
reg                              Ic7b6dae3017b55dd3cd27423d5f1b0ec;
wire [MAX_SUM_WDTH_L-1:0]        I0f7c32fc1548fb49b8041f55c157498a;
reg                              I4a91a7c9b2a0f3552b8f2ef4e2398be2;
wire [MAX_SUM_WDTH_L-1:0]        I89ffab735ee30423c82e079ed98216c5;
reg                              I99ff29c7ba68b5d0819f1e1bead51287;
wire [MAX_SUM_WDTH_L-1:0]        I9494921d8487ee0b314f75cf0380fd2f;
reg                              If06b00be0356a2be5074d958ddcdb2f9;
wire [MAX_SUM_WDTH_L-1:0]        If2b3e7d1541cbd8ffc2b4cfc3ad13a57;
reg                              I604283449f13c7b225ea03f99f2e296a;
wire [MAX_SUM_WDTH_L-1:0]        Idf3d79da44f2d686f5bd43c3c1427430;
reg                              I2b600e5f5c146ee97c4044c08e1f5ad5;
wire [MAX_SUM_WDTH_L-1:0]        If8125ad3c9e7f0a2b84106064d320996;
reg                              I9fe16403fc21bb1159a5e0305fd1ef69;
wire [MAX_SUM_WDTH_L-1:0]        Ic9018b88fa91fb638bbab0613795ae13;
reg                              Iabdb9374e5caee281c25b003624b2c4e;
wire [MAX_SUM_WDTH_L-1:0]        Iad4ea0196eb32f9a152c9e6fe5059e46;
reg                              Ibd12036702fe60b57354b3aac921559d;
wire [MAX_SUM_WDTH_L-1:0]        Ia8ff29ed728e7f2ae4213f00328b495d;
reg                              Ib1639811de6eb1c38257800c201fb704;
wire [MAX_SUM_WDTH_L-1:0]        I70717726200ec02929f679ef05496455;
reg                              If926d98f659e8fe4bbf36ad2c5c852c5;
wire [MAX_SUM_WDTH_L-1:0]        Iaf1e4c7dae6ad89567836877c08f57d2;
reg                              I211f8d7f97ebb8eb3e50313513abfb1b;
wire [MAX_SUM_WDTH_L-1:0]        Icd09aa81e9b43528af73e23b2f0f80cb;
reg                              I304ac9f96945546cdf1b6f1fa7136731;
wire [MAX_SUM_WDTH_L-1:0]        I6ebb2b94f0f80425f8401ae823d92a1d;
reg                              I7a9800418bd5c195fc47a72370680b56;
wire [MAX_SUM_WDTH_L-1:0]        I4a2c3204a6a9936d4a215b46c0ffd045;
reg                              I5f6a61c9f0c67510e148e596f553a4d6;
wire [MAX_SUM_WDTH_L-1:0]        Ib02c0694762c4815448b2c8d3df767c2;
reg                              I8e313ceb21359bcc44114ab217b1c394;
wire [MAX_SUM_WDTH_L-1:0]        I98cee6efbbe565d3a4de16703189782f;
reg                              I4c9518755c33d725221ad79ee6badba9;
wire [MAX_SUM_WDTH_L-1:0]        Ibf981c01a9d44cbea3c6d8ead92bc2ab;
reg                              I3c3cffec9f47c9979cb9503f222f370c;
wire [MAX_SUM_WDTH_L-1:0]        I864c33e8ea204d20a9baef4584f22d4e;
reg                              I68d6769541fdc3df321e192f645c667f;
wire [MAX_SUM_WDTH_L-1:0]        I6ad3228e0e2e1f19648d73e83ba5a229;
reg                              Ided55428cbb77f454c2607ac783d7548;
wire [MAX_SUM_WDTH_L-1:0]        Ie099210a99a4899c53baf39559592690;
reg                              Ifd3d4f3e2a388b3c70e7704d6351e0ba;
wire [MAX_SUM_WDTH_L-1:0]        Ieeec71d9df4613555fade2ced7b3baf1;
reg                              I17d32f292758416fe02527dfd938fa0d;
wire [MAX_SUM_WDTH_L-1:0]        I4931884e3544af182bcda9061091a42d;
reg                              I9ce3942aba354c1fd7d6b9a39c994d7b;
wire [MAX_SUM_WDTH_L-1:0]        Ib3fb10da528d450251764a9b9ede0dba;
reg                              I2c6c6041c9c69c84f4d64af6458955f5;
wire [MAX_SUM_WDTH_L-1:0]        Icdc9e676957b2223d60c413331fa982f;
reg                              I830a4fffe1244e071eb82c28ddc4a308;
wire [MAX_SUM_WDTH_L-1:0]        I381f6051282c062ccf53866830344cd4;
reg                              Ifad8e46fc3844bbfaf434a14f6b5869d;
wire [MAX_SUM_WDTH_L-1:0]        Icfc21935c007fbbceb2a67ebe1a68a0b;
reg                              I10a6c6a8fdb0003de1f360c148777d0f;
wire [MAX_SUM_WDTH_L-1:0]        I120d597a80158374726e064fb0f099fb;
reg                              I4cde586fc28f8d03fc9934d56f7ff7b8;
wire [MAX_SUM_WDTH_L-1:0]        I2520aa556aadf851f58f0b1820498730;
reg                              Ib83a067fb08e118dcf794902beef9405;
wire [MAX_SUM_WDTH_L-1:0]        I6203f49a08107f7185ebadeecf2c16b0;
reg                              I358cf9609272a4562423a85f9b2f56bf;
wire [MAX_SUM_WDTH_L-1:0]        Ia706fb593b63cebbee0321c154cb859b;
reg                              Ic1e9d9113150ad57954c0e369259dc62;
wire [MAX_SUM_WDTH_L-1:0]        Ia4b5f2b07556629673fc6576bc49a5dc;
reg                              If7fe3f5ccbb5b279e41fd183c8ff3974;
wire [MAX_SUM_WDTH_L-1:0]        Ic532c6b85b156f821e0742f47239a65c;

wire                             conv_Sgntin_row_00000_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00000_00000;
reg                              sign_qin_00000_00000;
wire                             conv_Sgntin_row_00000_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00000_00001;
reg                              sign_qin_00000_00001;
wire                             conv_Sgntin_row_00000_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00000_00002;
reg                              sign_qin_00000_00002;
wire                             conv_Sgntin_row_00000_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00000_00003;
reg                              sign_qin_00000_00003;
wire                             conv_Sgntin_row_00000_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00000_00004;
reg                              sign_qin_00000_00004;
wire                             conv_Sgntin_row_00000_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00000_00005;
reg                              sign_qin_00000_00005;
wire                             conv_Sgntin_row_00000_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00000_00006;
reg                              sign_qin_00000_00006;
wire                             conv_Sgntin_row_00000_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00000_00007;
reg                              sign_qin_00000_00007;
wire                             conv_Sgntin_row_00001_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00001_00000;
reg                              sign_qin_00001_00000;
wire                             conv_Sgntin_row_00001_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00001_00001;
reg                              sign_qin_00001_00001;
wire                             conv_Sgntin_row_00001_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00001_00002;
reg                              sign_qin_00001_00002;
wire                             conv_Sgntin_row_00001_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00001_00003;
reg                              sign_qin_00001_00003;
wire                             conv_Sgntin_row_00001_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00001_00004;
reg                              sign_qin_00001_00004;
wire                             conv_Sgntin_row_00001_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00001_00005;
reg                              sign_qin_00001_00005;
wire                             conv_Sgntin_row_00001_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00001_00006;
reg                              sign_qin_00001_00006;
wire                             conv_Sgntin_row_00001_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00001_00007;
reg                              sign_qin_00001_00007;
wire                             conv_Sgntin_row_00002_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00002_00000;
reg                              sign_qin_00002_00000;
wire                             conv_Sgntin_row_00002_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00002_00001;
reg                              sign_qin_00002_00001;
wire                             conv_Sgntin_row_00002_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00002_00002;
reg                              sign_qin_00002_00002;
wire                             conv_Sgntin_row_00002_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00002_00003;
reg                              sign_qin_00002_00003;
wire                             conv_Sgntin_row_00002_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00002_00004;
reg                              sign_qin_00002_00004;
wire                             conv_Sgntin_row_00002_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00002_00005;
reg                              sign_qin_00002_00005;
wire                             conv_Sgntin_row_00002_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00002_00006;
reg                              sign_qin_00002_00006;
wire                             conv_Sgntin_row_00002_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00002_00007;
reg                              sign_qin_00002_00007;
wire                             conv_Sgntin_row_00003_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00003_00000;
reg                              sign_qin_00003_00000;
wire                             conv_Sgntin_row_00003_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00003_00001;
reg                              sign_qin_00003_00001;
wire                             conv_Sgntin_row_00003_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00003_00002;
reg                              sign_qin_00003_00002;
wire                             conv_Sgntin_row_00003_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00003_00003;
reg                              sign_qin_00003_00003;
wire                             conv_Sgntin_row_00003_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00003_00004;
reg                              sign_qin_00003_00004;
wire                             conv_Sgntin_row_00003_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00003_00005;
reg                              sign_qin_00003_00005;
wire                             conv_Sgntin_row_00003_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00003_00006;
reg                              sign_qin_00003_00006;
wire                             conv_Sgntin_row_00003_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00003_00007;
reg                              sign_qin_00003_00007;
wire                             conv_Sgntin_row_00004_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00004_00000;
reg                              sign_qin_00004_00000;
wire                             conv_Sgntin_row_00004_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00004_00001;
reg                              sign_qin_00004_00001;
wire                             conv_Sgntin_row_00004_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00004_00002;
reg                              sign_qin_00004_00002;
wire                             conv_Sgntin_row_00004_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00004_00003;
reg                              sign_qin_00004_00003;
wire                             conv_Sgntin_row_00004_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00004_00004;
reg                              sign_qin_00004_00004;
wire                             conv_Sgntin_row_00004_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00004_00005;
reg                              sign_qin_00004_00005;
wire                             conv_Sgntin_row_00004_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00004_00006;
reg                              sign_qin_00004_00006;
wire                             conv_Sgntin_row_00004_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00004_00007;
reg                              sign_qin_00004_00007;
wire                             conv_Sgntin_row_00004_00008;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00004_00008;
reg                              sign_qin_00004_00008;
wire                             conv_Sgntin_row_00004_00009;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00004_00009;
reg                              sign_qin_00004_00009;
wire                             conv_Sgntin_row_00005_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00005_00000;
reg                              sign_qin_00005_00000;
wire                             conv_Sgntin_row_00005_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00005_00001;
reg                              sign_qin_00005_00001;
wire                             conv_Sgntin_row_00005_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00005_00002;
reg                              sign_qin_00005_00002;
wire                             conv_Sgntin_row_00005_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00005_00003;
reg                              sign_qin_00005_00003;
wire                             conv_Sgntin_row_00005_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00005_00004;
reg                              sign_qin_00005_00004;
wire                             conv_Sgntin_row_00005_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00005_00005;
reg                              sign_qin_00005_00005;
wire                             conv_Sgntin_row_00005_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00005_00006;
reg                              sign_qin_00005_00006;
wire                             conv_Sgntin_row_00005_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00005_00007;
reg                              sign_qin_00005_00007;
wire                             conv_Sgntin_row_00005_00008;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00005_00008;
reg                              sign_qin_00005_00008;
wire                             conv_Sgntin_row_00005_00009;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00005_00009;
reg                              sign_qin_00005_00009;
wire                             conv_Sgntin_row_00006_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00006_00000;
reg                              sign_qin_00006_00000;
wire                             conv_Sgntin_row_00006_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00006_00001;
reg                              sign_qin_00006_00001;
wire                             conv_Sgntin_row_00006_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00006_00002;
reg                              sign_qin_00006_00002;
wire                             conv_Sgntin_row_00006_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00006_00003;
reg                              sign_qin_00006_00003;
wire                             conv_Sgntin_row_00006_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00006_00004;
reg                              sign_qin_00006_00004;
wire                             conv_Sgntin_row_00006_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00006_00005;
reg                              sign_qin_00006_00005;
wire                             conv_Sgntin_row_00006_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00006_00006;
reg                              sign_qin_00006_00006;
wire                             conv_Sgntin_row_00006_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00006_00007;
reg                              sign_qin_00006_00007;
wire                             conv_Sgntin_row_00006_00008;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00006_00008;
reg                              sign_qin_00006_00008;
wire                             conv_Sgntin_row_00006_00009;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00006_00009;
reg                              sign_qin_00006_00009;
wire                             conv_Sgntin_row_00007_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00007_00000;
reg                              sign_qin_00007_00000;
wire                             conv_Sgntin_row_00007_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00007_00001;
reg                              sign_qin_00007_00001;
wire                             conv_Sgntin_row_00007_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00007_00002;
reg                              sign_qin_00007_00002;
wire                             conv_Sgntin_row_00007_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00007_00003;
reg                              sign_qin_00007_00003;
wire                             conv_Sgntin_row_00007_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00007_00004;
reg                              sign_qin_00007_00004;
wire                             conv_Sgntin_row_00007_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00007_00005;
reg                              sign_qin_00007_00005;
wire                             conv_Sgntin_row_00007_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00007_00006;
reg                              sign_qin_00007_00006;
wire                             conv_Sgntin_row_00007_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00007_00007;
reg                              sign_qin_00007_00007;
wire                             conv_Sgntin_row_00007_00008;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00007_00008;
reg                              sign_qin_00007_00008;
wire                             conv_Sgntin_row_00007_00009;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00007_00009;
reg                              sign_qin_00007_00009;
wire                             conv_Sgntin_row_00008_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00008_00000;
reg                              sign_qin_00008_00000;
wire                             conv_Sgntin_row_00008_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00008_00001;
reg                              sign_qin_00008_00001;
wire                             conv_Sgntin_row_00008_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00008_00002;
reg                              sign_qin_00008_00002;
wire                             conv_Sgntin_row_00008_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00008_00003;
reg                              sign_qin_00008_00003;
wire                             conv_Sgntin_row_00008_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00008_00004;
reg                              sign_qin_00008_00004;
wire                             conv_Sgntin_row_00008_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00008_00005;
reg                              sign_qin_00008_00005;
wire                             conv_Sgntin_row_00008_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00008_00006;
reg                              sign_qin_00008_00006;
wire                             conv_Sgntin_row_00008_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00008_00007;
reg                              sign_qin_00008_00007;
wire                             conv_Sgntin_row_00009_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00009_00000;
reg                              sign_qin_00009_00000;
wire                             conv_Sgntin_row_00009_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00009_00001;
reg                              sign_qin_00009_00001;
wire                             conv_Sgntin_row_00009_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00009_00002;
reg                              sign_qin_00009_00002;
wire                             conv_Sgntin_row_00009_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00009_00003;
reg                              sign_qin_00009_00003;
wire                             conv_Sgntin_row_00009_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00009_00004;
reg                              sign_qin_00009_00004;
wire                             conv_Sgntin_row_00009_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00009_00005;
reg                              sign_qin_00009_00005;
wire                             conv_Sgntin_row_00009_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00009_00006;
reg                              sign_qin_00009_00006;
wire                             conv_Sgntin_row_00009_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00009_00007;
reg                              sign_qin_00009_00007;
wire                             conv_Sgntin_row_00010_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00010_00000;
reg                              sign_qin_00010_00000;
wire                             conv_Sgntin_row_00010_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00010_00001;
reg                              sign_qin_00010_00001;
wire                             conv_Sgntin_row_00010_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00010_00002;
reg                              sign_qin_00010_00002;
wire                             conv_Sgntin_row_00010_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00010_00003;
reg                              sign_qin_00010_00003;
wire                             conv_Sgntin_row_00010_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00010_00004;
reg                              sign_qin_00010_00004;
wire                             conv_Sgntin_row_00010_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00010_00005;
reg                              sign_qin_00010_00005;
wire                             conv_Sgntin_row_00010_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00010_00006;
reg                              sign_qin_00010_00006;
wire                             conv_Sgntin_row_00010_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00010_00007;
reg                              sign_qin_00010_00007;
wire                             conv_Sgntin_row_00011_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00011_00000;
reg                              sign_qin_00011_00000;
wire                             conv_Sgntin_row_00011_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00011_00001;
reg                              sign_qin_00011_00001;
wire                             conv_Sgntin_row_00011_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00011_00002;
reg                              sign_qin_00011_00002;
wire                             conv_Sgntin_row_00011_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00011_00003;
reg                              sign_qin_00011_00003;
wire                             conv_Sgntin_row_00011_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00011_00004;
reg                              sign_qin_00011_00004;
wire                             conv_Sgntin_row_00011_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00011_00005;
reg                              sign_qin_00011_00005;
wire                             conv_Sgntin_row_00011_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00011_00006;
reg                              sign_qin_00011_00006;
wire                             conv_Sgntin_row_00011_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00011_00007;
reg                              sign_qin_00011_00007;
wire                             conv_Sgntin_row_00012_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00012_00000;
reg                              sign_qin_00012_00000;
wire                             conv_Sgntin_row_00012_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00012_00001;
reg                              sign_qin_00012_00001;
wire                             conv_Sgntin_row_00012_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00012_00002;
reg                              sign_qin_00012_00002;
wire                             conv_Sgntin_row_00012_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00012_00003;
reg                              sign_qin_00012_00003;
wire                             conv_Sgntin_row_00012_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00012_00004;
reg                              sign_qin_00012_00004;
wire                             conv_Sgntin_row_00012_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00012_00005;
reg                              sign_qin_00012_00005;
wire                             conv_Sgntin_row_00012_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00012_00006;
reg                              sign_qin_00012_00006;
wire                             conv_Sgntin_row_00012_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00012_00007;
reg                              sign_qin_00012_00007;
wire                             conv_Sgntin_row_00012_00008;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00012_00008;
reg                              sign_qin_00012_00008;
wire                             conv_Sgntin_row_00012_00009;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00012_00009;
reg                              sign_qin_00012_00009;
wire                             conv_Sgntin_row_00013_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00013_00000;
reg                              sign_qin_00013_00000;
wire                             conv_Sgntin_row_00013_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00013_00001;
reg                              sign_qin_00013_00001;
wire                             conv_Sgntin_row_00013_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00013_00002;
reg                              sign_qin_00013_00002;
wire                             conv_Sgntin_row_00013_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00013_00003;
reg                              sign_qin_00013_00003;
wire                             conv_Sgntin_row_00013_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00013_00004;
reg                              sign_qin_00013_00004;
wire                             conv_Sgntin_row_00013_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00013_00005;
reg                              sign_qin_00013_00005;
wire                             conv_Sgntin_row_00013_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00013_00006;
reg                              sign_qin_00013_00006;
wire                             conv_Sgntin_row_00013_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00013_00007;
reg                              sign_qin_00013_00007;
wire                             conv_Sgntin_row_00013_00008;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00013_00008;
reg                              sign_qin_00013_00008;
wire                             conv_Sgntin_row_00013_00009;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00013_00009;
reg                              sign_qin_00013_00009;
wire                             conv_Sgntin_row_00014_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00014_00000;
reg                              sign_qin_00014_00000;
wire                             conv_Sgntin_row_00014_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00014_00001;
reg                              sign_qin_00014_00001;
wire                             conv_Sgntin_row_00014_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00014_00002;
reg                              sign_qin_00014_00002;
wire                             conv_Sgntin_row_00014_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00014_00003;
reg                              sign_qin_00014_00003;
wire                             conv_Sgntin_row_00014_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00014_00004;
reg                              sign_qin_00014_00004;
wire                             conv_Sgntin_row_00014_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00014_00005;
reg                              sign_qin_00014_00005;
wire                             conv_Sgntin_row_00014_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00014_00006;
reg                              sign_qin_00014_00006;
wire                             conv_Sgntin_row_00014_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00014_00007;
reg                              sign_qin_00014_00007;
wire                             conv_Sgntin_row_00014_00008;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00014_00008;
reg                              sign_qin_00014_00008;
wire                             conv_Sgntin_row_00014_00009;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00014_00009;
reg                              sign_qin_00014_00009;
wire                             conv_Sgntin_row_00015_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00015_00000;
reg                              sign_qin_00015_00000;
wire                             conv_Sgntin_row_00015_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00015_00001;
reg                              sign_qin_00015_00001;
wire                             conv_Sgntin_row_00015_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00015_00002;
reg                              sign_qin_00015_00002;
wire                             conv_Sgntin_row_00015_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00015_00003;
reg                              sign_qin_00015_00003;
wire                             conv_Sgntin_row_00015_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00015_00004;
reg                              sign_qin_00015_00004;
wire                             conv_Sgntin_row_00015_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00015_00005;
reg                              sign_qin_00015_00005;
wire                             conv_Sgntin_row_00015_00006;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00015_00006;
reg                              sign_qin_00015_00006;
wire                             conv_Sgntin_row_00015_00007;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00015_00007;
reg                              sign_qin_00015_00007;
wire                             conv_Sgntin_row_00015_00008;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00015_00008;
reg                              sign_qin_00015_00008;
wire                             conv_Sgntin_row_00015_00009;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00015_00009;
reg                              sign_qin_00015_00009;
wire                             conv_Sgntin_row_00016_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00016_00000;
reg                              sign_qin_00016_00000;
wire                             conv_Sgntin_row_00016_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00016_00001;
reg                              sign_qin_00016_00001;
wire                             conv_Sgntin_row_00016_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00016_00002;
reg                              sign_qin_00016_00002;
wire                             conv_Sgntin_row_00016_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00016_00003;
reg                              sign_qin_00016_00003;
wire                             conv_Sgntin_row_00017_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00017_00000;
reg                              sign_qin_00017_00000;
wire                             conv_Sgntin_row_00017_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00017_00001;
reg                              sign_qin_00017_00001;
wire                             conv_Sgntin_row_00017_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00017_00002;
reg                              sign_qin_00017_00002;
wire                             conv_Sgntin_row_00017_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00017_00003;
reg                              sign_qin_00017_00003;
wire                             conv_Sgntin_row_00018_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00018_00000;
reg                              sign_qin_00018_00000;
wire                             conv_Sgntin_row_00018_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00018_00001;
reg                              sign_qin_00018_00001;
wire                             conv_Sgntin_row_00018_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00018_00002;
reg                              sign_qin_00018_00002;
wire                             conv_Sgntin_row_00018_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00018_00003;
reg                              sign_qin_00018_00003;
wire                             conv_Sgntin_row_00019_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00019_00000;
reg                              sign_qin_00019_00000;
wire                             conv_Sgntin_row_00019_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00019_00001;
reg                              sign_qin_00019_00001;
wire                             conv_Sgntin_row_00019_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00019_00002;
reg                              sign_qin_00019_00002;
wire                             conv_Sgntin_row_00019_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00019_00003;
reg                              sign_qin_00019_00003;
wire                             conv_Sgntin_row_00020_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00020_00000;
reg                              sign_qin_00020_00000;
wire                             conv_Sgntin_row_00020_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00020_00001;
reg                              sign_qin_00020_00001;
wire                             conv_Sgntin_row_00020_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00020_00002;
reg                              sign_qin_00020_00002;
wire                             conv_Sgntin_row_00020_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00020_00003;
reg                              sign_qin_00020_00003;
wire                             conv_Sgntin_row_00020_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00020_00004;
reg                              sign_qin_00020_00004;
wire                             conv_Sgntin_row_00020_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00020_00005;
reg                              sign_qin_00020_00005;
wire                             conv_Sgntin_row_00021_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00021_00000;
reg                              sign_qin_00021_00000;
wire                             conv_Sgntin_row_00021_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00021_00001;
reg                              sign_qin_00021_00001;
wire                             conv_Sgntin_row_00021_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00021_00002;
reg                              sign_qin_00021_00002;
wire                             conv_Sgntin_row_00021_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00021_00003;
reg                              sign_qin_00021_00003;
wire                             conv_Sgntin_row_00021_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00021_00004;
reg                              sign_qin_00021_00004;
wire                             conv_Sgntin_row_00021_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00021_00005;
reg                              sign_qin_00021_00005;
wire                             conv_Sgntin_row_00022_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00022_00000;
reg                              sign_qin_00022_00000;
wire                             conv_Sgntin_row_00022_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00022_00001;
reg                              sign_qin_00022_00001;
wire                             conv_Sgntin_row_00022_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00022_00002;
reg                              sign_qin_00022_00002;
wire                             conv_Sgntin_row_00022_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00022_00003;
reg                              sign_qin_00022_00003;
wire                             conv_Sgntin_row_00022_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00022_00004;
reg                              sign_qin_00022_00004;
wire                             conv_Sgntin_row_00022_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00022_00005;
reg                              sign_qin_00022_00005;
wire                             conv_Sgntin_row_00023_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00023_00000;
reg                              sign_qin_00023_00000;
wire                             conv_Sgntin_row_00023_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00023_00001;
reg                              sign_qin_00023_00001;
wire                             conv_Sgntin_row_00023_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00023_00002;
reg                              sign_qin_00023_00002;
wire                             conv_Sgntin_row_00023_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00023_00003;
reg                              sign_qin_00023_00003;
wire                             conv_Sgntin_row_00023_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00023_00004;
reg                              sign_qin_00023_00004;
wire                             conv_Sgntin_row_00023_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00023_00005;
reg                              sign_qin_00023_00005;
wire                             conv_Sgntin_row_00024_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00024_00000;
reg                              sign_qin_00024_00000;
wire                             conv_Sgntin_row_00024_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00024_00001;
reg                              sign_qin_00024_00001;
wire                             conv_Sgntin_row_00024_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00024_00002;
reg                              sign_qin_00024_00002;
wire                             conv_Sgntin_row_00024_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00024_00003;
reg                              sign_qin_00024_00003;
wire                             conv_Sgntin_row_00024_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00024_00004;
reg                              sign_qin_00024_00004;
wire                             conv_Sgntin_row_00024_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00024_00005;
reg                              sign_qin_00024_00005;
wire                             conv_Sgntin_row_00025_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00025_00000;
reg                              sign_qin_00025_00000;
wire                             conv_Sgntin_row_00025_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00025_00001;
reg                              sign_qin_00025_00001;
wire                             conv_Sgntin_row_00025_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00025_00002;
reg                              sign_qin_00025_00002;
wire                             conv_Sgntin_row_00025_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00025_00003;
reg                              sign_qin_00025_00003;
wire                             conv_Sgntin_row_00025_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00025_00004;
reg                              sign_qin_00025_00004;
wire                             conv_Sgntin_row_00025_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00025_00005;
reg                              sign_qin_00025_00005;
wire                             conv_Sgntin_row_00026_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00026_00000;
reg                              sign_qin_00026_00000;
wire                             conv_Sgntin_row_00026_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00026_00001;
reg                              sign_qin_00026_00001;
wire                             conv_Sgntin_row_00026_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00026_00002;
reg                              sign_qin_00026_00002;
wire                             conv_Sgntin_row_00026_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00026_00003;
reg                              sign_qin_00026_00003;
wire                             conv_Sgntin_row_00026_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00026_00004;
reg                              sign_qin_00026_00004;
wire                             conv_Sgntin_row_00026_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00026_00005;
reg                              sign_qin_00026_00005;
wire                             conv_Sgntin_row_00027_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00027_00000;
reg                              sign_qin_00027_00000;
wire                             conv_Sgntin_row_00027_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00027_00001;
reg                              sign_qin_00027_00001;
wire                             conv_Sgntin_row_00027_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00027_00002;
reg                              sign_qin_00027_00002;
wire                             conv_Sgntin_row_00027_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00027_00003;
reg                              sign_qin_00027_00003;
wire                             conv_Sgntin_row_00027_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00027_00004;
reg                              sign_qin_00027_00004;
wire                             conv_Sgntin_row_00027_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00027_00005;
reg                              sign_qin_00027_00005;
wire                             conv_Sgntin_row_00028_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00028_00000;
reg                              sign_qin_00028_00000;
wire                             conv_Sgntin_row_00028_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00028_00001;
reg                              sign_qin_00028_00001;
wire                             conv_Sgntin_row_00028_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00028_00002;
reg                              sign_qin_00028_00002;
wire                             conv_Sgntin_row_00028_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00028_00003;
reg                              sign_qin_00028_00003;
wire                             conv_Sgntin_row_00028_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00028_00004;
reg                              sign_qin_00028_00004;
wire                             conv_Sgntin_row_00028_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00028_00005;
reg                              sign_qin_00028_00005;
wire                             conv_Sgntin_row_00029_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00029_00000;
reg                              sign_qin_00029_00000;
wire                             conv_Sgntin_row_00029_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00029_00001;
reg                              sign_qin_00029_00001;
wire                             conv_Sgntin_row_00029_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00029_00002;
reg                              sign_qin_00029_00002;
wire                             conv_Sgntin_row_00029_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00029_00003;
reg                              sign_qin_00029_00003;
wire                             conv_Sgntin_row_00029_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00029_00004;
reg                              sign_qin_00029_00004;
wire                             conv_Sgntin_row_00029_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00029_00005;
reg                              sign_qin_00029_00005;
wire                             conv_Sgntin_row_00030_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00030_00000;
reg                              sign_qin_00030_00000;
wire                             conv_Sgntin_row_00030_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00030_00001;
reg                              sign_qin_00030_00001;
wire                             conv_Sgntin_row_00030_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00030_00002;
reg                              sign_qin_00030_00002;
wire                             conv_Sgntin_row_00030_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00030_00003;
reg                              sign_qin_00030_00003;
wire                             conv_Sgntin_row_00030_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00030_00004;
reg                              sign_qin_00030_00004;
wire                             conv_Sgntin_row_00030_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00030_00005;
reg                              sign_qin_00030_00005;
wire                             conv_Sgntin_row_00031_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00031_00000;
reg                              sign_qin_00031_00000;
wire                             conv_Sgntin_row_00031_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00031_00001;
reg                              sign_qin_00031_00001;
wire                             conv_Sgntin_row_00031_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00031_00002;
reg                              sign_qin_00031_00002;
wire                             conv_Sgntin_row_00031_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00031_00003;
reg                              sign_qin_00031_00003;
wire                             conv_Sgntin_row_00031_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00031_00004;
reg                              sign_qin_00031_00004;
wire                             conv_Sgntin_row_00031_00005;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00031_00005;
reg                              sign_qin_00031_00005;
wire                             conv_Sgntin_row_00032_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00032_00000;
reg                              sign_qin_00032_00000;
wire                             conv_Sgntin_row_00032_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00032_00001;
reg                              sign_qin_00032_00001;
wire                             conv_Sgntin_row_00032_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00032_00002;
reg                              sign_qin_00032_00002;
wire                             conv_Sgntin_row_00032_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00032_00003;
reg                              sign_qin_00032_00003;
wire                             conv_Sgntin_row_00033_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00033_00000;
reg                              sign_qin_00033_00000;
wire                             conv_Sgntin_row_00033_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00033_00001;
reg                              sign_qin_00033_00001;
wire                             conv_Sgntin_row_00033_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00033_00002;
reg                              sign_qin_00033_00002;
wire                             conv_Sgntin_row_00033_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00033_00003;
reg                              sign_qin_00033_00003;
wire                             conv_Sgntin_row_00034_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00034_00000;
reg                              sign_qin_00034_00000;
wire                             conv_Sgntin_row_00034_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00034_00001;
reg                              sign_qin_00034_00001;
wire                             conv_Sgntin_row_00034_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00034_00002;
reg                              sign_qin_00034_00002;
wire                             conv_Sgntin_row_00034_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00034_00003;
reg                              sign_qin_00034_00003;
wire                             conv_Sgntin_row_00035_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00035_00000;
reg                              sign_qin_00035_00000;
wire                             conv_Sgntin_row_00035_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00035_00001;
reg                              sign_qin_00035_00001;
wire                             conv_Sgntin_row_00035_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00035_00002;
reg                              sign_qin_00035_00002;
wire                             conv_Sgntin_row_00035_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00035_00003;
reg                              sign_qin_00035_00003;
wire                             conv_Sgntin_row_00036_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00036_00000;
reg                              sign_qin_00036_00000;
wire                             conv_Sgntin_row_00036_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00036_00001;
reg                              sign_qin_00036_00001;
wire                             conv_Sgntin_row_00036_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00036_00002;
reg                              sign_qin_00036_00002;
wire                             conv_Sgntin_row_00036_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00036_00003;
reg                              sign_qin_00036_00003;
wire                             conv_Sgntin_row_00036_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00036_00004;
reg                              sign_qin_00036_00004;
wire                             conv_Sgntin_row_00037_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00037_00000;
reg                              sign_qin_00037_00000;
wire                             conv_Sgntin_row_00037_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00037_00001;
reg                              sign_qin_00037_00001;
wire                             conv_Sgntin_row_00037_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00037_00002;
reg                              sign_qin_00037_00002;
wire                             conv_Sgntin_row_00037_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00037_00003;
reg                              sign_qin_00037_00003;
wire                             conv_Sgntin_row_00037_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00037_00004;
reg                              sign_qin_00037_00004;
wire                             conv_Sgntin_row_00038_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00038_00000;
reg                              sign_qin_00038_00000;
wire                             conv_Sgntin_row_00038_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00038_00001;
reg                              sign_qin_00038_00001;
wire                             conv_Sgntin_row_00038_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00038_00002;
reg                              sign_qin_00038_00002;
wire                             conv_Sgntin_row_00038_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00038_00003;
reg                              sign_qin_00038_00003;
wire                             conv_Sgntin_row_00038_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00038_00004;
reg                              sign_qin_00038_00004;
wire                             conv_Sgntin_row_00039_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00039_00000;
reg                              sign_qin_00039_00000;
wire                             conv_Sgntin_row_00039_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00039_00001;
reg                              sign_qin_00039_00001;
wire                             conv_Sgntin_row_00039_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00039_00002;
reg                              sign_qin_00039_00002;
wire                             conv_Sgntin_row_00039_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00039_00003;
reg                              sign_qin_00039_00003;
wire                             conv_Sgntin_row_00039_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00039_00004;
reg                              sign_qin_00039_00004;
wire                             conv_Sgntin_row_00040_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00040_00000;
reg                              sign_qin_00040_00000;
wire                             conv_Sgntin_row_00040_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00040_00001;
reg                              sign_qin_00040_00001;
wire                             conv_Sgntin_row_00040_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00040_00002;
reg                              sign_qin_00040_00002;
wire                             conv_Sgntin_row_00040_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00040_00003;
reg                              sign_qin_00040_00003;
wire                             conv_Sgntin_row_00040_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00040_00004;
reg                              sign_qin_00040_00004;
wire                             conv_Sgntin_row_00041_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00041_00000;
reg                              sign_qin_00041_00000;
wire                             conv_Sgntin_row_00041_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00041_00001;
reg                              sign_qin_00041_00001;
wire                             conv_Sgntin_row_00041_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00041_00002;
reg                              sign_qin_00041_00002;
wire                             conv_Sgntin_row_00041_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00041_00003;
reg                              sign_qin_00041_00003;
wire                             conv_Sgntin_row_00041_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00041_00004;
reg                              sign_qin_00041_00004;
wire                             conv_Sgntin_row_00042_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00042_00000;
reg                              sign_qin_00042_00000;
wire                             conv_Sgntin_row_00042_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00042_00001;
reg                              sign_qin_00042_00001;
wire                             conv_Sgntin_row_00042_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00042_00002;
reg                              sign_qin_00042_00002;
wire                             conv_Sgntin_row_00042_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00042_00003;
reg                              sign_qin_00042_00003;
wire                             conv_Sgntin_row_00042_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00042_00004;
reg                              sign_qin_00042_00004;
wire                             conv_Sgntin_row_00043_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00043_00000;
reg                              sign_qin_00043_00000;
wire                             conv_Sgntin_row_00043_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00043_00001;
reg                              sign_qin_00043_00001;
wire                             conv_Sgntin_row_00043_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00043_00002;
reg                              sign_qin_00043_00002;
wire                             conv_Sgntin_row_00043_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00043_00003;
reg                              sign_qin_00043_00003;
wire                             conv_Sgntin_row_00043_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00043_00004;
reg                              sign_qin_00043_00004;
wire                             conv_Sgntin_row_00044_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00044_00000;
reg                              sign_qin_00044_00000;
wire                             conv_Sgntin_row_00044_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00044_00001;
reg                              sign_qin_00044_00001;
wire                             conv_Sgntin_row_00044_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00044_00002;
reg                              sign_qin_00044_00002;
wire                             conv_Sgntin_row_00044_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00044_00003;
reg                              sign_qin_00044_00003;
wire                             conv_Sgntin_row_00044_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00044_00004;
reg                              sign_qin_00044_00004;
wire                             conv_Sgntin_row_00045_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00045_00000;
reg                              sign_qin_00045_00000;
wire                             conv_Sgntin_row_00045_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00045_00001;
reg                              sign_qin_00045_00001;
wire                             conv_Sgntin_row_00045_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00045_00002;
reg                              sign_qin_00045_00002;
wire                             conv_Sgntin_row_00045_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00045_00003;
reg                              sign_qin_00045_00003;
wire                             conv_Sgntin_row_00045_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00045_00004;
reg                              sign_qin_00045_00004;
wire                             conv_Sgntin_row_00046_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00046_00000;
reg                              sign_qin_00046_00000;
wire                             conv_Sgntin_row_00046_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00046_00001;
reg                              sign_qin_00046_00001;
wire                             conv_Sgntin_row_00046_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00046_00002;
reg                              sign_qin_00046_00002;
wire                             conv_Sgntin_row_00046_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00046_00003;
reg                              sign_qin_00046_00003;
wire                             conv_Sgntin_row_00046_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00046_00004;
reg                              sign_qin_00046_00004;
wire                             conv_Sgntin_row_00047_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00047_00000;
reg                              sign_qin_00047_00000;
wire                             conv_Sgntin_row_00047_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00047_00001;
reg                              sign_qin_00047_00001;
wire                             conv_Sgntin_row_00047_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00047_00002;
reg                              sign_qin_00047_00002;
wire                             conv_Sgntin_row_00047_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00047_00003;
reg                              sign_qin_00047_00003;
wire                             conv_Sgntin_row_00047_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00047_00004;
reg                              sign_qin_00047_00004;
wire                             conv_Sgntin_row_00048_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00048_00000;
reg                              sign_qin_00048_00000;
wire                             conv_Sgntin_row_00048_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00048_00001;
reg                              sign_qin_00048_00001;
wire                             conv_Sgntin_row_00048_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00048_00002;
reg                              sign_qin_00048_00002;
wire                             conv_Sgntin_row_00048_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00048_00003;
reg                              sign_qin_00048_00003;
wire                             conv_Sgntin_row_00049_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00049_00000;
reg                              sign_qin_00049_00000;
wire                             conv_Sgntin_row_00049_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00049_00001;
reg                              sign_qin_00049_00001;
wire                             conv_Sgntin_row_00049_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00049_00002;
reg                              sign_qin_00049_00002;
wire                             conv_Sgntin_row_00049_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00049_00003;
reg                              sign_qin_00049_00003;
wire                             conv_Sgntin_row_00050_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00050_00000;
reg                              sign_qin_00050_00000;
wire                             conv_Sgntin_row_00050_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00050_00001;
reg                              sign_qin_00050_00001;
wire                             conv_Sgntin_row_00050_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00050_00002;
reg                              sign_qin_00050_00002;
wire                             conv_Sgntin_row_00050_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00050_00003;
reg                              sign_qin_00050_00003;
wire                             conv_Sgntin_row_00051_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00051_00000;
reg                              sign_qin_00051_00000;
wire                             conv_Sgntin_row_00051_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00051_00001;
reg                              sign_qin_00051_00001;
wire                             conv_Sgntin_row_00051_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00051_00002;
reg                              sign_qin_00051_00002;
wire                             conv_Sgntin_row_00051_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00051_00003;
reg                              sign_qin_00051_00003;
wire                             conv_Sgntin_row_00052_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00052_00000;
reg                              sign_qin_00052_00000;
wire                             conv_Sgntin_row_00052_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00052_00001;
reg                              sign_qin_00052_00001;
wire                             conv_Sgntin_row_00052_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00052_00002;
reg                              sign_qin_00052_00002;
wire                             conv_Sgntin_row_00052_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00052_00003;
reg                              sign_qin_00052_00003;
wire                             conv_Sgntin_row_00052_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00052_00004;
reg                              sign_qin_00052_00004;
wire                             conv_Sgntin_row_00053_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00053_00000;
reg                              sign_qin_00053_00000;
wire                             conv_Sgntin_row_00053_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00053_00001;
reg                              sign_qin_00053_00001;
wire                             conv_Sgntin_row_00053_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00053_00002;
reg                              sign_qin_00053_00002;
wire                             conv_Sgntin_row_00053_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00053_00003;
reg                              sign_qin_00053_00003;
wire                             conv_Sgntin_row_00053_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00053_00004;
reg                              sign_qin_00053_00004;
wire                             conv_Sgntin_row_00054_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00054_00000;
reg                              sign_qin_00054_00000;
wire                             conv_Sgntin_row_00054_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00054_00001;
reg                              sign_qin_00054_00001;
wire                             conv_Sgntin_row_00054_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00054_00002;
reg                              sign_qin_00054_00002;
wire                             conv_Sgntin_row_00054_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00054_00003;
reg                              sign_qin_00054_00003;
wire                             conv_Sgntin_row_00054_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00054_00004;
reg                              sign_qin_00054_00004;
wire                             conv_Sgntin_row_00055_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00055_00000;
reg                              sign_qin_00055_00000;
wire                             conv_Sgntin_row_00055_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00055_00001;
reg                              sign_qin_00055_00001;
wire                             conv_Sgntin_row_00055_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00055_00002;
reg                              sign_qin_00055_00002;
wire                             conv_Sgntin_row_00055_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00055_00003;
reg                              sign_qin_00055_00003;
wire                             conv_Sgntin_row_00055_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00055_00004;
reg                              sign_qin_00055_00004;
wire                             conv_Sgntin_row_00056_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00056_00000;
reg                              sign_qin_00056_00000;
wire                             conv_Sgntin_row_00056_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00056_00001;
reg                              sign_qin_00056_00001;
wire                             conv_Sgntin_row_00056_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00056_00002;
reg                              sign_qin_00056_00002;
wire                             conv_Sgntin_row_00056_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00056_00003;
reg                              sign_qin_00056_00003;
wire                             conv_Sgntin_row_00056_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00056_00004;
reg                              sign_qin_00056_00004;
wire                             conv_Sgntin_row_00057_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00057_00000;
reg                              sign_qin_00057_00000;
wire                             conv_Sgntin_row_00057_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00057_00001;
reg                              sign_qin_00057_00001;
wire                             conv_Sgntin_row_00057_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00057_00002;
reg                              sign_qin_00057_00002;
wire                             conv_Sgntin_row_00057_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00057_00003;
reg                              sign_qin_00057_00003;
wire                             conv_Sgntin_row_00057_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00057_00004;
reg                              sign_qin_00057_00004;
wire                             conv_Sgntin_row_00058_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00058_00000;
reg                              sign_qin_00058_00000;
wire                             conv_Sgntin_row_00058_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00058_00001;
reg                              sign_qin_00058_00001;
wire                             conv_Sgntin_row_00058_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00058_00002;
reg                              sign_qin_00058_00002;
wire                             conv_Sgntin_row_00058_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00058_00003;
reg                              sign_qin_00058_00003;
wire                             conv_Sgntin_row_00058_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00058_00004;
reg                              sign_qin_00058_00004;
wire                             conv_Sgntin_row_00059_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00059_00000;
reg                              sign_qin_00059_00000;
wire                             conv_Sgntin_row_00059_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00059_00001;
reg                              sign_qin_00059_00001;
wire                             conv_Sgntin_row_00059_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00059_00002;
reg                              sign_qin_00059_00002;
wire                             conv_Sgntin_row_00059_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00059_00003;
reg                              sign_qin_00059_00003;
wire                             conv_Sgntin_row_00059_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00059_00004;
reg                              sign_qin_00059_00004;
wire                             conv_Sgntin_row_00060_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00060_00000;
reg                              sign_qin_00060_00000;
wire                             conv_Sgntin_row_00060_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00060_00001;
reg                              sign_qin_00060_00001;
wire                             conv_Sgntin_row_00060_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00060_00002;
reg                              sign_qin_00060_00002;
wire                             conv_Sgntin_row_00060_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00060_00003;
reg                              sign_qin_00060_00003;
wire                             conv_Sgntin_row_00061_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00061_00000;
reg                              sign_qin_00061_00000;
wire                             conv_Sgntin_row_00061_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00061_00001;
reg                              sign_qin_00061_00001;
wire                             conv_Sgntin_row_00061_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00061_00002;
reg                              sign_qin_00061_00002;
wire                             conv_Sgntin_row_00061_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00061_00003;
reg                              sign_qin_00061_00003;
wire                             conv_Sgntin_row_00062_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00062_00000;
reg                              sign_qin_00062_00000;
wire                             conv_Sgntin_row_00062_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00062_00001;
reg                              sign_qin_00062_00001;
wire                             conv_Sgntin_row_00062_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00062_00002;
reg                              sign_qin_00062_00002;
wire                             conv_Sgntin_row_00062_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00062_00003;
reg                              sign_qin_00062_00003;
wire                             conv_Sgntin_row_00063_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00063_00000;
reg                              sign_qin_00063_00000;
wire                             conv_Sgntin_row_00063_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00063_00001;
reg                              sign_qin_00063_00001;
wire                             conv_Sgntin_row_00063_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00063_00002;
reg                              sign_qin_00063_00002;
wire                             conv_Sgntin_row_00063_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00063_00003;
reg                              sign_qin_00063_00003;
wire                             conv_Sgntin_row_00064_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00064_00000;
reg                              sign_qin_00064_00000;
wire                             conv_Sgntin_row_00064_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00064_00001;
reg                              sign_qin_00064_00001;
wire                             conv_Sgntin_row_00064_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00064_00002;
reg                              sign_qin_00064_00002;
wire                             conv_Sgntin_row_00064_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00064_00003;
reg                              sign_qin_00064_00003;
wire                             conv_Sgntin_row_00064_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00064_00004;
reg                              sign_qin_00064_00004;
wire                             conv_Sgntin_row_00065_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00065_00000;
reg                              sign_qin_00065_00000;
wire                             conv_Sgntin_row_00065_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00065_00001;
reg                              sign_qin_00065_00001;
wire                             conv_Sgntin_row_00065_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00065_00002;
reg                              sign_qin_00065_00002;
wire                             conv_Sgntin_row_00065_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00065_00003;
reg                              sign_qin_00065_00003;
wire                             conv_Sgntin_row_00065_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00065_00004;
reg                              sign_qin_00065_00004;
wire                             conv_Sgntin_row_00066_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00066_00000;
reg                              sign_qin_00066_00000;
wire                             conv_Sgntin_row_00066_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00066_00001;
reg                              sign_qin_00066_00001;
wire                             conv_Sgntin_row_00066_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00066_00002;
reg                              sign_qin_00066_00002;
wire                             conv_Sgntin_row_00066_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00066_00003;
reg                              sign_qin_00066_00003;
wire                             conv_Sgntin_row_00066_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00066_00004;
reg                              sign_qin_00066_00004;
wire                             conv_Sgntin_row_00067_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00067_00000;
reg                              sign_qin_00067_00000;
wire                             conv_Sgntin_row_00067_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00067_00001;
reg                              sign_qin_00067_00001;
wire                             conv_Sgntin_row_00067_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00067_00002;
reg                              sign_qin_00067_00002;
wire                             conv_Sgntin_row_00067_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00067_00003;
reg                              sign_qin_00067_00003;
wire                             conv_Sgntin_row_00067_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00067_00004;
reg                              sign_qin_00067_00004;
wire                             conv_Sgntin_row_00068_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00068_00000;
reg                              sign_qin_00068_00000;
wire                             conv_Sgntin_row_00068_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00068_00001;
reg                              sign_qin_00068_00001;
wire                             conv_Sgntin_row_00068_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00068_00002;
reg                              sign_qin_00068_00002;
wire                             conv_Sgntin_row_00068_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00068_00003;
reg                              sign_qin_00068_00003;
wire                             conv_Sgntin_row_00068_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00068_00004;
reg                              sign_qin_00068_00004;
wire                             conv_Sgntin_row_00069_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00069_00000;
reg                              sign_qin_00069_00000;
wire                             conv_Sgntin_row_00069_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00069_00001;
reg                              sign_qin_00069_00001;
wire                             conv_Sgntin_row_00069_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00069_00002;
reg                              sign_qin_00069_00002;
wire                             conv_Sgntin_row_00069_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00069_00003;
reg                              sign_qin_00069_00003;
wire                             conv_Sgntin_row_00069_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00069_00004;
reg                              sign_qin_00069_00004;
wire                             conv_Sgntin_row_00070_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00070_00000;
reg                              sign_qin_00070_00000;
wire                             conv_Sgntin_row_00070_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00070_00001;
reg                              sign_qin_00070_00001;
wire                             conv_Sgntin_row_00070_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00070_00002;
reg                              sign_qin_00070_00002;
wire                             conv_Sgntin_row_00070_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00070_00003;
reg                              sign_qin_00070_00003;
wire                             conv_Sgntin_row_00070_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00070_00004;
reg                              sign_qin_00070_00004;
wire                             conv_Sgntin_row_00071_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00071_00000;
reg                              sign_qin_00071_00000;
wire                             conv_Sgntin_row_00071_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00071_00001;
reg                              sign_qin_00071_00001;
wire                             conv_Sgntin_row_00071_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00071_00002;
reg                              sign_qin_00071_00002;
wire                             conv_Sgntin_row_00071_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00071_00003;
reg                              sign_qin_00071_00003;
wire                             conv_Sgntin_row_00071_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00071_00004;
reg                              sign_qin_00071_00004;
wire                             conv_Sgntin_row_00072_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00072_00000;
reg                              sign_qin_00072_00000;
wire                             conv_Sgntin_row_00072_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00072_00001;
reg                              sign_qin_00072_00001;
wire                             conv_Sgntin_row_00072_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00072_00002;
reg                              sign_qin_00072_00002;
wire                             conv_Sgntin_row_00072_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00072_00003;
reg                              sign_qin_00072_00003;
wire                             conv_Sgntin_row_00073_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00073_00000;
reg                              sign_qin_00073_00000;
wire                             conv_Sgntin_row_00073_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00073_00001;
reg                              sign_qin_00073_00001;
wire                             conv_Sgntin_row_00073_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00073_00002;
reg                              sign_qin_00073_00002;
wire                             conv_Sgntin_row_00073_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00073_00003;
reg                              sign_qin_00073_00003;
wire                             conv_Sgntin_row_00074_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00074_00000;
reg                              sign_qin_00074_00000;
wire                             conv_Sgntin_row_00074_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00074_00001;
reg                              sign_qin_00074_00001;
wire                             conv_Sgntin_row_00074_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00074_00002;
reg                              sign_qin_00074_00002;
wire                             conv_Sgntin_row_00074_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00074_00003;
reg                              sign_qin_00074_00003;
wire                             conv_Sgntin_row_00075_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00075_00000;
reg                              sign_qin_00075_00000;
wire                             conv_Sgntin_row_00075_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00075_00001;
reg                              sign_qin_00075_00001;
wire                             conv_Sgntin_row_00075_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00075_00002;
reg                              sign_qin_00075_00002;
wire                             conv_Sgntin_row_00075_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00075_00003;
reg                              sign_qin_00075_00003;
wire                             conv_Sgntin_row_00076_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00076_00000;
reg                              sign_qin_00076_00000;
wire                             conv_Sgntin_row_00076_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00076_00001;
reg                              sign_qin_00076_00001;
wire                             conv_Sgntin_row_00076_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00076_00002;
reg                              sign_qin_00076_00002;
wire                             conv_Sgntin_row_00076_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00076_00003;
reg                              sign_qin_00076_00003;
wire                             conv_Sgntin_row_00077_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00077_00000;
reg                              sign_qin_00077_00000;
wire                             conv_Sgntin_row_00077_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00077_00001;
reg                              sign_qin_00077_00001;
wire                             conv_Sgntin_row_00077_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00077_00002;
reg                              sign_qin_00077_00002;
wire                             conv_Sgntin_row_00077_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00077_00003;
reg                              sign_qin_00077_00003;
wire                             conv_Sgntin_row_00078_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00078_00000;
reg                              sign_qin_00078_00000;
wire                             conv_Sgntin_row_00078_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00078_00001;
reg                              sign_qin_00078_00001;
wire                             conv_Sgntin_row_00078_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00078_00002;
reg                              sign_qin_00078_00002;
wire                             conv_Sgntin_row_00078_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00078_00003;
reg                              sign_qin_00078_00003;
wire                             conv_Sgntin_row_00079_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00079_00000;
reg                              sign_qin_00079_00000;
wire                             conv_Sgntin_row_00079_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00079_00001;
reg                              sign_qin_00079_00001;
wire                             conv_Sgntin_row_00079_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00079_00002;
reg                              sign_qin_00079_00002;
wire                             conv_Sgntin_row_00079_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00079_00003;
reg                              sign_qin_00079_00003;
wire                             conv_Sgntin_row_00080_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00080_00000;
reg                              sign_qin_00080_00000;
wire                             conv_Sgntin_row_00080_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00080_00001;
reg                              sign_qin_00080_00001;
wire                             conv_Sgntin_row_00080_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00080_00002;
reg                              sign_qin_00080_00002;
wire                             conv_Sgntin_row_00080_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00080_00003;
reg                              sign_qin_00080_00003;
wire                             conv_Sgntin_row_00081_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00081_00000;
reg                              sign_qin_00081_00000;
wire                             conv_Sgntin_row_00081_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00081_00001;
reg                              sign_qin_00081_00001;
wire                             conv_Sgntin_row_00081_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00081_00002;
reg                              sign_qin_00081_00002;
wire                             conv_Sgntin_row_00081_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00081_00003;
reg                              sign_qin_00081_00003;
wire                             conv_Sgntin_row_00082_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00082_00000;
reg                              sign_qin_00082_00000;
wire                             conv_Sgntin_row_00082_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00082_00001;
reg                              sign_qin_00082_00001;
wire                             conv_Sgntin_row_00082_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00082_00002;
reg                              sign_qin_00082_00002;
wire                             conv_Sgntin_row_00082_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00082_00003;
reg                              sign_qin_00082_00003;
wire                             conv_Sgntin_row_00083_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00083_00000;
reg                              sign_qin_00083_00000;
wire                             conv_Sgntin_row_00083_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00083_00001;
reg                              sign_qin_00083_00001;
wire                             conv_Sgntin_row_00083_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00083_00002;
reg                              sign_qin_00083_00002;
wire                             conv_Sgntin_row_00083_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00083_00003;
reg                              sign_qin_00083_00003;
wire                             conv_Sgntin_row_00084_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00084_00000;
reg                              sign_qin_00084_00000;
wire                             conv_Sgntin_row_00084_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00084_00001;
reg                              sign_qin_00084_00001;
wire                             conv_Sgntin_row_00084_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00084_00002;
reg                              sign_qin_00084_00002;
wire                             conv_Sgntin_row_00084_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00084_00003;
reg                              sign_qin_00084_00003;
wire                             conv_Sgntin_row_00085_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00085_00000;
reg                              sign_qin_00085_00000;
wire                             conv_Sgntin_row_00085_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00085_00001;
reg                              sign_qin_00085_00001;
wire                             conv_Sgntin_row_00085_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00085_00002;
reg                              sign_qin_00085_00002;
wire                             conv_Sgntin_row_00085_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00085_00003;
reg                              sign_qin_00085_00003;
wire                             conv_Sgntin_row_00086_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00086_00000;
reg                              sign_qin_00086_00000;
wire                             conv_Sgntin_row_00086_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00086_00001;
reg                              sign_qin_00086_00001;
wire                             conv_Sgntin_row_00086_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00086_00002;
reg                              sign_qin_00086_00002;
wire                             conv_Sgntin_row_00086_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00086_00003;
reg                              sign_qin_00086_00003;
wire                             conv_Sgntin_row_00087_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00087_00000;
reg                              sign_qin_00087_00000;
wire                             conv_Sgntin_row_00087_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00087_00001;
reg                              sign_qin_00087_00001;
wire                             conv_Sgntin_row_00087_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00087_00002;
reg                              sign_qin_00087_00002;
wire                             conv_Sgntin_row_00087_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00087_00003;
reg                              sign_qin_00087_00003;
wire                             conv_Sgntin_row_00088_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00088_00000;
reg                              sign_qin_00088_00000;
wire                             conv_Sgntin_row_00088_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00088_00001;
reg                              sign_qin_00088_00001;
wire                             conv_Sgntin_row_00088_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00088_00002;
reg                              sign_qin_00088_00002;
wire                             conv_Sgntin_row_00089_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00089_00000;
reg                              sign_qin_00089_00000;
wire                             conv_Sgntin_row_00089_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00089_00001;
reg                              sign_qin_00089_00001;
wire                             conv_Sgntin_row_00089_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00089_00002;
reg                              sign_qin_00089_00002;
wire                             conv_Sgntin_row_00090_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00090_00000;
reg                              sign_qin_00090_00000;
wire                             conv_Sgntin_row_00090_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00090_00001;
reg                              sign_qin_00090_00001;
wire                             conv_Sgntin_row_00090_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00090_00002;
reg                              sign_qin_00090_00002;
wire                             conv_Sgntin_row_00091_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00091_00000;
reg                              sign_qin_00091_00000;
wire                             conv_Sgntin_row_00091_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00091_00001;
reg                              sign_qin_00091_00001;
wire                             conv_Sgntin_row_00091_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00091_00002;
reg                              sign_qin_00091_00002;
wire                             conv_Sgntin_row_00092_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00092_00000;
reg                              sign_qin_00092_00000;
wire                             conv_Sgntin_row_00092_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00092_00001;
reg                              sign_qin_00092_00001;
wire                             conv_Sgntin_row_00092_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00092_00002;
reg                              sign_qin_00092_00002;
wire                             conv_Sgntin_row_00092_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00092_00003;
reg                              sign_qin_00092_00003;
wire                             conv_Sgntin_row_00093_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00093_00000;
reg                              sign_qin_00093_00000;
wire                             conv_Sgntin_row_00093_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00093_00001;
reg                              sign_qin_00093_00001;
wire                             conv_Sgntin_row_00093_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00093_00002;
reg                              sign_qin_00093_00002;
wire                             conv_Sgntin_row_00093_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00093_00003;
reg                              sign_qin_00093_00003;
wire                             conv_Sgntin_row_00094_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00094_00000;
reg                              sign_qin_00094_00000;
wire                             conv_Sgntin_row_00094_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00094_00001;
reg                              sign_qin_00094_00001;
wire                             conv_Sgntin_row_00094_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00094_00002;
reg                              sign_qin_00094_00002;
wire                             conv_Sgntin_row_00094_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00094_00003;
reg                              sign_qin_00094_00003;
wire                             conv_Sgntin_row_00095_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00095_00000;
reg                              sign_qin_00095_00000;
wire                             conv_Sgntin_row_00095_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00095_00001;
reg                              sign_qin_00095_00001;
wire                             conv_Sgntin_row_00095_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00095_00002;
reg                              sign_qin_00095_00002;
wire                             conv_Sgntin_row_00095_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00095_00003;
reg                              sign_qin_00095_00003;
wire                             conv_Sgntin_row_00096_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00096_00000;
reg                              sign_qin_00096_00000;
wire                             conv_Sgntin_row_00096_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00096_00001;
reg                              sign_qin_00096_00001;
wire                             conv_Sgntin_row_00096_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00096_00002;
reg                              sign_qin_00096_00002;
wire                             conv_Sgntin_row_00096_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00096_00003;
reg                              sign_qin_00096_00003;
wire                             conv_Sgntin_row_00097_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00097_00000;
reg                              sign_qin_00097_00000;
wire                             conv_Sgntin_row_00097_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00097_00001;
reg                              sign_qin_00097_00001;
wire                             conv_Sgntin_row_00097_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00097_00002;
reg                              sign_qin_00097_00002;
wire                             conv_Sgntin_row_00097_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00097_00003;
reg                              sign_qin_00097_00003;
wire                             conv_Sgntin_row_00098_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00098_00000;
reg                              sign_qin_00098_00000;
wire                             conv_Sgntin_row_00098_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00098_00001;
reg                              sign_qin_00098_00001;
wire                             conv_Sgntin_row_00098_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00098_00002;
reg                              sign_qin_00098_00002;
wire                             conv_Sgntin_row_00098_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00098_00003;
reg                              sign_qin_00098_00003;
wire                             conv_Sgntin_row_00099_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00099_00000;
reg                              sign_qin_00099_00000;
wire                             conv_Sgntin_row_00099_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00099_00001;
reg                              sign_qin_00099_00001;
wire                             conv_Sgntin_row_00099_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00099_00002;
reg                              sign_qin_00099_00002;
wire                             conv_Sgntin_row_00099_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00099_00003;
reg                              sign_qin_00099_00003;
wire                             conv_Sgntin_row_00100_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00100_00000;
reg                              sign_qin_00100_00000;
wire                             conv_Sgntin_row_00100_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00100_00001;
reg                              sign_qin_00100_00001;
wire                             conv_Sgntin_row_00100_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00100_00002;
reg                              sign_qin_00100_00002;
wire                             conv_Sgntin_row_00101_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00101_00000;
reg                              sign_qin_00101_00000;
wire                             conv_Sgntin_row_00101_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00101_00001;
reg                              sign_qin_00101_00001;
wire                             conv_Sgntin_row_00101_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00101_00002;
reg                              sign_qin_00101_00002;
wire                             conv_Sgntin_row_00102_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00102_00000;
reg                              sign_qin_00102_00000;
wire                             conv_Sgntin_row_00102_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00102_00001;
reg                              sign_qin_00102_00001;
wire                             conv_Sgntin_row_00102_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00102_00002;
reg                              sign_qin_00102_00002;
wire                             conv_Sgntin_row_00103_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00103_00000;
reg                              sign_qin_00103_00000;
wire                             conv_Sgntin_row_00103_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00103_00001;
reg                              sign_qin_00103_00001;
wire                             conv_Sgntin_row_00103_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00103_00002;
reg                              sign_qin_00103_00002;
wire                             conv_Sgntin_row_00104_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00104_00000;
reg                              sign_qin_00104_00000;
wire                             conv_Sgntin_row_00104_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00104_00001;
reg                              sign_qin_00104_00001;
wire                             conv_Sgntin_row_00104_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00104_00002;
reg                              sign_qin_00104_00002;
wire                             conv_Sgntin_row_00104_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00104_00003;
reg                              sign_qin_00104_00003;
wire                             conv_Sgntin_row_00104_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00104_00004;
reg                              sign_qin_00104_00004;
wire                             conv_Sgntin_row_00105_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00105_00000;
reg                              sign_qin_00105_00000;
wire                             conv_Sgntin_row_00105_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00105_00001;
reg                              sign_qin_00105_00001;
wire                             conv_Sgntin_row_00105_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00105_00002;
reg                              sign_qin_00105_00002;
wire                             conv_Sgntin_row_00105_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00105_00003;
reg                              sign_qin_00105_00003;
wire                             conv_Sgntin_row_00105_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00105_00004;
reg                              sign_qin_00105_00004;
wire                             conv_Sgntin_row_00106_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00106_00000;
reg                              sign_qin_00106_00000;
wire                             conv_Sgntin_row_00106_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00106_00001;
reg                              sign_qin_00106_00001;
wire                             conv_Sgntin_row_00106_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00106_00002;
reg                              sign_qin_00106_00002;
wire                             conv_Sgntin_row_00106_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00106_00003;
reg                              sign_qin_00106_00003;
wire                             conv_Sgntin_row_00106_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00106_00004;
reg                              sign_qin_00106_00004;
wire                             conv_Sgntin_row_00107_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00107_00000;
reg                              sign_qin_00107_00000;
wire                             conv_Sgntin_row_00107_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00107_00001;
reg                              sign_qin_00107_00001;
wire                             conv_Sgntin_row_00107_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00107_00002;
reg                              sign_qin_00107_00002;
wire                             conv_Sgntin_row_00107_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00107_00003;
reg                              sign_qin_00107_00003;
wire                             conv_Sgntin_row_00107_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00107_00004;
reg                              sign_qin_00107_00004;
wire                             conv_Sgntin_row_00108_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00108_00000;
reg                              sign_qin_00108_00000;
wire                             conv_Sgntin_row_00108_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00108_00001;
reg                              sign_qin_00108_00001;
wire                             conv_Sgntin_row_00108_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00108_00002;
reg                              sign_qin_00108_00002;
wire                             conv_Sgntin_row_00109_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00109_00000;
reg                              sign_qin_00109_00000;
wire                             conv_Sgntin_row_00109_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00109_00001;
reg                              sign_qin_00109_00001;
wire                             conv_Sgntin_row_00109_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00109_00002;
reg                              sign_qin_00109_00002;
wire                             conv_Sgntin_row_00110_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00110_00000;
reg                              sign_qin_00110_00000;
wire                             conv_Sgntin_row_00110_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00110_00001;
reg                              sign_qin_00110_00001;
wire                             conv_Sgntin_row_00110_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00110_00002;
reg                              sign_qin_00110_00002;
wire                             conv_Sgntin_row_00111_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00111_00000;
reg                              sign_qin_00111_00000;
wire                             conv_Sgntin_row_00111_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00111_00001;
reg                              sign_qin_00111_00001;
wire                             conv_Sgntin_row_00111_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00111_00002;
reg                              sign_qin_00111_00002;
wire                             conv_Sgntin_row_00112_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00112_00000;
reg                              sign_qin_00112_00000;
wire                             conv_Sgntin_row_00112_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00112_00001;
reg                              sign_qin_00112_00001;
wire                             conv_Sgntin_row_00112_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00112_00002;
reg                              sign_qin_00112_00002;
wire                             conv_Sgntin_row_00112_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00112_00003;
reg                              sign_qin_00112_00003;
wire                             conv_Sgntin_row_00113_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00113_00000;
reg                              sign_qin_00113_00000;
wire                             conv_Sgntin_row_00113_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00113_00001;
reg                              sign_qin_00113_00001;
wire                             conv_Sgntin_row_00113_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00113_00002;
reg                              sign_qin_00113_00002;
wire                             conv_Sgntin_row_00113_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00113_00003;
reg                              sign_qin_00113_00003;
wire                             conv_Sgntin_row_00114_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00114_00000;
reg                              sign_qin_00114_00000;
wire                             conv_Sgntin_row_00114_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00114_00001;
reg                              sign_qin_00114_00001;
wire                             conv_Sgntin_row_00114_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00114_00002;
reg                              sign_qin_00114_00002;
wire                             conv_Sgntin_row_00114_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00114_00003;
reg                              sign_qin_00114_00003;
wire                             conv_Sgntin_row_00115_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00115_00000;
reg                              sign_qin_00115_00000;
wire                             conv_Sgntin_row_00115_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00115_00001;
reg                              sign_qin_00115_00001;
wire                             conv_Sgntin_row_00115_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00115_00002;
reg                              sign_qin_00115_00002;
wire                             conv_Sgntin_row_00115_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00115_00003;
reg                              sign_qin_00115_00003;
wire                             conv_Sgntin_row_00116_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00116_00000;
reg                              sign_qin_00116_00000;
wire                             conv_Sgntin_row_00116_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00116_00001;
reg                              sign_qin_00116_00001;
wire                             conv_Sgntin_row_00116_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00116_00002;
reg                              sign_qin_00116_00002;
wire                             conv_Sgntin_row_00117_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00117_00000;
reg                              sign_qin_00117_00000;
wire                             conv_Sgntin_row_00117_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00117_00001;
reg                              sign_qin_00117_00001;
wire                             conv_Sgntin_row_00117_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00117_00002;
reg                              sign_qin_00117_00002;
wire                             conv_Sgntin_row_00118_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00118_00000;
reg                              sign_qin_00118_00000;
wire                             conv_Sgntin_row_00118_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00118_00001;
reg                              sign_qin_00118_00001;
wire                             conv_Sgntin_row_00118_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00118_00002;
reg                              sign_qin_00118_00002;
wire                             conv_Sgntin_row_00119_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00119_00000;
reg                              sign_qin_00119_00000;
wire                             conv_Sgntin_row_00119_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00119_00001;
reg                              sign_qin_00119_00001;
wire                             conv_Sgntin_row_00119_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00119_00002;
reg                              sign_qin_00119_00002;
wire                             conv_Sgntin_row_00120_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00120_00000;
reg                              sign_qin_00120_00000;
wire                             conv_Sgntin_row_00120_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00120_00001;
reg                              sign_qin_00120_00001;
wire                             conv_Sgntin_row_00120_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00120_00002;
reg                              sign_qin_00120_00002;
wire                             conv_Sgntin_row_00120_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00120_00003;
reg                              sign_qin_00120_00003;
wire                             conv_Sgntin_row_00120_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00120_00004;
reg                              sign_qin_00120_00004;
wire                             conv_Sgntin_row_00121_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00121_00000;
reg                              sign_qin_00121_00000;
wire                             conv_Sgntin_row_00121_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00121_00001;
reg                              sign_qin_00121_00001;
wire                             conv_Sgntin_row_00121_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00121_00002;
reg                              sign_qin_00121_00002;
wire                             conv_Sgntin_row_00121_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00121_00003;
reg                              sign_qin_00121_00003;
wire                             conv_Sgntin_row_00121_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00121_00004;
reg                              sign_qin_00121_00004;
wire                             conv_Sgntin_row_00122_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00122_00000;
reg                              sign_qin_00122_00000;
wire                             conv_Sgntin_row_00122_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00122_00001;
reg                              sign_qin_00122_00001;
wire                             conv_Sgntin_row_00122_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00122_00002;
reg                              sign_qin_00122_00002;
wire                             conv_Sgntin_row_00122_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00122_00003;
reg                              sign_qin_00122_00003;
wire                             conv_Sgntin_row_00122_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00122_00004;
reg                              sign_qin_00122_00004;
wire                             conv_Sgntin_row_00123_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00123_00000;
reg                              sign_qin_00123_00000;
wire                             conv_Sgntin_row_00123_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00123_00001;
reg                              sign_qin_00123_00001;
wire                             conv_Sgntin_row_00123_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00123_00002;
reg                              sign_qin_00123_00002;
wire                             conv_Sgntin_row_00123_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00123_00003;
reg                              sign_qin_00123_00003;
wire                             conv_Sgntin_row_00123_00004;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00123_00004;
reg                              sign_qin_00123_00004;
wire                             conv_Sgntin_row_00124_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00124_00000;
reg                              sign_qin_00124_00000;
wire                             conv_Sgntin_row_00124_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00124_00001;
reg                              sign_qin_00124_00001;
wire                             conv_Sgntin_row_00124_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00124_00002;
reg                              sign_qin_00124_00002;
wire                             conv_Sgntin_row_00125_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00125_00000;
reg                              sign_qin_00125_00000;
wire                             conv_Sgntin_row_00125_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00125_00001;
reg                              sign_qin_00125_00001;
wire                             conv_Sgntin_row_00125_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00125_00002;
reg                              sign_qin_00125_00002;
wire                             conv_Sgntin_row_00126_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00126_00000;
reg                              sign_qin_00126_00000;
wire                             conv_Sgntin_row_00126_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00126_00001;
reg                              sign_qin_00126_00001;
wire                             conv_Sgntin_row_00126_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00126_00002;
reg                              sign_qin_00126_00002;
wire                             conv_Sgntin_row_00127_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00127_00000;
reg                              sign_qin_00127_00000;
wire                             conv_Sgntin_row_00127_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00127_00001;
reg                              sign_qin_00127_00001;
wire                             conv_Sgntin_row_00127_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00127_00002;
reg                              sign_qin_00127_00002;
wire                             conv_Sgntin_row_00128_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00128_00000;
reg                              sign_qin_00128_00000;
wire                             conv_Sgntin_row_00128_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00128_00001;
reg                              sign_qin_00128_00001;
wire                             conv_Sgntin_row_00128_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00128_00002;
reg                              sign_qin_00128_00002;
wire                             conv_Sgntin_row_00128_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00128_00003;
reg                              sign_qin_00128_00003;
wire                             conv_Sgntin_row_00129_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00129_00000;
reg                              sign_qin_00129_00000;
wire                             conv_Sgntin_row_00129_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00129_00001;
reg                              sign_qin_00129_00001;
wire                             conv_Sgntin_row_00129_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00129_00002;
reg                              sign_qin_00129_00002;
wire                             conv_Sgntin_row_00129_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00129_00003;
reg                              sign_qin_00129_00003;
wire                             conv_Sgntin_row_00130_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00130_00000;
reg                              sign_qin_00130_00000;
wire                             conv_Sgntin_row_00130_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00130_00001;
reg                              sign_qin_00130_00001;
wire                             conv_Sgntin_row_00130_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00130_00002;
reg                              sign_qin_00130_00002;
wire                             conv_Sgntin_row_00130_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00130_00003;
reg                              sign_qin_00130_00003;
wire                             conv_Sgntin_row_00131_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00131_00000;
reg                              sign_qin_00131_00000;
wire                             conv_Sgntin_row_00131_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00131_00001;
reg                              sign_qin_00131_00001;
wire                             conv_Sgntin_row_00131_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00131_00002;
reg                              sign_qin_00131_00002;
wire                             conv_Sgntin_row_00131_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00131_00003;
reg                              sign_qin_00131_00003;
wire                             conv_Sgntin_row_00132_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00132_00000;
reg                              sign_qin_00132_00000;
wire                             conv_Sgntin_row_00132_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00132_00001;
reg                              sign_qin_00132_00001;
wire                             conv_Sgntin_row_00132_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00132_00002;
reg                              sign_qin_00132_00002;
wire                             conv_Sgntin_row_00132_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00132_00003;
reg                              sign_qin_00132_00003;
wire                             conv_Sgntin_row_00133_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00133_00000;
reg                              sign_qin_00133_00000;
wire                             conv_Sgntin_row_00133_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00133_00001;
reg                              sign_qin_00133_00001;
wire                             conv_Sgntin_row_00133_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00133_00002;
reg                              sign_qin_00133_00002;
wire                             conv_Sgntin_row_00133_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00133_00003;
reg                              sign_qin_00133_00003;
wire                             conv_Sgntin_row_00134_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00134_00000;
reg                              sign_qin_00134_00000;
wire                             conv_Sgntin_row_00134_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00134_00001;
reg                              sign_qin_00134_00001;
wire                             conv_Sgntin_row_00134_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00134_00002;
reg                              sign_qin_00134_00002;
wire                             conv_Sgntin_row_00134_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00134_00003;
reg                              sign_qin_00134_00003;
wire                             conv_Sgntin_row_00135_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00135_00000;
reg                              sign_qin_00135_00000;
wire                             conv_Sgntin_row_00135_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00135_00001;
reg                              sign_qin_00135_00001;
wire                             conv_Sgntin_row_00135_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00135_00002;
reg                              sign_qin_00135_00002;
wire                             conv_Sgntin_row_00135_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00135_00003;
reg                              sign_qin_00135_00003;
wire                             conv_Sgntin_row_00136_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00136_00000;
reg                              sign_qin_00136_00000;
wire                             conv_Sgntin_row_00136_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00136_00001;
reg                              sign_qin_00136_00001;
wire                             conv_Sgntin_row_00136_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00136_00002;
reg                              sign_qin_00136_00002;
wire                             conv_Sgntin_row_00136_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00136_00003;
reg                              sign_qin_00136_00003;
wire                             conv_Sgntin_row_00137_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00137_00000;
reg                              sign_qin_00137_00000;
wire                             conv_Sgntin_row_00137_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00137_00001;
reg                              sign_qin_00137_00001;
wire                             conv_Sgntin_row_00137_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00137_00002;
reg                              sign_qin_00137_00002;
wire                             conv_Sgntin_row_00137_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00137_00003;
reg                              sign_qin_00137_00003;
wire                             conv_Sgntin_row_00138_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00138_00000;
reg                              sign_qin_00138_00000;
wire                             conv_Sgntin_row_00138_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00138_00001;
reg                              sign_qin_00138_00001;
wire                             conv_Sgntin_row_00138_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00138_00002;
reg                              sign_qin_00138_00002;
wire                             conv_Sgntin_row_00138_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00138_00003;
reg                              sign_qin_00138_00003;
wire                             conv_Sgntin_row_00139_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00139_00000;
reg                              sign_qin_00139_00000;
wire                             conv_Sgntin_row_00139_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00139_00001;
reg                              sign_qin_00139_00001;
wire                             conv_Sgntin_row_00139_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00139_00002;
reg                              sign_qin_00139_00002;
wire                             conv_Sgntin_row_00139_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00139_00003;
reg                              sign_qin_00139_00003;
wire                             conv_Sgntin_row_00140_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00140_00000;
reg                              sign_qin_00140_00000;
wire                             conv_Sgntin_row_00140_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00140_00001;
reg                              sign_qin_00140_00001;
wire                             conv_Sgntin_row_00140_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00140_00002;
reg                              sign_qin_00140_00002;
wire                             conv_Sgntin_row_00140_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00140_00003;
reg                              sign_qin_00140_00003;
wire                             conv_Sgntin_row_00141_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00141_00000;
reg                              sign_qin_00141_00000;
wire                             conv_Sgntin_row_00141_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00141_00001;
reg                              sign_qin_00141_00001;
wire                             conv_Sgntin_row_00141_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00141_00002;
reg                              sign_qin_00141_00002;
wire                             conv_Sgntin_row_00141_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00141_00003;
reg                              sign_qin_00141_00003;
wire                             conv_Sgntin_row_00142_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00142_00000;
reg                              sign_qin_00142_00000;
wire                             conv_Sgntin_row_00142_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00142_00001;
reg                              sign_qin_00142_00001;
wire                             conv_Sgntin_row_00142_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00142_00002;
reg                              sign_qin_00142_00002;
wire                             conv_Sgntin_row_00142_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00142_00003;
reg                              sign_qin_00142_00003;
wire                             conv_Sgntin_row_00143_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00143_00000;
reg                              sign_qin_00143_00000;
wire                             conv_Sgntin_row_00143_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00143_00001;
reg                              sign_qin_00143_00001;
wire                             conv_Sgntin_row_00143_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00143_00002;
reg                              sign_qin_00143_00002;
wire                             conv_Sgntin_row_00143_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00143_00003;
reg                              sign_qin_00143_00003;
wire                             conv_Sgntin_row_00144_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00144_00000;
reg                              sign_qin_00144_00000;
wire                             conv_Sgntin_row_00144_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00144_00001;
reg                              sign_qin_00144_00001;
wire                             conv_Sgntin_row_00144_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00144_00002;
reg                              sign_qin_00144_00002;
wire                             conv_Sgntin_row_00144_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00144_00003;
reg                              sign_qin_00144_00003;
wire                             conv_Sgntin_row_00145_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00145_00000;
reg                              sign_qin_00145_00000;
wire                             conv_Sgntin_row_00145_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00145_00001;
reg                              sign_qin_00145_00001;
wire                             conv_Sgntin_row_00145_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00145_00002;
reg                              sign_qin_00145_00002;
wire                             conv_Sgntin_row_00145_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00145_00003;
reg                              sign_qin_00145_00003;
wire                             conv_Sgntin_row_00146_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00146_00000;
reg                              sign_qin_00146_00000;
wire                             conv_Sgntin_row_00146_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00146_00001;
reg                              sign_qin_00146_00001;
wire                             conv_Sgntin_row_00146_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00146_00002;
reg                              sign_qin_00146_00002;
wire                             conv_Sgntin_row_00146_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00146_00003;
reg                              sign_qin_00146_00003;
wire                             conv_Sgntin_row_00147_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00147_00000;
reg                              sign_qin_00147_00000;
wire                             conv_Sgntin_row_00147_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00147_00001;
reg                              sign_qin_00147_00001;
wire                             conv_Sgntin_row_00147_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00147_00002;
reg                              sign_qin_00147_00002;
wire                             conv_Sgntin_row_00147_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00147_00003;
reg                              sign_qin_00147_00003;
wire                             conv_Sgntin_row_00148_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00148_00000;
reg                              sign_qin_00148_00000;
wire                             conv_Sgntin_row_00148_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00148_00001;
reg                              sign_qin_00148_00001;
wire                             conv_Sgntin_row_00148_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00148_00002;
reg                              sign_qin_00148_00002;
wire                             conv_Sgntin_row_00149_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00149_00000;
reg                              sign_qin_00149_00000;
wire                             conv_Sgntin_row_00149_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00149_00001;
reg                              sign_qin_00149_00001;
wire                             conv_Sgntin_row_00149_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00149_00002;
reg                              sign_qin_00149_00002;
wire                             conv_Sgntin_row_00150_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00150_00000;
reg                              sign_qin_00150_00000;
wire                             conv_Sgntin_row_00150_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00150_00001;
reg                              sign_qin_00150_00001;
wire                             conv_Sgntin_row_00150_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00150_00002;
reg                              sign_qin_00150_00002;
wire                             conv_Sgntin_row_00151_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00151_00000;
reg                              sign_qin_00151_00000;
wire                             conv_Sgntin_row_00151_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00151_00001;
reg                              sign_qin_00151_00001;
wire                             conv_Sgntin_row_00151_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00151_00002;
reg                              sign_qin_00151_00002;
wire                             conv_Sgntin_row_00152_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00152_00000;
reg                              sign_qin_00152_00000;
wire                             conv_Sgntin_row_00152_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00152_00001;
reg                              sign_qin_00152_00001;
wire                             conv_Sgntin_row_00152_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00152_00002;
reg                              sign_qin_00152_00002;
wire                             conv_Sgntin_row_00152_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00152_00003;
reg                              sign_qin_00152_00003;
wire                             conv_Sgntin_row_00153_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00153_00000;
reg                              sign_qin_00153_00000;
wire                             conv_Sgntin_row_00153_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00153_00001;
reg                              sign_qin_00153_00001;
wire                             conv_Sgntin_row_00153_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00153_00002;
reg                              sign_qin_00153_00002;
wire                             conv_Sgntin_row_00153_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00153_00003;
reg                              sign_qin_00153_00003;
wire                             conv_Sgntin_row_00154_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00154_00000;
reg                              sign_qin_00154_00000;
wire                             conv_Sgntin_row_00154_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00154_00001;
reg                              sign_qin_00154_00001;
wire                             conv_Sgntin_row_00154_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00154_00002;
reg                              sign_qin_00154_00002;
wire                             conv_Sgntin_row_00154_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00154_00003;
reg                              sign_qin_00154_00003;
wire                             conv_Sgntin_row_00155_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00155_00000;
reg                              sign_qin_00155_00000;
wire                             conv_Sgntin_row_00155_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00155_00001;
reg                              sign_qin_00155_00001;
wire                             conv_Sgntin_row_00155_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00155_00002;
reg                              sign_qin_00155_00002;
wire                             conv_Sgntin_row_00155_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00155_00003;
reg                              sign_qin_00155_00003;
wire                             conv_Sgntin_row_00156_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00156_00000;
reg                              sign_qin_00156_00000;
wire                             conv_Sgntin_row_00156_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00156_00001;
reg                              sign_qin_00156_00001;
wire                             conv_Sgntin_row_00156_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00156_00002;
reg                              sign_qin_00156_00002;
wire                             conv_Sgntin_row_00156_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00156_00003;
reg                              sign_qin_00156_00003;
wire                             conv_Sgntin_row_00157_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00157_00000;
reg                              sign_qin_00157_00000;
wire                             conv_Sgntin_row_00157_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00157_00001;
reg                              sign_qin_00157_00001;
wire                             conv_Sgntin_row_00157_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00157_00002;
reg                              sign_qin_00157_00002;
wire                             conv_Sgntin_row_00157_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00157_00003;
reg                              sign_qin_00157_00003;
wire                             conv_Sgntin_row_00158_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00158_00000;
reg                              sign_qin_00158_00000;
wire                             conv_Sgntin_row_00158_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00158_00001;
reg                              sign_qin_00158_00001;
wire                             conv_Sgntin_row_00158_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00158_00002;
reg                              sign_qin_00158_00002;
wire                             conv_Sgntin_row_00158_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00158_00003;
reg                              sign_qin_00158_00003;
wire                             conv_Sgntin_row_00159_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00159_00000;
reg                              sign_qin_00159_00000;
wire                             conv_Sgntin_row_00159_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00159_00001;
reg                              sign_qin_00159_00001;
wire                             conv_Sgntin_row_00159_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00159_00002;
reg                              sign_qin_00159_00002;
wire                             conv_Sgntin_row_00159_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00159_00003;
reg                              sign_qin_00159_00003;
wire                             conv_Sgntin_row_00160_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00160_00000;
reg                              sign_qin_00160_00000;
wire                             conv_Sgntin_row_00160_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00160_00001;
reg                              sign_qin_00160_00001;
wire                             conv_Sgntin_row_00160_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00160_00002;
reg                              sign_qin_00160_00002;
wire                             conv_Sgntin_row_00160_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00160_00003;
reg                              sign_qin_00160_00003;
wire                             conv_Sgntin_row_00161_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00161_00000;
reg                              sign_qin_00161_00000;
wire                             conv_Sgntin_row_00161_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00161_00001;
reg                              sign_qin_00161_00001;
wire                             conv_Sgntin_row_00161_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00161_00002;
reg                              sign_qin_00161_00002;
wire                             conv_Sgntin_row_00161_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00161_00003;
reg                              sign_qin_00161_00003;
wire                             conv_Sgntin_row_00162_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00162_00000;
reg                              sign_qin_00162_00000;
wire                             conv_Sgntin_row_00162_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00162_00001;
reg                              sign_qin_00162_00001;
wire                             conv_Sgntin_row_00162_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00162_00002;
reg                              sign_qin_00162_00002;
wire                             conv_Sgntin_row_00162_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00162_00003;
reg                              sign_qin_00162_00003;
wire                             conv_Sgntin_row_00163_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00163_00000;
reg                              sign_qin_00163_00000;
wire                             conv_Sgntin_row_00163_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00163_00001;
reg                              sign_qin_00163_00001;
wire                             conv_Sgntin_row_00163_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00163_00002;
reg                              sign_qin_00163_00002;
wire                             conv_Sgntin_row_00163_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00163_00003;
reg                              sign_qin_00163_00003;
wire                             conv_Sgntin_row_00164_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00164_00000;
reg                              sign_qin_00164_00000;
wire                             conv_Sgntin_row_00164_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00164_00001;
reg                              sign_qin_00164_00001;
wire                             conv_Sgntin_row_00164_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00164_00002;
reg                              sign_qin_00164_00002;
wire                             conv_Sgntin_row_00164_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00164_00003;
reg                              sign_qin_00164_00003;
wire                             conv_Sgntin_row_00165_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00165_00000;
reg                              sign_qin_00165_00000;
wire                             conv_Sgntin_row_00165_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00165_00001;
reg                              sign_qin_00165_00001;
wire                             conv_Sgntin_row_00165_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00165_00002;
reg                              sign_qin_00165_00002;
wire                             conv_Sgntin_row_00165_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00165_00003;
reg                              sign_qin_00165_00003;
wire                             conv_Sgntin_row_00166_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00166_00000;
reg                              sign_qin_00166_00000;
wire                             conv_Sgntin_row_00166_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00166_00001;
reg                              sign_qin_00166_00001;
wire                             conv_Sgntin_row_00166_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00166_00002;
reg                              sign_qin_00166_00002;
wire                             conv_Sgntin_row_00166_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00166_00003;
reg                              sign_qin_00166_00003;
wire                             conv_Sgntin_row_00167_00000;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00167_00000;
reg                              sign_qin_00167_00000;
wire                             conv_Sgntin_row_00167_00001;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00167_00001;
reg                              sign_qin_00167_00001;
wire                             conv_Sgntin_row_00167_00002;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00167_00002;
reg                              sign_qin_00167_00002;
wire                             conv_Sgntin_row_00167_00003;
reg   [MAX_SUM_WDTH_L-1:0]       conv_qin_00167_00003;
reg                              sign_qin_00167_00003;







/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ic93835a022c46b7aa00a465c407d7da2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I2e30088bf29cedd7debc15b1e6ec4ada;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I38f512bfb84094d1e92a10a345d5505f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I1e878f00f056f637625cb013a93325a8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I25db27464b31fee41ccd7a3cfe4d403e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I19417a224c5cdf1211e9790aa29c4c5c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I16dcafa854ea9c67d8a080feb2ba9166;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I7f63338eee2663fbe61fffd248433310;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Icb1e3c56c8729c32d43c69710e345db2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I6ece8e3c1e89613879336936f77d732f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I72a646ae7e32a16af0f5930a6e95b36a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I7e72d119dd93a6ab05a23fde0a865866;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Ied4fdf5805039cd2fcd042fd13755fdc;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00013;
reg  [MAX_SUM_WDTH_L-1:0]        Id44c2293b765cff450dd1d747c47c1f3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00014;
reg  [MAX_SUM_WDTH_L-1:0]        I8f4ed02f7aeb823b745040f7f3f43ac7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00015;
reg  [MAX_SUM_WDTH_L-1:0]        I6488b9b8f405d7d81a4874fab2678102;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00016;
reg  [MAX_SUM_WDTH_L-1:0]        Ifff612d16828ec907a348479e19ddf31;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00017;
reg  [MAX_SUM_WDTH_L-1:0]        I268262076f22bc6b1507bc8f91b98a0a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00018;
reg  [MAX_SUM_WDTH_L-1:0]        If1f732841adb7c0cad1ba37c0f5fd517;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00019;
reg  [MAX_SUM_WDTH_L-1:0]        I0df8a24f31c027756d248c3bd1b9bf7b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00020;
reg  [MAX_SUM_WDTH_L-1:0]        I8ef901e733b12e76412eb36684e2b575;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00000_00021;
reg  [MAX_SUM_WDTH_L-1:0]        Ia48916a02f68b1b8f5fc7fece04677bb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ia37409944d9fdd3b16e7007e13d82a79;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Idd65f149afe9d5f63ddaf34b82b11e95;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00002;
reg  [MAX_SUM_WDTH_L-1:0]        If2886d560854faed32ebd8e33d868973;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I77778118bb3ea900c080754ff4c49c26;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I7292ed752d8741594d757730950feea4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I68cfd7868e061793ee8a41e69e80219b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I667ead814b303fca64ef047bb8246b19;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I4f25c7edb12e868cb5532e42b4ba5133;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I5aed2d82717f359bb5ac5a0ab91b7beb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I92835fd54631deaefa7b214e2c4b9bff;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I67e067da565635fcff166e3a7d0c446b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00011;
reg  [MAX_SUM_WDTH_L-1:0]        Ifdb0f307b1b9458c0487a1574ccc094b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00012;
reg  [MAX_SUM_WDTH_L-1:0]        I5c6b7d143e42fd3b8bcdb7d7ed4da2c2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00013;
reg  [MAX_SUM_WDTH_L-1:0]        Ie679a21d0136a08cc5e6526e9f8d1843;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00014;
reg  [MAX_SUM_WDTH_L-1:0]        I611942a72a5e12f6afaea6bde6699ef6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00015;
reg  [MAX_SUM_WDTH_L-1:0]        Ica9883c97f823a4491cbee5b45c43590;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00016;
reg  [MAX_SUM_WDTH_L-1:0]        I8e6addfc61f5bfb7af74fc2993639565;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00017;
reg  [MAX_SUM_WDTH_L-1:0]        I9d53619f10e2a426f7297bbf7c81158a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00018;
reg  [MAX_SUM_WDTH_L-1:0]        I8a055c27778913287ad951183fa0d4d6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00019;
reg  [MAX_SUM_WDTH_L-1:0]        I8f6ae5c80bb2f50084b5f5ee5ab0ffc3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00020;
reg  [MAX_SUM_WDTH_L-1:0]        I3db8b3a342e8e2f13a448246aa001c2f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00001_00021;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbee0996ea0f5e16b1f711345be7f2ae;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Idb777f1eb4c3cbba103b9b43f948ccf9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Id5e46b1f8844c7587f99d22170581a24;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I67aadabd3cf49456cace7392a1e7a35a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Id5635595d6b7b6dd7e6d510a27ad6702;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Ice783314a4868f0bba8bc3c5e3b65ae4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ib2d9b7f58cf571b904be02e6073f9b94;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I61b6effae91ae4bdcce4550eb5cf0796;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00007;
reg  [MAX_SUM_WDTH_L-1:0]        If5cf6e81b0e3b77f6a45f2555201acc2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I62fae5bf51588f28c3521715b834909d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00009;
reg  [MAX_SUM_WDTH_L-1:0]        If5cbdab78a4cf86b6285a400d0e0ac90;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I6e481cc49441c08bcd9fdcabbe90a000;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I3aa663be3dd604564ef68b9a2b9d7319;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00012;
reg  [MAX_SUM_WDTH_L-1:0]        I8031632ee8700c63c207e2d6a6bdb630;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00013;
reg  [MAX_SUM_WDTH_L-1:0]        If9be2701858da0bdffbf2dff7bcfd7e1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00014;
reg  [MAX_SUM_WDTH_L-1:0]        Ief209532f4cbf1c6a41bea414577f825;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00015;
reg  [MAX_SUM_WDTH_L-1:0]        I1c8953ad3f64f3c3cc506808aad29dab;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00016;
reg  [MAX_SUM_WDTH_L-1:0]        I1b519d88bbf86cfb080a50ea0480a128;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00017;
reg  [MAX_SUM_WDTH_L-1:0]        I5b8258f35d889071109216b464abb2a4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00018;
reg  [MAX_SUM_WDTH_L-1:0]        Id9681d4e0e4d375f9279de115a4337a3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00019;
reg  [MAX_SUM_WDTH_L-1:0]        Ib42144ece00b82debd70011724a29c91;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00020;
reg  [MAX_SUM_WDTH_L-1:0]        Ic5717058a1815f63f164de1b1defe8cb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00002_00021;
reg  [MAX_SUM_WDTH_L-1:0]        Iea41672f012f225d64d9c75b198c812f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I7a070bd014e1d2c5e55e5fcba88a5664;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I4a0a8b28429b708363458c74230b0fc2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00002;
reg  [MAX_SUM_WDTH_L-1:0]        If585e4075ac1740f3b141ae6a50200f7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1a68cf09bb21a1629369fde87f51bea;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I72b8547125d0ad6c1ad39a68b55c818c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ie14ba4a8657740f9a8d057258db2cb09;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I27490a69fb2a1f6f298639254c37cf9e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I49b9c212fbe74a5dd8b087e417296186;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I0a8e6f5cc8b6ea599b7605abe6479bec;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00009;
reg  [MAX_SUM_WDTH_L-1:0]        Ib6d94b34d3886717e4016fec196f277f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Id7e53d36da7171e036ebfc984dbcea6e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I2ec254d80fd0683d782302cf3839559b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbedaef61051d5df82cd6d55e05c80da;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00013;
reg  [MAX_SUM_WDTH_L-1:0]        I501336bb7ba172c05dd5840036e6228c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00014;
reg  [MAX_SUM_WDTH_L-1:0]        I8e5c4c6c63e42054359cee697cc0d026;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00015;
reg  [MAX_SUM_WDTH_L-1:0]        Id3daa6db921871b752bf92366446afcc;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00016;
reg  [MAX_SUM_WDTH_L-1:0]        Id8367ec60787bfad0da8aa76c6ed8ddb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00017;
reg  [MAX_SUM_WDTH_L-1:0]        I533649312ec995f1f9e514c59a8675b1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00018;
reg  [MAX_SUM_WDTH_L-1:0]        I0621d0b2c83e70b4afd65eb9dca4b514;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00019;
reg  [MAX_SUM_WDTH_L-1:0]        I2ae01892a3cd0432618d7280b31daddb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00020;
reg  [MAX_SUM_WDTH_L-1:0]        I5ed8a2f30bd2ea269341c2267ae3fe83;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00003_00021;
reg  [MAX_SUM_WDTH_L-1:0]        I2c819e7f62c0dc0aac650074b203163b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I30e20b58913d6fbe5817e1956ba8e570;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I1b922bed7f3c4a6705f3ce7a885a68cd;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I2f65f0917713ecc8585392d3b557c1bf;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I3301533e7d9e527118a67c462f1b4357;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I52a88bdb1f03da82730f7579b7b5305d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I644c730662b3725d26cd46fb46106104;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I3da3e36c76c4123bec6879bccb39e933;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Iebde55cddc8170f7dd8855ea55eff0ce;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Ie673e2d92a7090b2fa1c5e14a2e03be3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00009;
reg  [MAX_SUM_WDTH_L-1:0]        If90afe75714f8660ad0eb9f9ea06cd6b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Ifd96e3a6e0050c30a4308328cfecb21f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I68b92cc2d83e9a718edd2aea82314016;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00012;
reg  [MAX_SUM_WDTH_L-1:0]        I6bdbb92363f0e072ed04654e9aad17a5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00013;
reg  [MAX_SUM_WDTH_L-1:0]        I87a4267db59b97ef1b9bca8743cb0322;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00014;
reg  [MAX_SUM_WDTH_L-1:0]        I44eacb2bea725efab7c0dd560279f0f8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00015;
reg  [MAX_SUM_WDTH_L-1:0]        I87a2736466c5ee62b7cc55f17e715ffa;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00016;
reg  [MAX_SUM_WDTH_L-1:0]        I7a66c7713ba126fdc24940cd92f7e10b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00017;
reg  [MAX_SUM_WDTH_L-1:0]        I1f11c579f34c41aade41c53f53468057;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00018;
reg  [MAX_SUM_WDTH_L-1:0]        I651a438f70583d476ae10f066e035435;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00019;
reg  [MAX_SUM_WDTH_L-1:0]        Ibdf17fa73794c846e15fe0a915b071e5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00020;
reg  [MAX_SUM_WDTH_L-1:0]        I76d3221fbcefc0ee08655f7ba4919f3c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00021;
reg  [MAX_SUM_WDTH_L-1:0]        I3458f69c90ea8b20b3d1f67e9a13ec2e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00004_00022;
reg  [MAX_SUM_WDTH_L-1:0]        Ia2d6e9e1e92a30c7028af50ddfbb9bf9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I66c91b5133d9812a03daecc0b14211f8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ifb5986949e88167526d9fcfe07b417ca;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Iedada801ca6cd173ee523ef335e91ff6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I4e2722e547586da7565b2d91a7fc91e7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Ib321a8ceda62c64ab25dc1c718301bda;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I58daeebec4873e6c1c07c090ff81235c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I3f103fbbe49c86c9db46129bd4632cab;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Id6697ca17f1bd6ddd112951b9d89a8ea;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I445ede2983c7470b4418a2ec0cbbd5e1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I034e56cd77ee400ed81b78177b202930;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I08edadbd9366786f96b44268d096b4aa;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I8f86a7af86eb04c5df18e09888cdce7b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Ic00d037a11f8a27ab34e4daab8c9c2e6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00013;
reg  [MAX_SUM_WDTH_L-1:0]        I4d95ceccc6c3ad37f13c98339c59e5c4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00014;
reg  [MAX_SUM_WDTH_L-1:0]        I1ea967d377f462a0e06d7d0d4d95b342;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00015;
reg  [MAX_SUM_WDTH_L-1:0]        Ib0feec63123e66bd6ad6935e9b7fa6bf;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00016;
reg  [MAX_SUM_WDTH_L-1:0]        I7d120060ddae9ff8f7206b3ef63eda50;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00017;
reg  [MAX_SUM_WDTH_L-1:0]        Ib47f8f72386e2e65a88fbadd3a705225;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00018;
reg  [MAX_SUM_WDTH_L-1:0]        I4e0efc35346e2934f5bb4c34a4bc5f90;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00019;
reg  [MAX_SUM_WDTH_L-1:0]        I3ca1014802f58087e3434a1e0df19c01;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00020;
reg  [MAX_SUM_WDTH_L-1:0]        I688a3879b7be1544e6f94b4221c03213;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00021;
reg  [MAX_SUM_WDTH_L-1:0]        Ic22988138610c8671ec342f65f34c7ae;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00005_00022;
reg  [MAX_SUM_WDTH_L-1:0]        I0b85fdd83569e5cbb7d71eed50cb32fd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Idf55390c11e5b41ebc2a28e0af109913;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I6b48935ea25672ee9a42f49eae9e519f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I6a9e6c39c20e45773dab7823a7ff9486;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I42907182010c5889ddb7a700ead16525;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Ib6c26f3e3358cc2ed6fbda83eabd4bd3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ia50d85808790790450f87a5246874b3f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Id4a1744702d7808a80bc40697c864765;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I0cf3d2f3e6793a2dcf15949da16ad28d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I90bd9107f4c931fa1ccb92998ea8cdeb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00009;
reg  [MAX_SUM_WDTH_L-1:0]        Ida1c729e6bfcec2c31a92aa9002f2c68;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Ib848feeccd0ea78ebc8ba8368534c3d1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00011;
reg  [MAX_SUM_WDTH_L-1:0]        Icc11970bbae3adcfa33a0e5dba3e78f4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00012;
reg  [MAX_SUM_WDTH_L-1:0]        I86bb4ef4bdd7af8861280ef30fbeeeea;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00013;
reg  [MAX_SUM_WDTH_L-1:0]        I7e0c259c6c7bacdff5edc44a22e005ba;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00014;
reg  [MAX_SUM_WDTH_L-1:0]        I897ddba059b27f7ed009b0cb70cfb46f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00015;
reg  [MAX_SUM_WDTH_L-1:0]        I4496243eb0542a514b551b4d09bffd7d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00016;
reg  [MAX_SUM_WDTH_L-1:0]        Ic931fb08b2e8441321ebdeed84576a0d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00017;
reg  [MAX_SUM_WDTH_L-1:0]        Ieb6af5390b98e893ee05a939c16d2ffd;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00018;
reg  [MAX_SUM_WDTH_L-1:0]        Ic2a54bad4c5a8885dd24b8687c6db0de;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00019;
reg  [MAX_SUM_WDTH_L-1:0]        I6ecbad763d2b48b78a0584beaefc78ee;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00020;
reg  [MAX_SUM_WDTH_L-1:0]        I20556d23c873c71c7ebc8a961bf40251;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00021;
reg  [MAX_SUM_WDTH_L-1:0]        I79012e6351e6320c22437aa216ea4df1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00006_00022;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf74ab9af877d27c3a6f3881f00ddaf1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I843d35db35d7b42a87ce78d3772cec2f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I2b1398b4bfd374d7221b0a68da28e979;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I6f615d6e74b0c02f8e4265523ad16404;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Iae8a98dd4a7cbfbc56c1404b6a2020af;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Iad53375a54d01c559c74981bf279dfb5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I5db1307f922e0c742d7d9f3a79a4a4f3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I9f78172ed5bf73752196f9a8810005f3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00007;
reg  [MAX_SUM_WDTH_L-1:0]        If85a22d670d47f491dd7568d0453ba1d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Ib9e529170b2896e930a839295796fd31;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00009;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7af536846bac40c1f221d1f72c6c25c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Ib0eb61a2cb831dd35ce9850994e7c2da;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I89d338f59960af7a47595d6afa206abc;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Ib3c1176eb8991e3e85855a9fe845c303;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00013;
reg  [MAX_SUM_WDTH_L-1:0]        I93073d05d509b821a743998cf32c58ee;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00014;
reg  [MAX_SUM_WDTH_L-1:0]        Iab6dac1909c1564c3890ffecc13418df;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00015;
reg  [MAX_SUM_WDTH_L-1:0]        I1b75eeb29167a171d89f6e67039436d5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00016;
reg  [MAX_SUM_WDTH_L-1:0]        I3a31adc52a1405555017b2ddf219b407;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00017;
reg  [MAX_SUM_WDTH_L-1:0]        Iaadba89c6a370240fc0758029f7d8db0;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00018;
reg  [MAX_SUM_WDTH_L-1:0]        I4f4a64fb3ced7d9f7ee4513178e9655a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00019;
reg  [MAX_SUM_WDTH_L-1:0]        I0c76ca58f69c91758e755cd581241284;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00020;
reg  [MAX_SUM_WDTH_L-1:0]        I2312bce18958346149c868846e04643b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00021;
reg  [MAX_SUM_WDTH_L-1:0]        I3e154098cb0a48f1c23234f46613f406;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00007_00022;
reg  [MAX_SUM_WDTH_L-1:0]        I1645c1c588bcbf15dd62d47e08b8e139;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00008_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I4c25de66590e1745d37112e08d8c8e2c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00008_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ia03092ac621b8dd1c206fea1e8b0215f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00008_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I5c9bdb033436dc9f6069baca31f24c2d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00008_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I8f07cf4865480f18ad6945974ec2231c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00008_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I4a7119e8862fe4a6a4100dd9ac67dd24;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00008_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Id78fcfc6724a05f46d44d7c3e7d0c756;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00008_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I7cbd9d619623cbabf8ed6b1fece8f012;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00008_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I58951165d251e370b0f3b3fb537aed18;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00008_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I21daac106f526d84cb8fa5239c19499d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00008_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I178029cec3a5d6141abdfa91b91fdbf4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00009_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I96dfb2efbb55a644616e3474ed07c364;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00009_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I7a17d8f0e2d16c441044db68ee037731;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00009_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I2ced9bb3ae6bdc5b5ef2865fb46abf07;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00009_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I89a93384020d93cf4d26b3902e06cd9e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00009_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbb47d29b9a45559c13ffa3b046c66f5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00009_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I0034177eb1049577a3578b371527f34b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00009_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I22d9ea7bb5a1a3405bcd04b9af40fa62;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00009_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I8a632e7a911bf5726fee587189cb6f16;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00009_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I3765afc490b34e8a310998a4ebcff8cb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00009_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I7607e800ae46a96e016b303120da4247;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00010_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I29b2f1fddee5e32f217d25410bcfce4f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00010_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Iba5f8a31a81f6aa06f5e38c03dc6db54;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00010_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ifcb5c907ad503331317599e4e0ce7be8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00010_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I62d6f2ab4ec8b6ecfa544ad4d90eb30b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00010_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Ide65414c51b3cb182c0f2f238903d60a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00010_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I03a8dc2288eaeb619e746990e20cc868;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00010_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Id81c1b44d16ddbcd466382c60fe84986;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00010_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I503d72f4a2fd20dbf35aa27321d2ede7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00010_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Id6595a4cf33062d1f05cbcee2d0685f1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00010_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I83ebdd7331ca8fbcf5250851b346c0b0;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00011_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I7f6ea26cdfe5986065e7b5aa6842cc1c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00011_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Idab1ec32c20f93c4cc1acb38158f92d5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00011_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I0738add83419502e73674ded2f1ad6c7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00011_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I6c93e63a8e5a2dbd598f1565c7323b39;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00011_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I4aa57a9d46371f1680d5f95596f60b5d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00011_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I5369a7203b78951a3c006c2d3b22507c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00011_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ie72a79a6966cf198687b7c8a8bcdeb13;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00011_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Ie917ae4c44ab0f9c2f1747ff0d2a754e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00011_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I0b1a31ccb34a742552c11b1945e23dd8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00011_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I9a65a845cf2eced39050e8481665f557;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00012_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I3b402b35d38a9fde312c89b82297c1a5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00012_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I309fa33562370e339c19e2377e6a6a7a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00012_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I7d06aed81222a030837cad2074c68e19;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00012_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I835cc6af0cd8189035f2441c2e0d3100;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00012_00004;
reg  [MAX_SUM_WDTH_L-1:0]        If6f768d12f04087246a0d65de1aef99b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00013_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie4b180e1e2cadb865b0eaf6509f99dbb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00013_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ie329a11fc3f6f59f6f1790612fde3250;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00013_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Idb7ddbee4076f7bf49177e69f5e4d112;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00013_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I614d66a7dca2d08efdfdc157ca803d5c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00013_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Iea16eb0ab70ebb1bc47ae55e11ced62d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00014_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa8db43284d5bbebaed4f72d65cf9f92;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00014_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I365d9f3e8b2a9890427f07386deeb093;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00014_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I466aaa0b6cde2ade1901797b8c11e32c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00014_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I7057e329a65ab240ed6cfa824307af65;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00014_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I624e50e3457d33d12680eaf8e7c34aa3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00015_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I9f356fd6820c33fdb5baff05a781e192;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00015_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I39b9c7c664fe7017731877d145d55b44;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00015_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ic62ffbb9e58e0d08b0dec24bba1dc6f2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00015_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I8da2a532288fb817e7dc0cb7b4e3761c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00015_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I6a6e559f5c98f846014e8107fea5a5d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00016_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ibef9219f577b1a62dfdd77296fbfb24d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00016_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I52e6688b5bfff75529d18e20b22832ce;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00016_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Iff22c49354eefca0ea3c5959c14b782c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00016_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ie5377bbdb4111ed00356d5b7737102f3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00016_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I55bf0f3379a8c44634b8f0a3d06c049e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00017_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I9bc9541607f4f6aedb686cdde297bcda;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00017_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ia4620554fbb1d81a71a15a846e4be2f5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00017_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb31b35388ba8ba2ecf98449308ee67d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00017_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ia20410fb3d56587f89a54c00b943b305;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00017_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I9d268f3da12e35b9a4229b7340c0f018;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00018_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I2fce29bd666082eedb2fb3ec8b5ae4dd;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00018_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ia1e8b61e2579a90f5c88ded11c7322c2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00018_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I8cf3718ba65b7fed72e3955f190e34d1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00018_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I7e802d300af54d394b4ee041798c0513;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00018_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Id4fd5a4b97cfa1e176a26f3a823c5516;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00019_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Icbf8d4e75fc66c05eb49c5075696fb07;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00019_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I746a7e90adb2f213b75ae12a161aca0d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00019_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Icb1029aaaaed8c698862ea9c5e22132c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00019_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ib93ea7028c172373b53cdafecae32a67;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00019_00004;
reg  [MAX_SUM_WDTH_L-1:0]        If9628275b000e418f3903daebfdace92;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I830202fb6f08f98c7f71893a881bd555;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I6f38bc9359562f57c1603355e9ee312b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I4701b732d59c26e3790a63c1936f9a24;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ib5d28d8f73d17ab6df6a1291e50c04ab;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I81259f391db792339824ad5dd1a0057b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I6f09ac63effe67a86798b9b4e1690664;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I370b4b3a0048a93ba374a40e170c75a3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I3f8476d0aa0ea2439b67ea1a4adf36c5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I35b52dba10a8a5b22b518388fecac82d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00009;
reg  [MAX_SUM_WDTH_L-1:0]        Ic7db274ed18e6fdecf30381a31238777;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I2c4e538a8db759e9799541d9178ec61e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00011;
reg  [MAX_SUM_WDTH_L-1:0]        Ief6d4c3f5ef8663e111ef99347b023f5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Id95e964e5faecb52c72669b0d28a4bf5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00020_00013;
reg  [MAX_SUM_WDTH_L-1:0]        I0fcef4538102ac6d24aa7090d5405afa;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I055019e38eec6badd1739033d43d7d97;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I35c20a6e823da77a870b421eef2e0a95;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I32cc12cdacef1a4ef64577e0fa977f46;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I26b3f2360ca4a8caee61b2f3a3a08267;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I5ef9b7dc0c63e9ca6a5fb5f7ffa06041;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00005;
reg  [MAX_SUM_WDTH_L-1:0]        If881473b05090f40a027d7eeee7f7ed9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I23bd59ab5b038935301396aaf2acefc1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I874386d94dacf84e699d159af1a49836;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I95bfe51a759bf4165168e5e3b99d6b34;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I4ba5b2f9b7ec0937ecd2c9945cf6de87;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I0b08fb8db0e8a1de3d416907c87fe700;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00011;
reg  [MAX_SUM_WDTH_L-1:0]        Ie030d12e5acf9ef4975a17c83b2481c1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7a0e852d3dfcef950804ea0ebb0c80a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00021_00013;
reg  [MAX_SUM_WDTH_L-1:0]        Iaa4c38d030eab2b7899399aa0d7886d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Icce7ff1d652d4d9c2be5ecf679059bbe;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00001;
reg  [MAX_SUM_WDTH_L-1:0]        If816bc5eacaea23443602e575ddf60b8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I3b224a4ded05446cc5300d430bdd1947;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ia5fc5cfb0e52237b407b37a3858fccb5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I92f8ba6e7f8e9b30fb5b6973eb8fd03e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Icdfa60d2a024dd934f7e6639c6cb2c28;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ifff70b976513eaa42b6bd4b80c98611e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Ica12fa8b631b70a6bbe9f6e92bf73ea0;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Ie69c255335760f706c644b115887269b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00009;
reg  [MAX_SUM_WDTH_L-1:0]        Idb06676b41de19bc86eae34c292183d9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Ib21d2306d5ded3406fac754e69a10d20;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00011;
reg  [MAX_SUM_WDTH_L-1:0]        Ib41d1aa2dcf81879976fb8964cbf6f79;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00012;
reg  [MAX_SUM_WDTH_L-1:0]        I5f8f5e246f008b8d8c75f72828337bab;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00022_00013;
reg  [MAX_SUM_WDTH_L-1:0]        Id6625e78da0e14d2eeb19cc8ac6520e0;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I6d9ddc6afa559ac35c042df1a9390ce9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I9334055c7833676469670372d3c5cc31;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I0c97d772c737c6ff85b584bf69ccaf93;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ic6ce97ae85d91dd8a79f3f9d0da375a2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I83ff9a2750b298b0f7c9b6ce13f574af;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I85699a2a05c343a6a9e828af6d445e9e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I51f6e39b24b2554884e381be79f47ff2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I9f65fd05c6929300860c8cbbde5607f2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00008;
reg  [MAX_SUM_WDTH_L-1:0]        If09761d8f06051d4287ee29ac9c9fa19;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I33bfbe0bcca6d32c86b9576577e3f265;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00010;
reg  [MAX_SUM_WDTH_L-1:0]        If2921210b1c05ecbf00af3a2bcb96ef4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00011;
reg  [MAX_SUM_WDTH_L-1:0]        Ib074e38e280474a782da831a3e0028b4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00012;
reg  [MAX_SUM_WDTH_L-1:0]        I507449dde0bc0c8f53a10759436ec731;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00023_00013;
reg  [MAX_SUM_WDTH_L-1:0]        Id55a3e3f2d75baeba71a345fad695c69;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00024_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I20984f43d22671639a7a178ad15aec04;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00024_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I59f88336d6bdd50ded87d353fb5ce3e9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00024_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I488635e3f7ed77ea88199f5bffd4b1d6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00024_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ie6893017d21c050ba10d206854f4a9f4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00024_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Id3f68b4dc0ab60673208b7d2081f3533;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00024_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I433756b944e061a824a89bda241e879f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00024_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I2eb60a922aa4f7482dd92b9351d53a2d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00025_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I0867979e1b159c8ceae548930376f482;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00025_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I4accfbeae8a5ee0dbeab23ef3a116145;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00025_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ic7570b0b7c5bef5758f68562ae4c90f6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00025_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Iceadadc4456881fdeea85934a9bf4d6c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00025_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I7b2b617ae67424f54961eebce42de77e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00025_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I953f0f8af76f89b2d9ab4abf19fb411d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00025_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I915b4736dcb20f831d02e48f4e79f008;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00026_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7eec587348ae1ca1f00c0a3ad10ad27;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00026_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I001a212686304248c8359e5fc01227c0;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00026_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb7554e012c0fc1223c29b759c900666;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00026_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I9aeb9c42b54a05be6bf9b7b88b6860ba;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00026_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I6a5a5966965b0790b906c6fda71aef80;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00026_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ic943083ca65ace6c42d73f4234739a06;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00026_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Id0b321686d4c39621024cf0dd99822dc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00027_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I0839dd3787442f1b79b87e02436bfdce;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00027_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I89e6a9fd97d8aa4dd3b832c3be4697b2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00027_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I93d4157f48b132642752220059861e98;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00027_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I8fc4faa2891d7fd3479ac1f788f481dc;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00027_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I440f30e9cb4bc89233b46ea00b4cbeb4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00027_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I6568bfd8780c11e0b1b049a01f92abd8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00027_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf7dc4da07f9955d5d4c7e1f63f1ad68;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I7ec1a328587b72a39c462083efea0ee0;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Iaf028e7ab4dc77a7649f15d603834b5f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I58db79a8e9f0cd1ded379897ba2f27ae;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I6d3cb4ccb4e51c7e6603d0abd1a082c4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I79f75f49ea8a29d684af396014b2f3ab;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I9c5ecd86bedb189fada40fae9d751a68;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Iad5f06e1989ead7d306c70a3b02cb8f4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00007;
reg  [MAX_SUM_WDTH_L-1:0]        If6d1a410df5a4aea6a01337a6074fbd9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I3bc40a4db14566b5099b14cee5f61135;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I7e683fd8235d7cfbf4ff407a286f07de;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I97afcedf05e588b7976d6005191dc916;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00011;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8d8eec0aaa662adf2837c9b705fce7e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00028_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Icbd765be950123705955e2c5d7ace84b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I706e8f5617cfae1e6fc83db18c8b5fe3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I1dd8f8c7f1b673898096b1f3ae383197;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I10ca8978cf4659265ed25a27d09acc1c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Iec4656b32460def4a608b6b0f6486af9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I5f4475897d1d58965da1b35fe0ef8c01;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ife61469306df3cf220666b187f1496a9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ib49319b9dfa4914f92f423ceaf840014;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I93ff2f879233cac9b9f0dd2f4c082c09;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I44597d694e9c5d29280e503d72a27c8d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I04a19448c5e75af8021ad02d1a708bb0;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I71a3093121c2f19dcd1412b468652fa8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I3ae09c82029c617034fe6aacbe9e94e6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00029_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Ie7af6b3b441f910b000a333afad6c76f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I4d71dfea8407aa5b5cbb991bc4fea963;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I1a082caecc831a90e74674ba35da4183;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Iec1de44616a2354a56ab1f681059d4c5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ie3c2318e64d0e218c3db557404c4aac8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I9a251d50f41e51b1a5cc2475f267e8a0;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I9b5767a49f7b9dcb8fdaea924835033c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I6ca1e6700a19d03621a193c7240bff54;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I931c597ff12bffce581f653346202f83;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Ia3a2c5d59f6340917ca3933c05ba4678;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00009;
reg  [MAX_SUM_WDTH_L-1:0]        Ie83d0a8ee5ed214bc7577467748aaa04;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Iaac29552e5fc65aaf4f0116f917b707c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00011;
reg  [MAX_SUM_WDTH_L-1:0]        Ie2c8eac7204b98139c03b6fbfff9af36;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00030_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Ied7fcdaec662cb3c2f89f131986fa102;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ib16a17d6430570b45a304d847ee2b11c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I42169e454756fe4d1c5f17f2eeb2e091;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I6fde38a3a92e06fa77123e3279813c41;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Id8ee16437e8d6d6da6d37440e04097b6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf249d8e5acced9b064132575f40e001;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I580659084e3d17b48de6b1c66154fcf5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I7a14e45d43ab77b265501902152c8616;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I81ba868784103e0eb05a44d981d4d666;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Ic6b88783957cbaf253648a30b22f6b1c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I4103c218a85a1d08db5c4f4b5686b2e5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I0e6c0958af503e4a120a49d02a432863;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I8f76b31e8f15c0e5fe24dcb723418111;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00031_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Id1457221b58344b60070aa026436df2c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00032_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Icc31966508e03d8869e81d8aeb243705;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00032_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I9dcccf542ba434b6e0fde6f012f98f92;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00032_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I51ccbb824a5e1e340eefd173c4491728;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00032_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7ae1730dcd8bc708bbfcc6a9f97ac66;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00032_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I4714f5c91203fcfa552f0fcf71b87442;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00032_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I3b6d1e84fdd1019249886fa5fe65895b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00033_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ia8a7d4207dbabc7970bf36f3fe74f72d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00033_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I84047457b43ef33874f4550c3b773460;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00033_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I5e51563c3e69beca0b463742e6e5f9ee;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00033_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I6c8d14e31c80811ccab1b6ab09d28089;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00033_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I50b3b7490c9b65b6e662cc86b163a2df;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00033_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I8351a2110a3d73ad8803cf17e3317017;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00034_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I1e6c696951688d581f21ab2302593335;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00034_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9840e28133eebdca0be313552195c7b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00034_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I82812258a8032e273cab7139266be1b6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00034_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I27ab6fd9927518e29ed36d7a7a241498;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00034_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I05b0f33a3808ac53b29d8d8309447650;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00034_00005;
reg  [MAX_SUM_WDTH_L-1:0]        If150ebf242231f0d22c996a71552f6eb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00035_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If2d0a2b58510715e74787cb60719cb5b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00035_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ib6745a6d17034a29501e022bd846bf2f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00035_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Iae09c127dfe86c9f7bdbeff447c777f5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00035_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I742128de6b237ed48e3a7ccd3788f0d7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00035_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Id5e8fda13ba8f6d95d694d0f30da75bb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00035_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I1aa5a04e40f9b1685c77e4d101c3ccf4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00036_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ife1adea26d13bc299bb2de241ad4a6ea;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00036_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ifcf6c761f0f253921710af87ab1d2247;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00036_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I1478e6a9113c124bdc4361908af6643f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00036_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I0afd42151925883835844cf5deef6156;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00036_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I2b4ab0aadffb3a1bb86f45ebc8acf085;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00036_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Iffa867719ba9c31a8756cc5e6bf81147;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00036_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb62b6cb003f0d5549c864075f23d19b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00036_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I3690d101ae99f258cc58b4482cc378c8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00037_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Id597e95ce8a168ab67890085a26870d0;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00037_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I98df60eb8f65641f9cccce4023be905c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00037_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ibcb4fbdee372353b79c460cdeafdfe4e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00037_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I74dbf75966d047a4a9e91c1bc793666f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00037_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I79b8d9f9447c4c1b551ec6c1e8903040;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00037_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ib34b66548621fabe0753223712b1369f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00037_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ie5b3eb4c00bedfaecc3215d43ff28362;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00037_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Icf3a1b0b6dbcf959b44379024f3c4169;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00038_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I918c2bbe7c71f8c6a07b0bad8811f4e7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00038_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Iedd960a21b1c08b4a5293cff200218b3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00038_00002;
reg  [MAX_SUM_WDTH_L-1:0]        If9722c28747df3a59b0ecf8200907e98;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00038_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ib83df72c8b73a333d0699a8bbbec16be;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00038_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Ide3798a77f709a9f694523338b081f70;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00038_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I0a9722a805604433562f85c62b168b96;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00038_00006;
reg  [MAX_SUM_WDTH_L-1:0]        If9480ec13cd538ed03a43e56bd6264a6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00038_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I433ecf86b7704c5552e5fb5cafe0d529;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00039_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I8326f0b2d25139609e2c5e466724f224;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00039_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbe211d9955cdf2810c9003d1fb78074;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00039_00002;
reg  [MAX_SUM_WDTH_L-1:0]        If15e950b569a92b590127d0ca6f20a16;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00039_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I03e0532841ba39eb1d4ae823c4de2f7d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00039_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I1be81a7b73987ee023e396cec87312d1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00039_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I4ce1a767a78673590c4074f3f03bad8d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00039_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I57806bb7da625881e68ae315543f70d6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00039_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I8b0ab476b4790150575abb06bcdce2b3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00040_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I8846a8961b7d557df4fc62dada679c33;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00040_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I7909a0f96a92e93f95023cddc742a5eb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00040_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I43ac4857544c0fb79d04e850435ef673;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00040_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ia6dfa47c465325c1d9fb9b9c5ce08f01;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00040_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I2e9eda5bea0cc3d88359ce8a7a82f21f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00040_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I53ec2486418e41b2ccfa8fd82777eaf0;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00040_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I18387c05cef21970ecbc39c20a87aafb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00040_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I2b23eae78cb925008ad59f45e80e165b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00040_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Ic69eb7677638a90b7a54389d47be46de;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00041_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I8cb9a216f4da7c27f678386cb214c59d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00041_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I48cb720a6323697084ac3bbd8fcadfcb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00041_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8dc3c1885c92cdcce7fcb58d65d03e7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00041_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ic3aa51a5c758405fa6e2dbed707555b2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00041_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I4d418179c859feb8bc7d750416bb1004;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00041_00005;
reg  [MAX_SUM_WDTH_L-1:0]        If207b2adc6f668f85cb76bf54673fe18;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00041_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ib08b8067ea75e210e83526ca4a37217e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00041_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I95b30f641cbf7bec1886643c4468017d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00041_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I1978531a6f8d1d25ee6d404025ec4753;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00042_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I6c9698ba88db16b8d22ccebd58cc541d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00042_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I0d8ac5e09b200a55bf5ba6f834cc9174;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00042_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ib58b7d3d77a54ff1a180c6fa5f1400e6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00042_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Icf6b990098b7ab91800bfcf1e643153c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00042_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Ie4308b9ac6fb6de9329ba02b1eeb0e8a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00042_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I01d4f02a356c51d7e4e1993de0d8eebd;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00042_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I36c351e3641b01cc43e1dd5de0a649e5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00042_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I4fc983e94c5b8f7bafca61fb0d351c08;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00042_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I1fcb82fdf96cda14a55fa6358cb62c1e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00043_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I665e54ea6bdca483149d3b7f3ee42a2b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00043_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I925df2307b5af6d1b166e5435641d3bd;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00043_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I9b14f48aa357d09e460a445da86cdf89;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00043_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I78e94ecb6c92fa8ee24edaff33b6f82d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00043_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I5ebeb9ce5adee72a7c9527ea6d3a3028;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00043_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I90d7b28ec09142ca8086836fc0c5ea0d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00043_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I27d9985415e6d0b117e5a4c2863aa7f8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00043_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Idf9b563e5d10c2bdbcc07e81d74467eb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00043_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Ie351922194483938302ff6cafc477e4a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ifb2da5faf236ca8636677bc1dc35c4db;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ie15825d216685ae241b528fa9c158ff3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Id92c2d8bc61245c0c8e40bec2424c3c8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Icd9fd8d7114b6e894dbee493b6797df6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I29ff688c085f2b18e7a3af969f18af76;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I6d56db9fcfe69dfcd747521a1ff62297;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I2f17f7c79a0118b39a63894917c6affa;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I7350af5d5ee09ad28c459e3674a829ab;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I67b6415c5135e3d6a41d56d98d3f8315;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I4a6fffd8bb7244599383f2aa3a1c8916;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I7dbcd21016231546b76aab175cac9f74;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I9aeff3dc44ed0d0f32518590a900dcc9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00012;
reg  [MAX_SUM_WDTH_L-1:0]        I988b7d5d56d22d2c77c5c8c125129a50;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00013;
reg  [MAX_SUM_WDTH_L-1:0]        Iff35cd97f2a6d37a7861b9cc1a655ef5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00014;
reg  [MAX_SUM_WDTH_L-1:0]        Ifb3f2a1bedfe41c73d198046a2a3f177;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00044_00015;
reg  [MAX_SUM_WDTH_L-1:0]        I37ddc6ccbc188a3eb8c33a501de820be;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ica608f1136da397e2ab61bd4a5d83201;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I80636a3df4541bf29780bcb4d0ee48f9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I9ad99d544187db3cc7090b92c9933a31;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Iaa8a2b6fcd469869efcf0b75ca38e68f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I9a171d2d8eee362a0073ab7b139d3037;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I84cdcba86bc5991feb391003cd7be40b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00006;
reg  [MAX_SUM_WDTH_L-1:0]        If9e5c3a848acce5daf570458f78f6aad;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I73247d4348333f67a491fc607b15af0e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I021c745eee4b85a2cd91d9d8d2b18b2c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I1381c0a0bd28b1c5542992084635b355;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Ie74eeddc21428254a8fc4c3e293b5eb7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00011;
reg  [MAX_SUM_WDTH_L-1:0]        Ib1d0f94258b45de4bfe610086d8990c5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00012;
reg  [MAX_SUM_WDTH_L-1:0]        I138d6d5d60df37870cdbb1d9c51a94af;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00013;
reg  [MAX_SUM_WDTH_L-1:0]        I706378735e63e15c8d5395446ea41db8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00014;
reg  [MAX_SUM_WDTH_L-1:0]        If8680a7fc4f5532a660006bf4ca6a66e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00045_00015;
reg  [MAX_SUM_WDTH_L-1:0]        Ic59d1ff3051a95166c3c2d5a2881221b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I54a551af28c505601cdfaf8faaa94afb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I6a3124c03eb83d41c16704133bd1cfde;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9ee27b9761af611ab96f0010abd47a3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I305436919f84066a22ab1417ebabd737;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I78e63717f436493b756efa32d66cdefd;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ic965ba971642db19ca773eb68dc0b9bf;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I579480a66a5f6331fb46de13090ce888;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I38d78b447217271a63f30f78b424e2ae;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I4c8d7e5474b19a7c63444d0cb6143728;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00009;
reg  [MAX_SUM_WDTH_L-1:0]        Ia4bc4b7414bf31305ec8f63e7eda61e7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbebe287d56c7d627f3ffcf706575e77;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I83867e6ee369fff7e39ef5c8d5398fef;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00012;
reg  [MAX_SUM_WDTH_L-1:0]        I1d40df7dbf99674f987bd06db714a702;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00013;
reg  [MAX_SUM_WDTH_L-1:0]        I92f42789cb81760ff2973e3a5fe915c3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00014;
reg  [MAX_SUM_WDTH_L-1:0]        Idbd5f2a25ab05808721cf9c403017565;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00046_00015;
reg  [MAX_SUM_WDTH_L-1:0]        I7ca5f07d6d3c2a045dfd55ae5214dd65;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I7f4e1445c68abbadce23944b99d206f9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Id9f28016678e5e2127d9f0aa93e0b534;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I6b939c57a8b7c7c51ab43e1b1df12f6a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ic5d0df586d56bf4cb322d4c3ad677385;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I2e287724873cf6761799eaf464ed6302;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7a10cffe31a53aafa1104b97543280b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ieeb089c6a18791a2227c8571913d689a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Ib29b00328971c3cd67209a5ea5b63b0a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I517e0868f2bb9a22c287a1f3eeaad2f3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I2bc9f76469e2a3f9846560ad1975cf54;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I9f089315e435cd69d2929fdd936a8a77;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I9b54c9fb4179423c731217286e329930;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00012;
reg  [MAX_SUM_WDTH_L-1:0]        I82fb41ab743146badfd2e82258afb310;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00013;
reg  [MAX_SUM_WDTH_L-1:0]        I5619b91de99eead78befdcba1c62411e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00014;
reg  [MAX_SUM_WDTH_L-1:0]        I83dd2047dece99cd841b2e7955819d57;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00047_00015;
reg  [MAX_SUM_WDTH_L-1:0]        I8c927e66ccbf4d19f07af5ef9fbfe3fb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00048_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I0793fa8938acdf65486e5582d01b9e5a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00048_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ied68d7ba0ee9974eb33767e737760b4d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00048_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I95ba37056659b29fd4318a68d85445e8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00048_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I08d7051a18f358d08728f1c401c15c47;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00048_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I768b6f55827ac49eb6ac2655e9397be1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00048_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ic66f737fe60c55d4c10e5d72b307a061;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00048_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I5653779f15c6c9b0f3b26927c48d6234;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00048_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Iac550729fc437fd67151fab57134ec88;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00048_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I853b03c5826eedc3c67a2fae7a640212;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00049_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If46a6b47c1c52243cc0bc92d1edb594f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00049_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I75b36a9b429cd657afc8151b9613aca6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00049_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ife682dd9f677da4d27294fb61b141948;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00049_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ic2b6177a9c586b274b68b25584e6df2c;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00049_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I0d23011c4381496a19cced7bf7960546;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00049_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ic5992d5eaeafd5dded641a7d9801e763;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00049_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ic9e7fe68b9045c6c9eb86185b5f5872e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00049_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I51ad746720b5e6e09ab50f0283552f1a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00049_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I0c8964888a1315507f5d71959dd24cf0;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00050_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Id4d4f814a0bb3418cbf70c306acf048f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00050_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Ic91bd7b4bd148e526ca21d4a5ba87be9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00050_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I7959dddc32f0f181b3ba39149afe1016;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00050_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I087263600b5f38be072a4f1db787aea7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00050_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I78d17a56de5cbe08191ef23b9731c485;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00050_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I82f713a43596df3b935d6da6f8041dc2;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00050_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I422987396853a6a39dabb6e7ddbf91fb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00050_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb6556671e104141dd33188ea5fc024d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00050_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Ie42ce76076a2a5e887e0112086012da6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00051_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I4aea430599b9c0702b3bebd5960b5c91;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00051_00001;
reg  [MAX_SUM_WDTH_L-1:0]        Icbe11a3970136e485eee1bc5053e7273;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00051_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I0a7f1ea1719c1f5ff104445a4130a5a8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00051_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I1802d759f26dd919bc315bfd4156238d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00051_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I2148493e253783fad70f4f2807b83008;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00051_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I39e7f78d33aa7f50264908d2efe23634;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00051_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I844be5874def16af98de935019f35fe8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00051_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Iee5172ba70a6e368b4903f9ff1d93471;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00051_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I1f34b473283291e0970879465c005e2f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1e0b5120737a7f4bf845618ccd22239;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I8abec3020ee5358f8768e5595e9992b4;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I6fe683073211a484cb6e3c416b365d9f;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Id7d764da58ade36853e8a45b5ee19dc3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I3cee2fdf353643deac7d6bca20c8fb52;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00005;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9b8f8f0434fe3783c3d8f68fef30e50;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00006;
reg  [MAX_SUM_WDTH_L-1:0]        I68cba8ad7742cbb34d0b1fb16be4a58a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Idcea56657d40e0fdf9a1c2d920938fd6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Ic549ffab8f0ce161a177faa2ffd1326d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I4d463d500f93f74b2724972ec1d62439;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Iba2f362e263953331649c726afa9c481;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00052_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I6a053d931fb030e03d4882856d3bda75;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I27ede93004e0c240efaa56cc8c570910;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I61a11c1711ca10eefea3438722b40bff;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7924c88692cfddf24fb1eff66eacb7e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00003;
reg  [MAX_SUM_WDTH_L-1:0]        Ibcfd01e622f7f5a5156dd9b335b4e5e0;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I7f6f418ea51b4298da8758bda3f6a21b;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I7185da8937449e23abdd0f39a4b3ed7d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Idc3e3ffa31d9b76c7cf9358a5b2e65d7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I31fe8c887c4aff7c69336676cd31aaa1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I59684d5fe6bbb4b54ac097bd25fceef5;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I86a7cd69148f9590ce91d0aa270d6c54;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Iabce1ccdd968980f622f0e137b159d11;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00053_00011;
reg  [MAX_SUM_WDTH_L-1:0]        Iff02977d7b4c733cca1794246f630931;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I9026c904e5ead7ff2994c4f781d61466;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I99d7489ba87c629c6dd9702a9bbfd3c8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Ifaf191e0d00ba6da7019c2efcf08e1d9;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I4c295991fb08c90862a2f3ba6489000a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Iee61d179da125934298400256788cbb8;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00005;
reg  [MAX_SUM_WDTH_L-1:0]        If87c84440426fb24070372dc1d4bf315;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ib9259a807b31c1b7a528d336bfc403ee;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I411c4d909b2a571e685cd703245516d7;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00008;
reg  [MAX_SUM_WDTH_L-1:0]        If8425453cca8fc8623cb85375c4b8a1d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I654b497f62df75fa283127b5de29b1ad;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I2768519342f7b8a1ee40c1d5ac502b66;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00054_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I8e354c1c5ba44fe5430887248ce0c43b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I8970d8a8aea29913e8696c14c153d16e;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00001;
reg  [MAX_SUM_WDTH_L-1:0]        I3555c6e2fd480a6be11549bf95a9b0b1;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00002;
reg  [MAX_SUM_WDTH_L-1:0]        I8d5600a352e8ba4756f917f912fda6dd;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I7e99d73c95e7ae5c3fe07a3c60ef52eb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00004;
reg  [MAX_SUM_WDTH_L-1:0]        I831633aebe5c6a52b98d630205376f3a;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I82e35482de74223be0d2558334ac2dfb;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Iae2a6f9649ef1bb193e4f0ab5ecbc3e3;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00007;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8eca65d791ad2f6e8f4ed244f22ae3d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00008;
reg  [MAX_SUM_WDTH_L-1:0]        Ic24146b01094df9b9ccd455a791f239d;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I1c9031fd54ff9417d44c9fb17dc1fc63;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00010;
reg  [MAX_SUM_WDTH_L-1:0]        Idefa20487bc5ba6daff03e6b327d76c6;
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00055_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I6f984fd9ea27b40ab3afeac8afd29ade;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00056_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I0be92debced4961df5f461fe81e80bf1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00057_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7bdaba4c6601b7146498aea6c9a3e07;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00058_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Id450c0a1cabe087be051fbf4158e6016;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00059_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I656d0d69f6e243746b87ad67764dbc3d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00060_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Iab9d870dc1ad159bbaecb20a9b72f005;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00061_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Id53b60854f19e095c38f2c255dc57f29;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00062_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If9ba44a2e4a8f0b61692fc69ebeb82bd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00063_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ief95e8620a1c8ddfd6df673a3a223bd8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00064_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I61519bc0aa02ed461dbb91851d0ae19e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00065_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie0c11d584811174a66ca221baf87c36b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00066_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If10f4f45ff0fd17541735934ad20f187;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00067_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I445919f07a6fa8654211301a9a6126bd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00068_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I64102b82893352549abd2e2132b19476;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00069_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I1fc1933fe891ac26f35a42a1b242d919;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00070_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I84dfba8bcf8ad3b85f9472fd60d607b5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00071_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I4302fccefe5ee13161f9ad49f9ddf43c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00072_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I59d7153724d3b3805af799692fbe245a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00073_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Id1650d0e39be078027493f58e9bbcbdd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00074_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If40ad4aca8dbb3bf7dde8c2ff2e5b8f2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00075_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie49f173549396caeab1d13da36e37c65;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00076_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I3002a0e0cdf8e79bc7186a876410d106;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00077_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I2b50fa03f584d10e9af3be085a02a12c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00078_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If473d172a7bff5aeae99245bbb72978d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00079_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ib89f7b5625995290a64bcfb143d978ca;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00080_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Iebe0c9b4a87d58a1c55e2ee6b01603c4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00081_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I104411bb641d2445c7e1385a809bb682;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00082_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I47dd28b4ae4f7151aff5bb271e35b716;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00083_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I3a27d5573b748df459b90a5a347f9d09;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00084_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I2dbef85d2b2b95af39c3a98c4e143253;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00085_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I510d39830ae7b0a857ac11baa7c144d3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00086_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I2751a94a66ea4cb44c512df4c509937f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00087_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ic9a003bfb70ac2da6c229fcad09246d4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00088_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I34ed986182a3311a8cb005b3dccc224b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00089_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ic79281755397f6099ff30c5d07d7e6de;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00090_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I8d6559ccc33cbc663584923a55b928b5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00091_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I4f0a4c241844e390318f11899a0f2c5a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00092_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I45fffa266ce3838f82d755b59216a4d6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00093_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I8f0e65f5db47d5460d4ec2172807a3e1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00094_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I34127c0d1af2438e13b6f4709ece80ba;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00095_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I3a67de0e76bbf29d8c77c21865abda2f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00096_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ic64e64aeb754249b868e14311ea19759;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00097_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ic4aa0dc9014c8445f8d9a7723d7263f5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00098_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I47b988d017580bdfe8f443904b1f3aac;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00099_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ica9ff13e8c3850be6c70b0b06c1d9fbf;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00100_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If2efeb489911f295dd7722cb22ea521d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00101_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Iaa16dffcc01e41e6ff17e92bdefe3df5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00102_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8857b9841fbd795a4192976ef7ecc25;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00103_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If12aef69eea28052aa3bdb6ac31af205;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00104_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I0b3c6162ae2b9221738a18a29489887f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00105_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I08211bba29e87faf4079152bcc973e7d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00106_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ibff3da265f1c3f21548f5b019e1a9dc1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00107_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9fa1762d7844b0d781afdfb0771cea9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00108_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ia677d504b9f7fc2698c0345f236428ba;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00109_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Idebce29121c0481df83d755b60ff632c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00110_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Iad2c780a6386674d50cca54d8c4ebd86;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00111_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If1d7944e7c4828ddb91ffea28609cbc7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00112_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I843a68ceb0adab829091f31d0de56eb6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00113_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I59701b9eb54dda2744a79cebe7d73f3b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00114_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If63cf5e8f47e4e51176401f0d954ea23;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00115_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Id09454844b525697de3e3727d89551e4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00116_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I6d1b2ce4368945b56eee7814638471cc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00117_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I6079945faa57335b1c902ccf7f960a70;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00118_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie7752906ac55cf51f3e96e8c0046f1aa;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00119_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I2d7d4135a94f5df949283c043228791f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00120_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I99c75e3d26c5d01f6ae9abcd05407d8c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00121_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I81e6f97621dbfb2fed6fc236005a2b19;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00122_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ieac60532dcfc916a65054e35cf31d6d2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00123_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7eb83ba73e0dc17f69c357b6ca555bf;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00124_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I5139d8a7a099e3c619c60647c15b7420;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00125_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I6ccd2e11ebd5b2de80b120e20650a602;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00126_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie669cebe5fe39e1a841f8dd3c1f6bc57;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00127_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If32acb9fc212c4af34099acf6df2bc5a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00128_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I075ce236a181bf925c8ccce91d9bc8cd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00129_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I541d4e422b999a0dfca44d275178e1d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00130_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I3e02657f3d9f79338cd083ed024bf96c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00131_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ia5e5537405ab8edcc7cd43c86837d43d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00132_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I07ff388e3b6c7288f0f6c35a345023fe;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00133_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I56cb3b3e193ca5068734417fd0ec4e02;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00134_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I5bbf1765d8f81581d0cf31c0bc755fb3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00135_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Iaa1643095e518846cdede4d5a90dff84;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00136_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Iee6e12f4717a3279dd31b874eabae69e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00137_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ic52a9edbbc5283844d2514ea142ca6e2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00138_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ice3e978c8da2a7de5b28542a5589f0a2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00139_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I336a425aed221c85ca80b9a97d21d6b1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00140_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie477c0f3b77bb299ba8b1a410d211ef7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00141_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie62920d089ae762603cd33fbf97d92bb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00142_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I2ca952e4e676537fd5a8fc71ecfa10e9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00143_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Iefd31e7ff3c829c88f60bc89d70afcf7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00144_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Iafa987a413fd8fcacfe872bc0f5bc2d6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00145_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I305c1ea420d666f258e38c5a65847367;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00146_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I9f040c4088bfab72d74e5332e9710d1a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00147_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ia2f41f9778324a06daeb185c736516a4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00148_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Id9778ba5fbdbed4d33a092da6b68c414;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00149_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I27c2c79d0d719c71c8e28218d1174a13;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00150_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I2a9d6a774769b12ae20bc0cee0c36f5c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00151_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I2c567b75f1399c069b95284f4c36b6d1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00152_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If3d3eb609abfd6e315eec803d2e94490;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00153_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I9c58aea7ce986b1d28f5808b347c015d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00154_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Id139c7a783196941100003b6cb0cd1e7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00155_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I524d7614b01460778da3ce98f6aaa3d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00156_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I8acda65f116d5c91cbe2662ac282aa31;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00157_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If67dbe22f8d22b3430215fb0deae8204;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00158_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I9a35cd7512787263abedd6d9913cf507;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00159_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If9cca23469c5e6001650f1f8b1360ae8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00160_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Icc2606ae8f9a3b425225ae7339112b9d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00161_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I34aa1802d24e074ae54563898929abfa;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00162_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Icb85b3464dc40e8504c53c377e889c45;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00163_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie595a7d10b5ac84c0301fb55bebd3680;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00164_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I9c217a672cabc05efbdff218637123ba;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00165_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If20f3780b4af857ffe8083056085517a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00166_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ic2e275bfa8ab3d2002d2aa374ac9bfe2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00167_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Iac5798fd9915b6778700da6a14f6a381;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00168_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ide3204bf317fdfb993410d338085b174;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00169_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ic3a95140fc1029efa17a6557bc977719;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00170_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I647d3a46bb2c7ed0f1ec08760b3858be;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00171_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I4816747af9d9fc8dc85fd831336ec710;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00172_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I1f66c026a5437320bd1f4df2ff71663d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00173_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If347c58c328193f420286ea27a4afa20;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00174_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I7a126c8304be920f2a920315dc61ba7f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00175_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I237327d6a74df1fb05537dc3691ebf11;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00176_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I64a3e8bb4c87b066806d33a5306a2c53;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00177_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbca6ec39234473fb517447a8beacafc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00178_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I78327356176a16fc996188b83b058cbc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00179_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ifec496c87a7a2474855067305ac8cba3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00180_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I41584165a62caaa37ddebbf79bb8b617;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00181_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Idf0916d6b025aad6eccb98ada5ba3aca;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00182_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I00ef133d5a53f8f99f35b50327e5272b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00183_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I6f0e302d38d75982d0761e306ce9f146;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00184_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I127eed5de00e10a020717e796de76c7d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00185_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If9aad73aefb1b225f35e8c813b85fe87;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00186_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I00a89ac37676521a081a21b1ec1a0798;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00187_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I06f3a34f2b1770ef82ddc2a732b3d4fb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00188_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I4744d64a746f16004e3bedaaa41465f1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00189_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ifae0cc6cc1c65d24bbe84c4ba938e2ea;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00190_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I1223c21129382d41e4f38ef4bbe60c2f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00191_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I14e36e16df00adcd7dc1973d3852d2d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00192_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I0d05ae27b53fb6939e4c2f862a8d20b2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00193_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I97a6fcc08929c3b7d15e36d7706ed13d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00194_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I1f04e86bf27596718836d0a09adbe120;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00195_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie40873cfd6d10a61a94a761becf588a8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00196_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I61960ed74fee948cc12bd1fd8384559a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00197_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I8533a3ec4be4c49166184c94761eaebc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00198_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I00be319b5bdb85ffaf3bb0eca0b348b6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00199_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ie889c916b5af185b52ff5e2e3cc23045;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00200_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I89697be6dcb2e7f972db498c1b1dea71;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00201_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If13dfbfff7cd8e197bb44006a3db73bf;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00202_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I87ed6c3e172c7a06bf6aefe7bf718d70;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00203_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I0db87adc849839fab3a4c9884d5a4882;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00204_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I535e01a6c35fd7b455e4b79b1d4bb414;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00205_00000;
reg  [MAX_SUM_WDTH_L-1:0]        Ia2d1c752cc4b405adb97a815e90a7b96;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00206_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I9ac12eb3878f6fc7dc428fe5e7f35d97;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        wire_qout_00207_00000;
reg  [MAX_SUM_WDTH_L-1:0]        If46fa11dfadb0691eaaa0a40836e08d8;


reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00000;
wire                             tmp_bit_0;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00001;
wire                             tmp_bit_1;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00002;
wire                             tmp_bit_2;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00003;
wire                             tmp_bit_3;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00004;
wire                             tmp_bit_4;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00005;
wire                             tmp_bit_5;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00006;
wire                             tmp_bit_6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00007;
wire                             tmp_bit_7;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00008;
wire                             tmp_bit_8;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00009;
wire                             tmp_bit_9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00010;
wire                             tmp_bit_10;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00011;
wire                             tmp_bit_11;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00012;
wire                             tmp_bit_12;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00013;
wire                             tmp_bit_13;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00014;
wire                             tmp_bit_14;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00015;
wire                             tmp_bit_15;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00016;
wire                             tmp_bit_16;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00017;
wire                             tmp_bit_17;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00018;
wire                             tmp_bit_18;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00019;
wire                             tmp_bit_19;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00020;
wire                             tmp_bit_20;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00021;
wire                             tmp_bit_21;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00022;
wire                             tmp_bit_22;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00023;
wire                             tmp_bit_23;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00024;
wire                             tmp_bit_24;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00025;
wire                             tmp_bit_25;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00026;
wire                             tmp_bit_26;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00027;
wire                             tmp_bit_27;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00028;
wire                             tmp_bit_28;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00029;
wire                             tmp_bit_29;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00030;
wire                             tmp_bit_30;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00031;
wire                             tmp_bit_31;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00032;
wire                             tmp_bit_32;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00033;
wire                             tmp_bit_33;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00034;
wire                             tmp_bit_34;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00035;
wire                             tmp_bit_35;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00036;
wire                             tmp_bit_36;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00037;
wire                             tmp_bit_37;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00038;
wire                             tmp_bit_38;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00039;
wire                             tmp_bit_39;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00040;
wire                             tmp_bit_40;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00041;
wire                             tmp_bit_41;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00042;
wire                             tmp_bit_42;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00043;
wire                             tmp_bit_43;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00044;
wire                             tmp_bit_44;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00045;
wire                             tmp_bit_45;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00046;
wire                             tmp_bit_46;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00047;
wire                             tmp_bit_47;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00048;
wire                             tmp_bit_48;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00049;
wire                             tmp_bit_49;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00050;
wire                             tmp_bit_50;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00051;
wire                             tmp_bit_51;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00052;
wire                             tmp_bit_52;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00053;
wire                             tmp_bit_53;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00054;
wire                             tmp_bit_54;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00055;
wire                             tmp_bit_55;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00056;
wire                             tmp_bit_56;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00057;
wire                             tmp_bit_57;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00058;
wire                             tmp_bit_58;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00059;
wire                             tmp_bit_59;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00060;
wire                             tmp_bit_60;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00061;
wire                             tmp_bit_61;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00062;
wire                             tmp_bit_62;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00063;
wire                             tmp_bit_63;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00064;
wire                             tmp_bit_64;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00065;
wire                             tmp_bit_65;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00066;
wire                             tmp_bit_66;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00067;
wire                             tmp_bit_67;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00068;
wire                             tmp_bit_68;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00069;
wire                             tmp_bit_69;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00070;
wire                             tmp_bit_70;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00071;
wire                             tmp_bit_71;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00072;
wire                             tmp_bit_72;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00073;
wire                             tmp_bit_73;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00074;
wire                             tmp_bit_74;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00075;
wire                             tmp_bit_75;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00076;
wire                             tmp_bit_76;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00077;
wire                             tmp_bit_77;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00078;
wire                             tmp_bit_78;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00079;
wire                             tmp_bit_79;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00080;
wire                             tmp_bit_80;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00081;
wire                             tmp_bit_81;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00082;
wire                             tmp_bit_82;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00083;
wire                             tmp_bit_83;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00084;
wire                             tmp_bit_84;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00085;
wire                             tmp_bit_85;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00086;
wire                             tmp_bit_86;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00087;
wire                             tmp_bit_87;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00088;
wire                             tmp_bit_88;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00089;
wire                             tmp_bit_89;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00090;
wire                             tmp_bit_90;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00091;
wire                             tmp_bit_91;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00092;
wire                             tmp_bit_92;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00093;
wire                             tmp_bit_93;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00094;
wire                             tmp_bit_94;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00095;
wire                             tmp_bit_95;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00096;
wire                             tmp_bit_96;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00097;
wire                             tmp_bit_97;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00098;
wire                             tmp_bit_98;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00099;
wire                             tmp_bit_99;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00100;
wire                             tmp_bit_100;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00101;
wire                             tmp_bit_101;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00102;
wire                             tmp_bit_102;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00103;
wire                             tmp_bit_103;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00104;
wire                             tmp_bit_104;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00105;
wire                             tmp_bit_105;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00106;
wire                             tmp_bit_106;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00107;
wire                             tmp_bit_107;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00108;
wire                             tmp_bit_108;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00109;
wire                             tmp_bit_109;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00110;
wire                             tmp_bit_110;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00111;
wire                             tmp_bit_111;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00112;
wire                             tmp_bit_112;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00113;
wire                             tmp_bit_113;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00114;
wire                             tmp_bit_114;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00115;
wire                             tmp_bit_115;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00116;
wire                             tmp_bit_116;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00117;
wire                             tmp_bit_117;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00118;
wire                             tmp_bit_118;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00119;
wire                             tmp_bit_119;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00120;
wire                             tmp_bit_120;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00121;
wire                             tmp_bit_121;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00122;
wire                             tmp_bit_122;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00123;
wire                             tmp_bit_123;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00124;
wire                             tmp_bit_124;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00125;
wire                             tmp_bit_125;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00126;
wire                             tmp_bit_126;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00127;
wire                             tmp_bit_127;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00128;
wire                             tmp_bit_128;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00129;
wire                             tmp_bit_129;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00130;
wire                             tmp_bit_130;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00131;
wire                             tmp_bit_131;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00132;
wire                             tmp_bit_132;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00133;
wire                             tmp_bit_133;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00134;
wire                             tmp_bit_134;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00135;
wire                             tmp_bit_135;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00136;
wire                             tmp_bit_136;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00137;
wire                             tmp_bit_137;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00138;
wire                             tmp_bit_138;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00139;
wire                             tmp_bit_139;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00140;
wire                             tmp_bit_140;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00141;
wire                             tmp_bit_141;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00142;
wire                             tmp_bit_142;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00143;
wire                             tmp_bit_143;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00144;
wire                             tmp_bit_144;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00145;
wire                             tmp_bit_145;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00146;
wire                             tmp_bit_146;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00147;
wire                             tmp_bit_147;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00148;
wire                             tmp_bit_148;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00149;
wire                             tmp_bit_149;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00150;
wire                             tmp_bit_150;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00151;
wire                             tmp_bit_151;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00152;
wire                             tmp_bit_152;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00153;
wire                             tmp_bit_153;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00154;
wire                             tmp_bit_154;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00155;
wire                             tmp_bit_155;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00156;
wire                             tmp_bit_156;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00157;
wire                             tmp_bit_157;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00158;
wire                             tmp_bit_158;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00159;
wire                             tmp_bit_159;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00160;
wire                             tmp_bit_160;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00161;
wire                             tmp_bit_161;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00162;
wire                             tmp_bit_162;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00163;
wire                             tmp_bit_163;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00164;
wire                             tmp_bit_164;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00165;
wire                             tmp_bit_165;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00166;
wire                             tmp_bit_166;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00167;
wire                             tmp_bit_167;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00168;
wire                             tmp_bit_168;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00169;
wire                             tmp_bit_169;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00170;
wire                             tmp_bit_170;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00171;
wire                             tmp_bit_171;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00172;
wire                             tmp_bit_172;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00173;
wire                             tmp_bit_173;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00174;
wire                             tmp_bit_174;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00175;
wire                             tmp_bit_175;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00176;
wire                             tmp_bit_176;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00177;
wire                             tmp_bit_177;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00178;
wire                             tmp_bit_178;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00179;
wire                             tmp_bit_179;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00180;
wire                             tmp_bit_180;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00181;
wire                             tmp_bit_181;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00182;
wire                             tmp_bit_182;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00183;
wire                             tmp_bit_183;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00184;
wire                             tmp_bit_184;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00185;
wire                             tmp_bit_185;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00186;
wire                             tmp_bit_186;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00187;
wire                             tmp_bit_187;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00188;
wire                             tmp_bit_188;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00189;
wire                             tmp_bit_189;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00190;
wire                             tmp_bit_190;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00191;
wire                             tmp_bit_191;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00192;
wire                             tmp_bit_192;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00193;
wire                             tmp_bit_193;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00194;
wire                             tmp_bit_194;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00195;
wire                             tmp_bit_195;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00196;
wire                             tmp_bit_196;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00197;
wire                             tmp_bit_197;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00198;
wire                             tmp_bit_198;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00199;
wire                             tmp_bit_199;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00200;
wire                             tmp_bit_200;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00201;
wire                             tmp_bit_201;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00202;
wire                             tmp_bit_202;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00203;
wire                             tmp_bit_203;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00204;
wire                             tmp_bit_204;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00205;
wire                             tmp_bit_205;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00206;
wire                             tmp_bit_206;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    sum0_00207;
wire                             tmp_bit_207;

reg  [ 0:0]                      sgnprod_00000;
reg  [MAX_SUM_WDTH_L-1:0]        I5033323484d90d6bfbe03749019fc6dd;
wire  [MAX_SUM_WDTH_L-1:0]       I97afe24956b7f87cd431f048202bab67;
wire  [MAX_SUM_WDTH_L-1:0]       I117235e3ac8e68e4c1ab34db1612aba0;
wire  [MAX_SUM_WDTH_L-1:0]       Ifd700cc9d18f99b63f1947f3ae631976;
wire  [MAX_SUM_WDTH_L-1:0]       Ifffbe3d1007fb07a20d3b37902b3ec95;
wire  [MAX_SUM_WDTH_L-1:0]       If5443777169422ea6e1e3f709b970e05;
wire  [MAX_SUM_WDTH_L-1:0]       Ifaf9fc93e4609d818aa46751754c17f1;
wire  [MAX_SUM_WDTH_L-1:0]       I419caf964986c655df84d043badc37c9;
wire  [MAX_SUM_WDTH_L-1:0]       I3095214ac0e6c1323e75ee4ec85e6821;
reg  [ 0:0]                      sgnprod_00001;
reg  [MAX_SUM_WDTH_L-1:0]        If5dad13ac41b3034bdb034bc86c9b348;
wire  [MAX_SUM_WDTH_L-1:0]       Ided9739bf63937933250a6d0c37535f9;
wire  [MAX_SUM_WDTH_L-1:0]       Id0f139b9f3848b45554ac8429230eea2;
wire  [MAX_SUM_WDTH_L-1:0]       Id9feed58cf9565255abfd0bf7e3ec068;
wire  [MAX_SUM_WDTH_L-1:0]       I30a3be3b5f6ad1880a917eb35659a1bf;
wire  [MAX_SUM_WDTH_L-1:0]       Ie8148d9aa962a733eb65877b902a187d;
wire  [MAX_SUM_WDTH_L-1:0]       I69e98cf3e679183aef6005bb582b18dc;
wire  [MAX_SUM_WDTH_L-1:0]       I7f42a504fc61c9548acebdd8b1858eaa;
wire  [MAX_SUM_WDTH_L-1:0]       I08b1b4639b5a9ca509b943b977f6d4bb;
reg  [ 0:0]                      sgnprod_00002;
reg  [MAX_SUM_WDTH_L-1:0]        Iac428f9f798618e1ef495c626c41892b;
wire  [MAX_SUM_WDTH_L-1:0]       I8d7296627d886566783e79c01b9fa423;
wire  [MAX_SUM_WDTH_L-1:0]       I4fc4c97229a8b1f631a3b505941159e4;
wire  [MAX_SUM_WDTH_L-1:0]       Ib9b16bf51891c328dba2699eb9bcef95;
wire  [MAX_SUM_WDTH_L-1:0]       I6c30501ec81fce286817788d614a7824;
wire  [MAX_SUM_WDTH_L-1:0]       Ia4d4f37baec48121a88808075dd655ef;
wire  [MAX_SUM_WDTH_L-1:0]       I385495ea2bf6442a95ab7561456254ac;
wire  [MAX_SUM_WDTH_L-1:0]       I5128e03d383c226befa6f7422f3a6f04;
wire  [MAX_SUM_WDTH_L-1:0]       Ib208908bab4c20713cd17e20139c8db3;
reg  [ 0:0]                      sgnprod_00003;
reg  [MAX_SUM_WDTH_L-1:0]        I5a6427c8f18b36d2ea18fe60a0831ef1;
wire  [MAX_SUM_WDTH_L-1:0]       Id939992b99a11c09f4688c10ca1a34d1;
wire  [MAX_SUM_WDTH_L-1:0]       I823453ccb90d5b2b2d9dfc6e8358224d;
wire  [MAX_SUM_WDTH_L-1:0]       I279c5c00b92eb1b872b5afa168b0306e;
wire  [MAX_SUM_WDTH_L-1:0]       I66f25b1c3c0eb226295179adcca2c3d2;
wire  [MAX_SUM_WDTH_L-1:0]       I3068627e91b667d14cd3e55a9371931a;
wire  [MAX_SUM_WDTH_L-1:0]       I44c4e0a2d8a7289f8660b81a9ecfa19b;
wire  [MAX_SUM_WDTH_L-1:0]       Ibe868e258dc87f0dd1460ba6b8354671;
wire  [MAX_SUM_WDTH_L-1:0]       Idc3083c3021200345e3edd35a9d4725a;
reg  [ 0:0]                      sgnprod_00004;
reg  [MAX_SUM_WDTH_L-1:0]        Icc29441eac6ca7a138d45743d37505e3;
wire  [MAX_SUM_WDTH_L-1:0]       I320d4f19a5b18c23ff407508d47caa77;
wire  [MAX_SUM_WDTH_L-1:0]       I16becf3c92615d98d5ec51ee9641cc0a;
wire  [MAX_SUM_WDTH_L-1:0]       Ifbfacc3b3a0128119943bcbf80176612;
wire  [MAX_SUM_WDTH_L-1:0]       I6b4f670c9e8e25984e8891f2440322ab;
wire  [MAX_SUM_WDTH_L-1:0]       I19bf0990a30c72421f231772b8627e8e;
wire  [MAX_SUM_WDTH_L-1:0]       I3ec3eb096ebe3ee8a47e1cba6487b997;
wire  [MAX_SUM_WDTH_L-1:0]       I7379ef16405c461ac44b66c4315df831;
wire  [MAX_SUM_WDTH_L-1:0]       I79db45b23d21d533a1f9a6e8f94d403d;
wire  [MAX_SUM_WDTH_L-1:0]       I0979534730cc2b53547d413dbb6b75f4;
wire  [MAX_SUM_WDTH_L-1:0]       I5aa2f9c0667d1a6e871efbd4d2bad3a8;
reg  [ 0:0]                      sgnprod_00005;
reg  [MAX_SUM_WDTH_L-1:0]        I0e7754dcbc04a4850e052ae4a2fbe328;
wire  [MAX_SUM_WDTH_L-1:0]       Iadb28dc990ccf2dd3099544de16b8f16;
wire  [MAX_SUM_WDTH_L-1:0]       I1f71aebf698788d6ada66891e9ea756f;
wire  [MAX_SUM_WDTH_L-1:0]       Ib234e9cf7e7616a1ebc6ab99df2a7ccb;
wire  [MAX_SUM_WDTH_L-1:0]       I297d1edcc583ea4d69da780150f0620c;
wire  [MAX_SUM_WDTH_L-1:0]       Ib0a717cbb4fe38a3fc85520ca0826fd9;
wire  [MAX_SUM_WDTH_L-1:0]       I037ecd5945b1f1280b4469d73fe1c7ff;
wire  [MAX_SUM_WDTH_L-1:0]       I367ff6b11b884e02a3065fc7fe811e15;
wire  [MAX_SUM_WDTH_L-1:0]       I6fab19692b512166fe9c74b5e987788d;
wire  [MAX_SUM_WDTH_L-1:0]       I04dd73af505f618ccdb209b3cf97ceec;
wire  [MAX_SUM_WDTH_L-1:0]       If8c559905d4120488d431719c4e8ce24;
reg  [ 0:0]                      sgnprod_00006;
reg  [MAX_SUM_WDTH_L-1:0]        Ia30c019ed8ce395556494a92e7b42a92;
wire  [MAX_SUM_WDTH_L-1:0]       I20ed4f6f14e20ce3f0e106d1b7782fcd;
wire  [MAX_SUM_WDTH_L-1:0]       Ib10626ffa126188c5bf1fc8399107b26;
wire  [MAX_SUM_WDTH_L-1:0]       I29007c52357ac7afbda39d72a5bb60af;
wire  [MAX_SUM_WDTH_L-1:0]       I66d367c046611f145e607a90911cf499;
wire  [MAX_SUM_WDTH_L-1:0]       I9c4c2556f6170a8df61d909855a846ed;
wire  [MAX_SUM_WDTH_L-1:0]       I6fadc3e8d995bb4317bf7b4377c3c2c5;
wire  [MAX_SUM_WDTH_L-1:0]       I99b20e911c189e0616f02376ab736e91;
wire  [MAX_SUM_WDTH_L-1:0]       I5793c12f5dbdd8245dbb202d550ca960;
wire  [MAX_SUM_WDTH_L-1:0]       Id0660e9637cad1ce1a73d37188060154;
wire  [MAX_SUM_WDTH_L-1:0]       If5a7af7ca023e1393526e888f4220a44;
reg  [ 0:0]                      sgnprod_00007;
reg  [MAX_SUM_WDTH_L-1:0]        I9799695ea8244992a6694eaf5c8ae64d;
wire  [MAX_SUM_WDTH_L-1:0]       Id043eb50634e803e53adc1168379a5d0;
wire  [MAX_SUM_WDTH_L-1:0]       I1f866dd0b129267550aea1a267d9c91e;
wire  [MAX_SUM_WDTH_L-1:0]       I8c4da05c08210fe33139c3d3e5d75d58;
wire  [MAX_SUM_WDTH_L-1:0]       Ib41f7b823681fdd084b6d8436a407aa8;
wire  [MAX_SUM_WDTH_L-1:0]       Ic5b50a785b7acac7e3be4095aa92e50a;
wire  [MAX_SUM_WDTH_L-1:0]       I3ffbe03796b66d00d47fd918be60ab89;
wire  [MAX_SUM_WDTH_L-1:0]       Ifc92a916da938ef6164db250be635f88;
wire  [MAX_SUM_WDTH_L-1:0]       I8ccd42508ce7d5bd897c2cf0c54caeb3;
wire  [MAX_SUM_WDTH_L-1:0]       I4920e7e82749cc036b58a7cd0a03e327;
wire  [MAX_SUM_WDTH_L-1:0]       Ie1040b2aa91f272e4449c4b5f9f8f575;
reg  [ 0:0]                      sgnprod_00008;
reg  [MAX_SUM_WDTH_L-1:0]        I4524cd664b4cb41f642c675fa484c84b;
wire  [MAX_SUM_WDTH_L-1:0]       I65968fb0f63d52ad96cd8fa270126a1b;
wire  [MAX_SUM_WDTH_L-1:0]       I839ac8ee59f51d4c3de92ba5cb26e788;
wire  [MAX_SUM_WDTH_L-1:0]       I33cd95f1919318a0f3df5df7310d64c6;
wire  [MAX_SUM_WDTH_L-1:0]       I4933e8d16fba26cd797b25a9ac2a2de8;
wire  [MAX_SUM_WDTH_L-1:0]       I218f7578eb748e31d0002052f30c5842;
wire  [MAX_SUM_WDTH_L-1:0]       I2a808d1c42ad758ae3baaaee8129dfb2;
wire  [MAX_SUM_WDTH_L-1:0]       I4e851fd3c114af87f5e8c68c02594e3a;
wire  [MAX_SUM_WDTH_L-1:0]       I0da40f88adc46e90f616acdcdb8e0e2c;
reg  [ 0:0]                      sgnprod_00009;
reg  [MAX_SUM_WDTH_L-1:0]        I64e959d80af111ed2fcd54a5407d21bf;
wire  [MAX_SUM_WDTH_L-1:0]       I0dee7767e472a5fd71250ae6c57cc8b5;
wire  [MAX_SUM_WDTH_L-1:0]       I9f40be7552b3dd625e5bce0befc5a548;
wire  [MAX_SUM_WDTH_L-1:0]       I8fdf98ffd757c8845ed6ffa4ddd1a16b;
wire  [MAX_SUM_WDTH_L-1:0]       I8103b777314a4fa471e0898fde9cde08;
wire  [MAX_SUM_WDTH_L-1:0]       If6c3ee8e0d7dea58043d5be0f4630873;
wire  [MAX_SUM_WDTH_L-1:0]       I711a5171f591f472cdbfc9a0f5e1aa17;
wire  [MAX_SUM_WDTH_L-1:0]       Ic30bc38184dfbbd694af52640692709d;
wire  [MAX_SUM_WDTH_L-1:0]       I422f6fd1d273a3834d04b04ab8e2812d;
reg  [ 0:0]                      sgnprod_00010;
reg  [MAX_SUM_WDTH_L-1:0]        I3e0da4bcbab4804b5397fb3aa2c94f51;
wire  [MAX_SUM_WDTH_L-1:0]       Ia0fdc60b90ad18b6585ec1ad4e89e80b;
wire  [MAX_SUM_WDTH_L-1:0]       I7809fe7a30d041a7e569ffe890242df8;
wire  [MAX_SUM_WDTH_L-1:0]       I672b14ec1b3c4797545f266727505a85;
wire  [MAX_SUM_WDTH_L-1:0]       If9620d20ebaae6245a2c386d9bf5fdb1;
wire  [MAX_SUM_WDTH_L-1:0]       Ic74e22bffd88f32eefe499cde0fafa8a;
wire  [MAX_SUM_WDTH_L-1:0]       I76d38ce67387bd76ab45c9cba7d18b31;
wire  [MAX_SUM_WDTH_L-1:0]       I44413c6f6f6493f8a86abf6eb32604f6;
wire  [MAX_SUM_WDTH_L-1:0]       I67f632fca617fe06565ddcaaee8fa8b8;
reg  [ 0:0]                      sgnprod_00011;
reg  [MAX_SUM_WDTH_L-1:0]        I3740b30d31f3c61d93a14a46e3199c4d;
wire  [MAX_SUM_WDTH_L-1:0]       I3fd38a71ce6aa3db1d7a5a9f8a991e12;
wire  [MAX_SUM_WDTH_L-1:0]       I63e5718bf7d8771ef90b91be73d73264;
wire  [MAX_SUM_WDTH_L-1:0]       Ie385e1aeb2b0dcf6d2454be3d7708b27;
wire  [MAX_SUM_WDTH_L-1:0]       Ib2d1b7e105b25b492b45da72536d7578;
wire  [MAX_SUM_WDTH_L-1:0]       I588abf5ef4c583f0fec422736a0ce6a0;
wire  [MAX_SUM_WDTH_L-1:0]       I58bb95c56c7be17c263a2161210d7d8d;
wire  [MAX_SUM_WDTH_L-1:0]       Ifaf0e1f21b3bd7393c475b5126540a72;
wire  [MAX_SUM_WDTH_L-1:0]       I7027db9e0450724a6d417d708f1043f2;
reg  [ 0:0]                      sgnprod_00012;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf0a30abfec9031737eada436ac1a0d4;
wire  [MAX_SUM_WDTH_L-1:0]       Iebcb7206d8860b5094459c5d10b4efed;
wire  [MAX_SUM_WDTH_L-1:0]       I6bbf2b47a7dc50e66a3d8d258d6e31fb;
wire  [MAX_SUM_WDTH_L-1:0]       I8459abaa907f5afcd11884b1ec8c06c5;
wire  [MAX_SUM_WDTH_L-1:0]       Ia16ae2f6ef5000d47b6b84ed058252aa;
wire  [MAX_SUM_WDTH_L-1:0]       Ica32690dbc9ea110fefdce92260b125c;
wire  [MAX_SUM_WDTH_L-1:0]       Ic431d9383cce30b1889c92e2be4cb9d0;
wire  [MAX_SUM_WDTH_L-1:0]       Ib9cca4c0e58373c26d5fd9f51f793898;
wire  [MAX_SUM_WDTH_L-1:0]       I99bf0bc8ac20832b3724b2753f6ca449;
wire  [MAX_SUM_WDTH_L-1:0]       Ie701008f3c60c51ed72c5f964a8fc36e;
wire  [MAX_SUM_WDTH_L-1:0]       I3e2d78f8307a1787f8b2eccba94c7557;
reg  [ 0:0]                      sgnprod_00013;
reg  [MAX_SUM_WDTH_L-1:0]        Id36e8953a02400a5ab1f4dfdb0422e6d;
wire  [MAX_SUM_WDTH_L-1:0]       Ic1b4444ab0df9745d29bf893d9b83168;
wire  [MAX_SUM_WDTH_L-1:0]       I5f52dbf600656a8f5dc6b6b8a45ccebe;
wire  [MAX_SUM_WDTH_L-1:0]       I7f307af79f45ad4b9511e3961c917078;
wire  [MAX_SUM_WDTH_L-1:0]       Ie17a5be2a16d2efb98c976d7ee882535;
wire  [MAX_SUM_WDTH_L-1:0]       I5f19d2adff2f34a4bebe03f929a09c49;
wire  [MAX_SUM_WDTH_L-1:0]       I3cd69aeed9e869a2096d6dced5c209a0;
wire  [MAX_SUM_WDTH_L-1:0]       I359b6a22c9568a13b81670c741281393;
wire  [MAX_SUM_WDTH_L-1:0]       I24ba99614df383c38bbac50ae8b4487e;
wire  [MAX_SUM_WDTH_L-1:0]       I7498bee46de6b1c946ce95fdcc89f6e5;
wire  [MAX_SUM_WDTH_L-1:0]       I0f644f42cabf871b71e5a82871bc7b5d;
reg  [ 0:0]                      sgnprod_00014;
reg  [MAX_SUM_WDTH_L-1:0]        Ica71108a53bfcfd1892b4d03ef68110c;
wire  [MAX_SUM_WDTH_L-1:0]       I71f9e059726a6cac8bdf0efcc0eadd2b;
wire  [MAX_SUM_WDTH_L-1:0]       I0c9b2c1da30bfab514bbb556ae7bd4c4;
wire  [MAX_SUM_WDTH_L-1:0]       I7918b2e37e96aee94fbccca7e0f75fc4;
wire  [MAX_SUM_WDTH_L-1:0]       I76eebd77eb77e0abcbc727d2c511370a;
wire  [MAX_SUM_WDTH_L-1:0]       Ibb2288e62110bae5b2d3fe901974e5c7;
wire  [MAX_SUM_WDTH_L-1:0]       I080f931dfef9d8adfb1dc1ee073eb64c;
wire  [MAX_SUM_WDTH_L-1:0]       Ide1106431e3565158bd81ccd6b18f3a1;
wire  [MAX_SUM_WDTH_L-1:0]       I63df19931e8d28666cccd79922cbd418;
wire  [MAX_SUM_WDTH_L-1:0]       I9a7e4a59447048de90446f877eb06627;
wire  [MAX_SUM_WDTH_L-1:0]       I0917e92ed84363ca92fd2074acd74eba;
reg  [ 0:0]                      sgnprod_00015;
reg  [MAX_SUM_WDTH_L-1:0]        I7c97629ec6e594f9b2160815ddd133cc;
wire  [MAX_SUM_WDTH_L-1:0]       Ie3eefdf7b5561a90a6ddd9e6aa432509;
wire  [MAX_SUM_WDTH_L-1:0]       I56eeb10d11e886cff629457a640a1c76;
wire  [MAX_SUM_WDTH_L-1:0]       I7a9eea89c4e76d856df44b6bdc332840;
wire  [MAX_SUM_WDTH_L-1:0]       If8d8f4333e893788fcb9ec54256e5b7a;
wire  [MAX_SUM_WDTH_L-1:0]       Ie4af0e7e04778d85f5dee73da33376a8;
wire  [MAX_SUM_WDTH_L-1:0]       I019a4e997adf54f5f5ca651f80b7901b;
wire  [MAX_SUM_WDTH_L-1:0]       I10294667f09abbfd4e2f757c414072fc;
wire  [MAX_SUM_WDTH_L-1:0]       Id4e8ab8f15b36bd27d1e4ebc5cbe1495;
wire  [MAX_SUM_WDTH_L-1:0]       I6c93588ca9e7c623d75314da39e89a91;
wire  [MAX_SUM_WDTH_L-1:0]       I1020412efc78d12a9ebcbaeb83e5dcea;
reg  [ 0:0]                      sgnprod_00016;
reg  [MAX_SUM_WDTH_L-1:0]        I4823c8239ace86dc399e906c1b5a0d74;
wire  [MAX_SUM_WDTH_L-1:0]       Id0b574f35a83dcfd4481a10043cd1884;
wire  [MAX_SUM_WDTH_L-1:0]       Ifc577e5c2c7288373a8c5e3969ac1589;
wire  [MAX_SUM_WDTH_L-1:0]       Id18a1a17c1cf6e8a2492aa73b62898f2;
wire  [MAX_SUM_WDTH_L-1:0]       Id8ce8f636723b9f119bb86c25017e6b3;
reg  [ 0:0]                      sgnprod_00017;
reg  [MAX_SUM_WDTH_L-1:0]        I10ad572ca72c2ea991487c39f7eabd7b;
wire  [MAX_SUM_WDTH_L-1:0]       Ic29a18d8d504a2d5280c1d7771346518;
wire  [MAX_SUM_WDTH_L-1:0]       I96a79193aa2956b8f901d5fcc9cf65cf;
wire  [MAX_SUM_WDTH_L-1:0]       I8c97a246c749fbef029f8b1671c772bd;
wire  [MAX_SUM_WDTH_L-1:0]       If9ba9d221909ce7499725f6fd7d519f8;
reg  [ 0:0]                      sgnprod_00018;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9f3fd3a6d16316e55addbe0e336519f;
wire  [MAX_SUM_WDTH_L-1:0]       I53a7878f44253f0f1a82d9d27b1a44c3;
wire  [MAX_SUM_WDTH_L-1:0]       Ie0e928125f9d3d17d123d97e00f1fc34;
wire  [MAX_SUM_WDTH_L-1:0]       I2bd0f77efeca09eebe82ea234e9fe638;
wire  [MAX_SUM_WDTH_L-1:0]       I94f2e7ef9b3463bd598dc9049f6fb0ef;
reg  [ 0:0]                      sgnprod_00019;
reg  [MAX_SUM_WDTH_L-1:0]        I07965bca84276dd56da1af98e64b0adc;
wire  [MAX_SUM_WDTH_L-1:0]       I6dc16510af6b61b79b339d0fce77ac24;
wire  [MAX_SUM_WDTH_L-1:0]       Ic655e213ab81f5d61a018d3ed7016b12;
wire  [MAX_SUM_WDTH_L-1:0]       I2ffc4a604025a2f5c4e273c1d070a725;
wire  [MAX_SUM_WDTH_L-1:0]       I1c76818a9a3b688ca897aa479f7d807f;
reg  [ 0:0]                      sgnprod_00020;
reg  [MAX_SUM_WDTH_L-1:0]        Ic2ade31b8bcf68c4dcc1a371ff14074b;
wire  [MAX_SUM_WDTH_L-1:0]       I3bfee9d3d88f0569010a4e0101200c19;
wire  [MAX_SUM_WDTH_L-1:0]       I5d4738755a26beb6d0f61dd3dec0f804;
wire  [MAX_SUM_WDTH_L-1:0]       I2f3c800091275bcb72d1a2a38fba53f3;
wire  [MAX_SUM_WDTH_L-1:0]       I378e67cca7c4ff6325683f8346963210;
wire  [MAX_SUM_WDTH_L-1:0]       I04c8915a7f4bbde003f7facc84435c1a;
wire  [MAX_SUM_WDTH_L-1:0]       I3f50b10072f38b6addee6845e6df9118;
reg  [ 0:0]                      sgnprod_00021;
reg  [MAX_SUM_WDTH_L-1:0]        Ic0edcf240048fbfde4e938c3e4c5e281;
wire  [MAX_SUM_WDTH_L-1:0]       Icc60eb18ba740036d2a17f98f15cfb98;
wire  [MAX_SUM_WDTH_L-1:0]       I1677daa18aa8b226753b1a887b9420d1;
wire  [MAX_SUM_WDTH_L-1:0]       I36bc2d4c9a4480daa9b0944c08b50738;
wire  [MAX_SUM_WDTH_L-1:0]       I38419a6905f50135a6783aacca0384dd;
wire  [MAX_SUM_WDTH_L-1:0]       Ib48892dcb0715987289662a14672611e;
wire  [MAX_SUM_WDTH_L-1:0]       Icd9c94f929dbc71c9b836fda3019630b;
reg  [ 0:0]                      sgnprod_00022;
reg  [MAX_SUM_WDTH_L-1:0]        I8b42e89ff5f780d4ef8cd1cd5c99ef61;
wire  [MAX_SUM_WDTH_L-1:0]       I5d0249d9a772805b3fba3f3c7f5d35bd;
wire  [MAX_SUM_WDTH_L-1:0]       Ie97341deb6fb24d49eb8b96bd0fd3f35;
wire  [MAX_SUM_WDTH_L-1:0]       I17dd788f9d8e91307b6b1ab7488f9ce2;
wire  [MAX_SUM_WDTH_L-1:0]       I92ae370022ed107b152b10fd0aa3d2b7;
wire  [MAX_SUM_WDTH_L-1:0]       Iebb39f0d19ec1208bbfba6cf67a3bfc7;
wire  [MAX_SUM_WDTH_L-1:0]       I81861f6bb8bbbab6e93407cfb4a852b8;
reg  [ 0:0]                      sgnprod_00023;
reg  [MAX_SUM_WDTH_L-1:0]        I70b1b8521b36920707e95fc9418eb8a9;
wire  [MAX_SUM_WDTH_L-1:0]       I217b2e3ca0a534fc5b1910adf3c1b57d;
wire  [MAX_SUM_WDTH_L-1:0]       I8429b08891dc56af24c72ce1b7725457;
wire  [MAX_SUM_WDTH_L-1:0]       If96747262303f6c5c6b129e39224bd23;
wire  [MAX_SUM_WDTH_L-1:0]       If7012457af15c405baeaa1710319b541;
wire  [MAX_SUM_WDTH_L-1:0]       Ia0a0229ef71b85195352bb664ea4e4e3;
wire  [MAX_SUM_WDTH_L-1:0]       I42aeb7c23accc2ca874c7f8221c3af93;
reg  [ 0:0]                      sgnprod_00024;
reg  [MAX_SUM_WDTH_L-1:0]        I4fb1c32a62cbbaeb585c6564a3c938f9;
wire  [MAX_SUM_WDTH_L-1:0]       I7df6a95bf51f40693c439c6df36510d4;
wire  [MAX_SUM_WDTH_L-1:0]       I8fe65f9c344d7ec8657f192abefc3fb6;
wire  [MAX_SUM_WDTH_L-1:0]       I4d75c95d34d8d8aeeb528456bbe136e1;
wire  [MAX_SUM_WDTH_L-1:0]       I43746054a38c9521f8da9db9d0e91f99;
wire  [MAX_SUM_WDTH_L-1:0]       I0430ac2a4b2b2e2fc7f8154bf946553c;
wire  [MAX_SUM_WDTH_L-1:0]       I25dc807fd55b81c9f24fd0d1edcaa758;
reg  [ 0:0]                      sgnprod_00025;
reg  [MAX_SUM_WDTH_L-1:0]        Iefc37daeec14e14ef2fe0716f73109dc;
wire  [MAX_SUM_WDTH_L-1:0]       I7881184f1779b9fd4fdf329c5f7664da;
wire  [MAX_SUM_WDTH_L-1:0]       I8e6de2d692a307ee8a5a4b2a9265a633;
wire  [MAX_SUM_WDTH_L-1:0]       I54b2b18ab051b468808a3d0fc4bc893f;
wire  [MAX_SUM_WDTH_L-1:0]       I37ee86e2ca32832862cb57efe76bbedf;
wire  [MAX_SUM_WDTH_L-1:0]       Ic95f2fc697574803c0f7fa35c2609f0c;
wire  [MAX_SUM_WDTH_L-1:0]       I933a30c52c9bec5172530b2d739a3b63;
reg  [ 0:0]                      sgnprod_00026;
reg  [MAX_SUM_WDTH_L-1:0]        Ibd15f164f6d2ac9e5721a21464bc2c5c;
wire  [MAX_SUM_WDTH_L-1:0]       I7bbd7df18f85197c22fe8cfe37312af6;
wire  [MAX_SUM_WDTH_L-1:0]       I50d5ada7c91c7af16492c6b41151b68f;
wire  [MAX_SUM_WDTH_L-1:0]       I32c8e7996b3473d4906c40018799a16b;
wire  [MAX_SUM_WDTH_L-1:0]       Ic0eacd5a4812ad7ae3fa251ab2db4694;
wire  [MAX_SUM_WDTH_L-1:0]       Ideecf8ab87d28a840cd93851169ab05b;
wire  [MAX_SUM_WDTH_L-1:0]       I1ac6775eb38457b7962241d2e7336b0d;
reg  [ 0:0]                      sgnprod_00027;
reg  [MAX_SUM_WDTH_L-1:0]        I951dfff9507bb70214d48e03a0ebb3a7;
wire  [MAX_SUM_WDTH_L-1:0]       I2ecaa89698604fddd863d7e28d643a57;
wire  [MAX_SUM_WDTH_L-1:0]       I273e0fe9c51c8549c8dfff393ca2e4e1;
wire  [MAX_SUM_WDTH_L-1:0]       Ifb1fc76002f6920a1f44c7b1bbcd0020;
wire  [MAX_SUM_WDTH_L-1:0]       Idf6d4e3aa753aa396a9bffb27732f851;
wire  [MAX_SUM_WDTH_L-1:0]       If14ca1f5d1c2977f9da79eaebaad1bf9;
wire  [MAX_SUM_WDTH_L-1:0]       If8f1505d9f10e30bd3320f500d34932f;
reg  [ 0:0]                      sgnprod_00028;
reg  [MAX_SUM_WDTH_L-1:0]        Ie78e30b2a2eda75d0df7d10fd67b5e36;
wire  [MAX_SUM_WDTH_L-1:0]       Id32aa77c6406b35a00168bb5452b12fb;
wire  [MAX_SUM_WDTH_L-1:0]       I9a73686acefeb361337511f6943b036b;
wire  [MAX_SUM_WDTH_L-1:0]       Ib6eb7ce5a070f3a87bcf0e18be8c855d;
wire  [MAX_SUM_WDTH_L-1:0]       If69b0b717c35d33fc8c0e59b07eb9edc;
wire  [MAX_SUM_WDTH_L-1:0]       Ibb0d73078b779585e6b0e228391ecb96;
wire  [MAX_SUM_WDTH_L-1:0]       I2894546e399fe3e33d7579772a1310df;
reg  [ 0:0]                      sgnprod_00029;
reg  [MAX_SUM_WDTH_L-1:0]        Ia0b83a372dd4115dc4d61eb8ff0811b9;
wire  [MAX_SUM_WDTH_L-1:0]       I97f99a266267859aed199b278a430417;
wire  [MAX_SUM_WDTH_L-1:0]       Ie18cc792329941a3654322376a937d8d;
wire  [MAX_SUM_WDTH_L-1:0]       Ie914a99f08d60b74c3c36a632a4ca9b0;
wire  [MAX_SUM_WDTH_L-1:0]       I82916e9dc3894ad88e12de01a68d6aa5;
wire  [MAX_SUM_WDTH_L-1:0]       I6cbf576b3d652e34c0221f8316b5a392;
wire  [MAX_SUM_WDTH_L-1:0]       I9141b2516d7f855cd186472780af7b67;
reg  [ 0:0]                      sgnprod_00030;
reg  [MAX_SUM_WDTH_L-1:0]        If5c5bcbbea01aa22f242b913f0d01929;
wire  [MAX_SUM_WDTH_L-1:0]       I07bf32ed72de9c02abf700c64853af61;
wire  [MAX_SUM_WDTH_L-1:0]       I52663a2999fb9571834d517538691b6f;
wire  [MAX_SUM_WDTH_L-1:0]       I8dcb88c94506367aabe8d7ed62cc56c2;
wire  [MAX_SUM_WDTH_L-1:0]       Ie676a4bee61154145391d9cc473fe91d;
wire  [MAX_SUM_WDTH_L-1:0]       I9502c8fbf6b48749bf9f84a89a937dfe;
wire  [MAX_SUM_WDTH_L-1:0]       I0c91e540e7106f32ae59491d8ed1853e;
reg  [ 0:0]                      sgnprod_00031;
reg  [MAX_SUM_WDTH_L-1:0]        Iccba58cd3519fb4cc75a61b50da1d562;
wire  [MAX_SUM_WDTH_L-1:0]       Iddfb8a8e261389eb4a2a10880c19446a;
wire  [MAX_SUM_WDTH_L-1:0]       If0d55f861d4b3f0970c529024ca142d5;
wire  [MAX_SUM_WDTH_L-1:0]       Ib054f5d3f5cbb29a053d0e50c23cb3a8;
wire  [MAX_SUM_WDTH_L-1:0]       I1d65e9f97e93de8cc2a5dd532f8e482a;
wire  [MAX_SUM_WDTH_L-1:0]       I3bdeab8c87325d46e45d9e2d44756934;
wire  [MAX_SUM_WDTH_L-1:0]       If9228f7ecf19c41f4bbd8dabd0d5816c;
reg  [ 0:0]                      sgnprod_00032;
reg  [MAX_SUM_WDTH_L-1:0]        Ibc0999e4d0b3cc2650f9348b8c204b14;
wire  [MAX_SUM_WDTH_L-1:0]       I9e3edee214c4937d2aa462d3cffa624b;
wire  [MAX_SUM_WDTH_L-1:0]       I9fcbbd2e81b006b50e2d35ed2627bf83;
wire  [MAX_SUM_WDTH_L-1:0]       Ie16f3d50ad5e5581ca099549db7232d2;
wire  [MAX_SUM_WDTH_L-1:0]       I6345e93f3fa7f5eb2008dd41742afc2d;
reg  [ 0:0]                      sgnprod_00033;
reg  [MAX_SUM_WDTH_L-1:0]        I2aeff1fb4b839a581acaf26f90f9113c;
wire  [MAX_SUM_WDTH_L-1:0]       I698b93e10073b5d29357cde4bcac9dbe;
wire  [MAX_SUM_WDTH_L-1:0]       Ie7ced910d84655790823e6173a5a314a;
wire  [MAX_SUM_WDTH_L-1:0]       If6e3b6fd1810f6964e9024329d7cb3e3;
wire  [MAX_SUM_WDTH_L-1:0]       If1045908c6d7476bd5507e57d08c406c;
reg  [ 0:0]                      sgnprod_00034;
reg  [MAX_SUM_WDTH_L-1:0]        I7d60d53f883f8187700c4e78b4c22f1c;
wire  [MAX_SUM_WDTH_L-1:0]       I4d4f6705ed77a16ff31b34bae0d8b6d9;
wire  [MAX_SUM_WDTH_L-1:0]       I70a492396580ac1143d8a2f4b181e873;
wire  [MAX_SUM_WDTH_L-1:0]       I2fade32b5bdf245fa15289620dae2670;
wire  [MAX_SUM_WDTH_L-1:0]       Ie0dc166f57fea074496241a32cdb6015;
reg  [ 0:0]                      sgnprod_00035;
reg  [MAX_SUM_WDTH_L-1:0]        Id6fcf4b7af4a37c854a12e2ae80851fa;
wire  [MAX_SUM_WDTH_L-1:0]       If6a2518891412caa6d6d507082501f1e;
wire  [MAX_SUM_WDTH_L-1:0]       Ic9912e5a838a377b26a19d22148a64df;
wire  [MAX_SUM_WDTH_L-1:0]       Ibc0fca22d16444bc17877106ca772c31;
wire  [MAX_SUM_WDTH_L-1:0]       Ie4291d233597d5d676a80fd62d9bd208;
reg  [ 0:0]                      sgnprod_00036;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa5e5f7d753964f14f0f16dbe552fd85;
wire  [MAX_SUM_WDTH_L-1:0]       Ifc13b798d76aa70ec1877c275fb31d36;
wire  [MAX_SUM_WDTH_L-1:0]       I57d6637f0bdab578a790e4a12ccaa16b;
wire  [MAX_SUM_WDTH_L-1:0]       If8ea04fe685b4f20cdaf9a84984d56fe;
wire  [MAX_SUM_WDTH_L-1:0]       Ie0c86f20c28bcbe410b191b90d29bf76;
wire  [MAX_SUM_WDTH_L-1:0]       I3dc5d3f66726e15968a70cbf3d3b656a;
reg  [ 0:0]                      sgnprod_00037;
reg  [MAX_SUM_WDTH_L-1:0]        I900d471b087cf5a436c2ad66a84d8280;
wire  [MAX_SUM_WDTH_L-1:0]       Id674686e7ac37fd6f63846f9a9cede19;
wire  [MAX_SUM_WDTH_L-1:0]       Ie2ed9668d13d219c60f2e0614488cd42;
wire  [MAX_SUM_WDTH_L-1:0]       I98abc995ff89934534543be93c6e3ffa;
wire  [MAX_SUM_WDTH_L-1:0]       I579cf9386ab7b08efa204d735335e462;
wire  [MAX_SUM_WDTH_L-1:0]       I9efa4d729d10a6b7cc335fb765ed032c;
reg  [ 0:0]                      sgnprod_00038;
reg  [MAX_SUM_WDTH_L-1:0]        I6d1434907f0292ea2ee47cbc5b52bfb9;
wire  [MAX_SUM_WDTH_L-1:0]       If9191ebc8e88d4e75f0f35897ebb1421;
wire  [MAX_SUM_WDTH_L-1:0]       I3511287cfe69d5cedc5a8fbcad708437;
wire  [MAX_SUM_WDTH_L-1:0]       I91812179d44cb675b90d477f33ec48ad;
wire  [MAX_SUM_WDTH_L-1:0]       Idb04a1aae91fdc477ca38ed66789ee88;
wire  [MAX_SUM_WDTH_L-1:0]       I566054aece562960590ee28b157e4a3e;
reg  [ 0:0]                      sgnprod_00039;
reg  [MAX_SUM_WDTH_L-1:0]        I938bef7ba7ae1739d8e6a6a7c117a1b1;
wire  [MAX_SUM_WDTH_L-1:0]       I7b2ffb762cd9ef7aa8ba224efb75c46c;
wire  [MAX_SUM_WDTH_L-1:0]       Id90bbb642b0f4434d8a148a28b6b2f65;
wire  [MAX_SUM_WDTH_L-1:0]       Ia4e297e35d484b15adce7e1d67f582b0;
wire  [MAX_SUM_WDTH_L-1:0]       I84996b1d03b692f6f736fb04c7f91e83;
wire  [MAX_SUM_WDTH_L-1:0]       I83078cc7857fc17b30f640854a4d6be5;
reg  [ 0:0]                      sgnprod_00040;
reg  [MAX_SUM_WDTH_L-1:0]        I6384a9416b2d1da01df1b2d7b16c5390;
wire  [MAX_SUM_WDTH_L-1:0]       I94bb467129904032736fb13dd636c600;
wire  [MAX_SUM_WDTH_L-1:0]       Ifa76758b50f439170ecd6d86ff898bc4;
wire  [MAX_SUM_WDTH_L-1:0]       I9d831dd976e8cd5d8f6a6818601e6424;
wire  [MAX_SUM_WDTH_L-1:0]       I474774ae149804412ed4aaf1cdcaba88;
wire  [MAX_SUM_WDTH_L-1:0]       I964cdcb4e6b49a62d30c2a2540851317;
reg  [ 0:0]                      sgnprod_00041;
reg  [MAX_SUM_WDTH_L-1:0]        I5097a79e7cf7a30d38ba198d1407119c;
wire  [MAX_SUM_WDTH_L-1:0]       I6df268bc9f85ce88674a9165664ea84a;
wire  [MAX_SUM_WDTH_L-1:0]       I74fdcbe9f49f7bce1f5e31d956c5883c;
wire  [MAX_SUM_WDTH_L-1:0]       I4a1b8453cb7a21745d5f74ad05653ed2;
wire  [MAX_SUM_WDTH_L-1:0]       I9c53b478b2011fac0615a152fe60d5b6;
wire  [MAX_SUM_WDTH_L-1:0]       Id75dbed8f1a5befda32c60b994681013;
reg  [ 0:0]                      sgnprod_00042;
reg  [MAX_SUM_WDTH_L-1:0]        Ib113c26c8dcf49c972c41a938059a787;
wire  [MAX_SUM_WDTH_L-1:0]       I378a59323b74623c5524f854d6e11226;
wire  [MAX_SUM_WDTH_L-1:0]       I080bf885464a0cc948a4450e9f7d1d26;
wire  [MAX_SUM_WDTH_L-1:0]       If769e73adea227de1fd85c2e89d0ba08;
wire  [MAX_SUM_WDTH_L-1:0]       Ifa6a34b83225e9d9b28b14874c4444e3;
wire  [MAX_SUM_WDTH_L-1:0]       I584b1d4d6fb7ee4f20ad9c96715cdf90;
reg  [ 0:0]                      sgnprod_00043;
reg  [MAX_SUM_WDTH_L-1:0]        I970c4a25a8bce82a9d2846679029fcab;
wire  [MAX_SUM_WDTH_L-1:0]       I265f9b91fbb62164e589dcf96818c4f5;
wire  [MAX_SUM_WDTH_L-1:0]       I3d59a47c88227734cf6fc0d6fd30db11;
wire  [MAX_SUM_WDTH_L-1:0]       I6144b6df2c87ea0948d730343b42129f;
wire  [MAX_SUM_WDTH_L-1:0]       Ia7ca7400e36ea572fba8e19bcc81ecbd;
wire  [MAX_SUM_WDTH_L-1:0]       I302e61b49accf5db556b87517f2341f5;
reg  [ 0:0]                      sgnprod_00044;
reg  [MAX_SUM_WDTH_L-1:0]        Ibe2af096ad2db26e54d8b4b3bb05175c;
wire  [MAX_SUM_WDTH_L-1:0]       I5d9af1abff6efe3a55c6568d936b6ec7;
wire  [MAX_SUM_WDTH_L-1:0]       I8cde0aa611c476b5112edeb8f17f15bf;
wire  [MAX_SUM_WDTH_L-1:0]       Icaa40ec40d6d26cdf70bb5ae7d492e47;
wire  [MAX_SUM_WDTH_L-1:0]       I8346f15d822cacfeecbe5d75412cb53f;
wire  [MAX_SUM_WDTH_L-1:0]       I5ee364aab320ab40c0f65feda6f53b18;
reg  [ 0:0]                      sgnprod_00045;
reg  [MAX_SUM_WDTH_L-1:0]        Ie48569c467fba0c1291f71d6080ebedc;
wire  [MAX_SUM_WDTH_L-1:0]       I1f0ecba054900f96cd7100741191c5f4;
wire  [MAX_SUM_WDTH_L-1:0]       I4faf2caf62966416118a54015908c889;
wire  [MAX_SUM_WDTH_L-1:0]       Idd0329980a36f87859150530ab44b52d;
wire  [MAX_SUM_WDTH_L-1:0]       Ie66bc10dde27f08813d4d347fd7cf6ce;
wire  [MAX_SUM_WDTH_L-1:0]       Ie1d8b3ea7c6603cebf2f9adb776910b7;
reg  [ 0:0]                      sgnprod_00046;
reg  [MAX_SUM_WDTH_L-1:0]        I90e7ded06617b49cdb8b5301fe9c6a20;
wire  [MAX_SUM_WDTH_L-1:0]       Ia37488e9a50cf5cc08de74ade676db96;
wire  [MAX_SUM_WDTH_L-1:0]       I08aa45211cab01d567cd5eb172fd2f0c;
wire  [MAX_SUM_WDTH_L-1:0]       If4ff0c63ec1deb46412858e496451a01;
wire  [MAX_SUM_WDTH_L-1:0]       Ife7bfd15fc4c392b5d2288d9a4e879b3;
wire  [MAX_SUM_WDTH_L-1:0]       I24ac26debafd03c7333d174e8725afd6;
reg  [ 0:0]                      sgnprod_00047;
reg  [MAX_SUM_WDTH_L-1:0]        I4920014f5d017f4e840dc3b88526955f;
wire  [MAX_SUM_WDTH_L-1:0]       I99d80ad68e2563d0f78a0e3bb82c5328;
wire  [MAX_SUM_WDTH_L-1:0]       I9943733ef305983c629565c881054bbf;
wire  [MAX_SUM_WDTH_L-1:0]       I7cb4420bc55c03a6500f5228d31fe43c;
wire  [MAX_SUM_WDTH_L-1:0]       Ic4d19dec464359c0a9fa75148fe90c73;
wire  [MAX_SUM_WDTH_L-1:0]       I44993416e1d22613dbd78402c37a934d;
reg  [ 0:0]                      sgnprod_00048;
reg  [MAX_SUM_WDTH_L-1:0]        I03b70553f1c501609400574ae7cd73f5;
wire  [MAX_SUM_WDTH_L-1:0]       Ibc9b94a9dea471805cb442ac6904bc97;
wire  [MAX_SUM_WDTH_L-1:0]       I917d9f9b144d3bffafc77bddae7fba6b;
wire  [MAX_SUM_WDTH_L-1:0]       Ibc91c6c3d56bb8a14e22909c43ffec51;
wire  [MAX_SUM_WDTH_L-1:0]       If7c2d3eddd96b47b6c2aea8b27c8c7f4;
reg  [ 0:0]                      sgnprod_00049;
reg  [MAX_SUM_WDTH_L-1:0]        I63c9bf68b43ed66c51b0f4c0ed92e9ab;
wire  [MAX_SUM_WDTH_L-1:0]       I4df093ed94d26b058e97db550e347e3c;
wire  [MAX_SUM_WDTH_L-1:0]       Ie90303b0326bee4ab203a8cf1e643da9;
wire  [MAX_SUM_WDTH_L-1:0]       I19030d352fd059156ee42c66f9270beb;
wire  [MAX_SUM_WDTH_L-1:0]       I36767a902c53a384128ae1443cf88963;
reg  [ 0:0]                      sgnprod_00050;
reg  [MAX_SUM_WDTH_L-1:0]        If408dfead07757878cc878131bc7d6a3;
wire  [MAX_SUM_WDTH_L-1:0]       I868dffa3f07407f7996bb5bc596939b7;
wire  [MAX_SUM_WDTH_L-1:0]       I7d928be164d0dce8b1322ff230c053e9;
wire  [MAX_SUM_WDTH_L-1:0]       I98be4971a8a9a08abb3ebe474d7f0c6d;
wire  [MAX_SUM_WDTH_L-1:0]       I779e70dea33201e9237f29681ffd5e27;
reg  [ 0:0]                      sgnprod_00051;
reg  [MAX_SUM_WDTH_L-1:0]        Ia0857d63d309807789b6ff4f6028f1b3;
wire  [MAX_SUM_WDTH_L-1:0]       Ie2262914042172ab7e08599278f36af5;
wire  [MAX_SUM_WDTH_L-1:0]       I4001323da8f7956cdd480ac2d56df929;
wire  [MAX_SUM_WDTH_L-1:0]       Ib1cd6731034887a0a55e405c9db3e8de;
wire  [MAX_SUM_WDTH_L-1:0]       I51aa496e8c03944c28a908102514e6f8;
reg  [ 0:0]                      sgnprod_00052;
reg  [MAX_SUM_WDTH_L-1:0]        I53921b825c5e434b63bee0e1ecb7a517;
wire  [MAX_SUM_WDTH_L-1:0]       I6415f3996318472532e161510ccc8ca3;
wire  [MAX_SUM_WDTH_L-1:0]       Ia11b671b59240988737979328c472812;
wire  [MAX_SUM_WDTH_L-1:0]       Id4fabe0165a117a402dc14f2f3ec626a;
wire  [MAX_SUM_WDTH_L-1:0]       I57238f501ab7278b308d76211ced8cf7;
wire  [MAX_SUM_WDTH_L-1:0]       I9b257f8556ca4e5402637f01081b78e1;
reg  [ 0:0]                      sgnprod_00053;
reg  [MAX_SUM_WDTH_L-1:0]        I5e68f84e123c37f19a03c13892c77e19;
wire  [MAX_SUM_WDTH_L-1:0]       I2e093412a9fa3972cea01664389d8c27;
wire  [MAX_SUM_WDTH_L-1:0]       I17907fd8c6975c8c642535ff929221a6;
wire  [MAX_SUM_WDTH_L-1:0]       I3c6577b04ad56d864bbaa2c048323c11;
wire  [MAX_SUM_WDTH_L-1:0]       I6f0c341c05eaa8f35bbce4521f6e8f94;
wire  [MAX_SUM_WDTH_L-1:0]       Ib72ba950ecf9ae2668374f6633a67ca7;
reg  [ 0:0]                      sgnprod_00054;
reg  [MAX_SUM_WDTH_L-1:0]        Id5270b57c6fb4b18db3bbd0a523e467e;
wire  [MAX_SUM_WDTH_L-1:0]       I3d7c72d725f4563bb562e2992093cb02;
wire  [MAX_SUM_WDTH_L-1:0]       I813c881ac61a59041be3be78f6a466c8;
wire  [MAX_SUM_WDTH_L-1:0]       I866510e7dc721fa5aac312bc5ab5ba0a;
wire  [MAX_SUM_WDTH_L-1:0]       Ib4432359f97849dff6ad3e0f044157bd;
wire  [MAX_SUM_WDTH_L-1:0]       Ic86aa6eb1b4dcc2520309089b43292e6;
reg  [ 0:0]                      sgnprod_00055;
reg  [MAX_SUM_WDTH_L-1:0]        I3c18a84617eb21472d53e598700d7f4c;
wire  [MAX_SUM_WDTH_L-1:0]       I0731115afe5c15bcf131f7ef4f05802b;
wire  [MAX_SUM_WDTH_L-1:0]       Ib080b8fd34385aa7986dace4afd95267;
wire  [MAX_SUM_WDTH_L-1:0]       I134890b77451d0b78afc7402a6a28048;
wire  [MAX_SUM_WDTH_L-1:0]       I956da75f13433c1dd7a3cbd3b78922c1;
wire  [MAX_SUM_WDTH_L-1:0]       I440b26c9f1b9ccf70f97c9d5f732d38e;
reg  [ 0:0]                      sgnprod_00056;
reg  [MAX_SUM_WDTH_L-1:0]        Id36663e7a01fff3170833ecfecac1321;
wire  [MAX_SUM_WDTH_L-1:0]       I5e3a441faca44bffc4368d96d8fb0bfd;
wire  [MAX_SUM_WDTH_L-1:0]       I21d7ba25247a87a1a9c245d0d1f553b0;
wire  [MAX_SUM_WDTH_L-1:0]       I55aafa8162cfc4fccfae68cf78cd1c2b;
wire  [MAX_SUM_WDTH_L-1:0]       Ib99c25f0d8d6493cac4d5c816884c704;
wire  [MAX_SUM_WDTH_L-1:0]       Iee7c9f0a0e8ca127efee008b4874edbd;
reg  [ 0:0]                      sgnprod_00057;
reg  [MAX_SUM_WDTH_L-1:0]        I8d3be15109c7007a79fecaac0d891626;
wire  [MAX_SUM_WDTH_L-1:0]       I17b4a3baae65161387f472037ffc6fc4;
wire  [MAX_SUM_WDTH_L-1:0]       Ie7b7b202a968fe73f6b1e02a044414c5;
wire  [MAX_SUM_WDTH_L-1:0]       I479ab5c0e483c36267d8248340006666;
wire  [MAX_SUM_WDTH_L-1:0]       I777bfe165e25d7fde4fc950f23db7b84;
wire  [MAX_SUM_WDTH_L-1:0]       I146d505a34ddb8d65e0a1769f623a7fd;
reg  [ 0:0]                      sgnprod_00058;
reg  [MAX_SUM_WDTH_L-1:0]        I92169cc57291f20d336a479e392ec271;
wire  [MAX_SUM_WDTH_L-1:0]       Ia85239bddc04bf50bcf037ed2f76d7ac;
wire  [MAX_SUM_WDTH_L-1:0]       Ia7306bacf3c2b180d3261a5c1f0f4a30;
wire  [MAX_SUM_WDTH_L-1:0]       I2018147b86e47af5842c4f29d047d157;
wire  [MAX_SUM_WDTH_L-1:0]       Id17a85459845f8a8be694c4bf1fc29c9;
wire  [MAX_SUM_WDTH_L-1:0]       Ic012b15584d9d25af38f83d0526503da;
reg  [ 0:0]                      sgnprod_00059;
reg  [MAX_SUM_WDTH_L-1:0]        I6178b220b469b40dac39168057023a1c;
wire  [MAX_SUM_WDTH_L-1:0]       I7f09bd4a45143a036ce04af11b9927f9;
wire  [MAX_SUM_WDTH_L-1:0]       Ica32f94af6e6f3eaf2b724a2173fa463;
wire  [MAX_SUM_WDTH_L-1:0]       Ib750bb83ddfbbad2a2be8d1c8392b4ff;
wire  [MAX_SUM_WDTH_L-1:0]       I3906ece39480f96020717c6243e8ba4c;
wire  [MAX_SUM_WDTH_L-1:0]       Ie68ce21ade07fa53c30ebf27216b03f9;
reg  [ 0:0]                      sgnprod_00060;
reg  [MAX_SUM_WDTH_L-1:0]        I55342938216a0ea0889f96c2f6c05ce5;
wire  [MAX_SUM_WDTH_L-1:0]       I6cc6fa167c0d2b4b62ddbeecea175ed2;
wire  [MAX_SUM_WDTH_L-1:0]       Ibddf3468ae7c27d5a4b1388e524aa9c2;
wire  [MAX_SUM_WDTH_L-1:0]       Iadcb2b3acaac2e1bb505c65d3cbe4235;
wire  [MAX_SUM_WDTH_L-1:0]       I37cd96b8b0a4939d9a70098fd8bcf452;
reg  [ 0:0]                      sgnprod_00061;
reg  [MAX_SUM_WDTH_L-1:0]        Idf28431c76a84a48dd895979d2b11a63;
wire  [MAX_SUM_WDTH_L-1:0]       Ib34b169dcc76daee2d1aa2b2a7513af3;
wire  [MAX_SUM_WDTH_L-1:0]       If36fc316d6ec7c7e09eae77807b37099;
wire  [MAX_SUM_WDTH_L-1:0]       Ifd214c332218ac5c0fe5aded4b952711;
wire  [MAX_SUM_WDTH_L-1:0]       Idcd0fc8f86e2b6f03606b818b8346e5a;
reg  [ 0:0]                      sgnprod_00062;
reg  [MAX_SUM_WDTH_L-1:0]        I1ef61124c8d62e8f6a82a729fb091694;
wire  [MAX_SUM_WDTH_L-1:0]       If486aa8ac2cfb46f936714812cc760df;
wire  [MAX_SUM_WDTH_L-1:0]       I2d8e5b5fdbda7d599423c38aaace6658;
wire  [MAX_SUM_WDTH_L-1:0]       I6d0878fb7ec75c0a26be4dbba62f80dc;
wire  [MAX_SUM_WDTH_L-1:0]       I16a16ff0e8a6685a09803634da429fd2;
reg  [ 0:0]                      sgnprod_00063;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8bb96f0372323e6a8072ca56fb9396d;
wire  [MAX_SUM_WDTH_L-1:0]       Idb211abaa54ac26e7379c64a63f7d07c;
wire  [MAX_SUM_WDTH_L-1:0]       I351205eb71acb31b59d2b4470f0ba28c;
wire  [MAX_SUM_WDTH_L-1:0]       If5660c495bf7690252783d888d1ad6e8;
wire  [MAX_SUM_WDTH_L-1:0]       I3a5229cb8e44a15560b5c7bef96e65cc;
reg  [ 0:0]                      sgnprod_00064;
reg  [MAX_SUM_WDTH_L-1:0]        I432f74dda4f6b1cebdf5ad59c659080b;
wire  [MAX_SUM_WDTH_L-1:0]       I889b9b0828e97fe44d8366c5ef71a8f2;
wire  [MAX_SUM_WDTH_L-1:0]       Ie23062e00e39ead706f5b6ead233747d;
wire  [MAX_SUM_WDTH_L-1:0]       I8a2589544c75ecfdc31d28912c639695;
wire  [MAX_SUM_WDTH_L-1:0]       I5c21c59147e9c3a74c7cbbb6f2a23919;
wire  [MAX_SUM_WDTH_L-1:0]       Idacd78e24408e432abbbfb0c447fdde5;
reg  [ 0:0]                      sgnprod_00065;
reg  [MAX_SUM_WDTH_L-1:0]        Idc689442305acd00f0f32416d8fb3773;
wire  [MAX_SUM_WDTH_L-1:0]       I0e8b171fe5080485a7f4fef83f1f1528;
wire  [MAX_SUM_WDTH_L-1:0]       Ib22c2bd76e6c29cc2f1440885bf24b7b;
wire  [MAX_SUM_WDTH_L-1:0]       I149559fccd9def4ec1ead1fdcff3c7fd;
wire  [MAX_SUM_WDTH_L-1:0]       Icfa8fed3239748abca27a5fc17de79c0;
wire  [MAX_SUM_WDTH_L-1:0]       I2ff115fa483f080d93bada49a9566b33;
reg  [ 0:0]                      sgnprod_00066;
reg  [MAX_SUM_WDTH_L-1:0]        Ida03738adc101c03c2229756bed2469d;
wire  [MAX_SUM_WDTH_L-1:0]       Ibee4f3cd2f516c29ab68e07a640ab65e;
wire  [MAX_SUM_WDTH_L-1:0]       Ie495ab560f59ad038992c573de7d2f5b;
wire  [MAX_SUM_WDTH_L-1:0]       Ibd812def78c3a9c02f9ba45cc0413711;
wire  [MAX_SUM_WDTH_L-1:0]       I98166634dc80201b0cefb01d9559c228;
wire  [MAX_SUM_WDTH_L-1:0]       Ic2f03a980b5f0b042853ca746abab22b;
reg  [ 0:0]                      sgnprod_00067;
reg  [MAX_SUM_WDTH_L-1:0]        I4d14c75f28f3e516c259ea288996131b;
wire  [MAX_SUM_WDTH_L-1:0]       I2807a88097d2683ebdb9e0e785e3af02;
wire  [MAX_SUM_WDTH_L-1:0]       I8bebbb3a676c8506af0768516abcd740;
wire  [MAX_SUM_WDTH_L-1:0]       I31d380f34691c9fe9022035f233b77e2;
wire  [MAX_SUM_WDTH_L-1:0]       I1ffb5675c98ab5b3c62b24eb23441473;
wire  [MAX_SUM_WDTH_L-1:0]       If56424546ec4f3445853538207ea864e;
reg  [ 0:0]                      sgnprod_00068;
reg  [MAX_SUM_WDTH_L-1:0]        I6e6cbbf430d57f347a0d70558af143d8;
wire  [MAX_SUM_WDTH_L-1:0]       I31a49be4a34d9bac2e0d815097439772;
wire  [MAX_SUM_WDTH_L-1:0]       I6b96a2498078953e87de223aa2236d50;
wire  [MAX_SUM_WDTH_L-1:0]       I79bf36e298a85a42c7432f877055f0b4;
wire  [MAX_SUM_WDTH_L-1:0]       I90c070b9bde5da05e8a5d25d2de3ba6b;
wire  [MAX_SUM_WDTH_L-1:0]       I28d0e4e6d772dd58d845d91952ada300;
reg  [ 0:0]                      sgnprod_00069;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7487df45118e44acec6b9d07bbd5969;
wire  [MAX_SUM_WDTH_L-1:0]       I7232b4e277acc6f1acefcb606ca24508;
wire  [MAX_SUM_WDTH_L-1:0]       I32da124c433c55f692ffa4734d0dc8fc;
wire  [MAX_SUM_WDTH_L-1:0]       I56e487db14eeb8d93f494d2f11b57a49;
wire  [MAX_SUM_WDTH_L-1:0]       I94d3c02bd5b8e84926d4b3c2f56efeac;
wire  [MAX_SUM_WDTH_L-1:0]       I0c35b2e9176f9a06e26ca67d036411b4;
reg  [ 0:0]                      sgnprod_00070;
reg  [MAX_SUM_WDTH_L-1:0]        I492f382fea500462b3d0866240fb91b2;
wire  [MAX_SUM_WDTH_L-1:0]       Ia6ee7b70d0b7fe7c346760b1784e50b9;
wire  [MAX_SUM_WDTH_L-1:0]       I7ce57c278c683ad045526e49bcc47412;
wire  [MAX_SUM_WDTH_L-1:0]       Ie3d3e681cac0bb919946ac27057409e2;
wire  [MAX_SUM_WDTH_L-1:0]       I8ea0a8cdd6506c982ad75f23136bcebe;
wire  [MAX_SUM_WDTH_L-1:0]       Ic812f8bc775c5ee6a83e2b9aeb22b2a4;
reg  [ 0:0]                      sgnprod_00071;
reg  [MAX_SUM_WDTH_L-1:0]        I3fb3ebddaf28efb56092d19a1b4695de;
wire  [MAX_SUM_WDTH_L-1:0]       I0f0adf7fe957b9a68772bd8a1bc163d4;
wire  [MAX_SUM_WDTH_L-1:0]       If09562f8d82bc1dea7c38ed51523a889;
wire  [MAX_SUM_WDTH_L-1:0]       Ib0fd21d66cd89c4e5c95fbc9c7680b62;
wire  [MAX_SUM_WDTH_L-1:0]       I5a2b2bfadc638fe3fdc31136a8f09a8d;
wire  [MAX_SUM_WDTH_L-1:0]       Ica914d8c556285d6b90b35747065a6e5;
reg  [ 0:0]                      sgnprod_00072;
reg  [MAX_SUM_WDTH_L-1:0]        I22a26b7f0b1c8c16b00597732ce2ab23;
wire  [MAX_SUM_WDTH_L-1:0]       I00c5d739bccb0ab6d05da70fe51aafea;
wire  [MAX_SUM_WDTH_L-1:0]       I18e448761bc014ce490b766183350312;
wire  [MAX_SUM_WDTH_L-1:0]       I1b5920f488e9469bd416a6af3072a30b;
wire  [MAX_SUM_WDTH_L-1:0]       I70b41ffed4b6d88ddff219c567b8e968;
reg  [ 0:0]                      sgnprod_00073;
reg  [MAX_SUM_WDTH_L-1:0]        I2ac08a2d8c917ecb37fbaf5325cb0473;
wire  [MAX_SUM_WDTH_L-1:0]       I935e083b4561da7d015e98ca7f02854e;
wire  [MAX_SUM_WDTH_L-1:0]       Iaca9ef263bf220d786242b88c994fd21;
wire  [MAX_SUM_WDTH_L-1:0]       I92169291959eb33452b79bfd32618cbc;
wire  [MAX_SUM_WDTH_L-1:0]       I126dabc3ebb9c4157adf62b57f217bd0;
reg  [ 0:0]                      sgnprod_00074;
reg  [MAX_SUM_WDTH_L-1:0]        I50ff8f51e75fb9ce3db983c2a0f57196;
wire  [MAX_SUM_WDTH_L-1:0]       If4433b1ef2eb963cd301946958b69884;
wire  [MAX_SUM_WDTH_L-1:0]       I67ac5b9b794787b3c4738c3366689871;
wire  [MAX_SUM_WDTH_L-1:0]       I4f022d70078c412bdbef158f750d3da3;
wire  [MAX_SUM_WDTH_L-1:0]       I6be6165385f6a77aeedb88f2baaa9cab;
reg  [ 0:0]                      sgnprod_00075;
reg  [MAX_SUM_WDTH_L-1:0]        I444bc340ffb7ef7b72d4d2e761d58872;
wire  [MAX_SUM_WDTH_L-1:0]       Id1f7fe91547e158e1d39edffb1421ff3;
wire  [MAX_SUM_WDTH_L-1:0]       I7a51924134902612db53941390891245;
wire  [MAX_SUM_WDTH_L-1:0]       I45128b9e29dd2fdd94a78fc5ffdff2b1;
wire  [MAX_SUM_WDTH_L-1:0]       I7f1082408c8ebb5be18e8f71ff9510e5;
reg  [ 0:0]                      sgnprod_00076;
reg  [MAX_SUM_WDTH_L-1:0]        I039c6cac5830759529595a958b7f65c9;
wire  [MAX_SUM_WDTH_L-1:0]       I655ebf19c2f4b3dde716668f9ce12e59;
wire  [MAX_SUM_WDTH_L-1:0]       Ibc9d493a507122d92af42d858cdc4c61;
wire  [MAX_SUM_WDTH_L-1:0]       Ib3d3103e5ee4feb160a97c7e26f7102b;
wire  [MAX_SUM_WDTH_L-1:0]       I6cc56b119e72175df3b7ce64dc3d9305;
reg  [ 0:0]                      sgnprod_00077;
reg  [MAX_SUM_WDTH_L-1:0]        I0584de7d919236ab138e288a27d08ff1;
wire  [MAX_SUM_WDTH_L-1:0]       I57cf4a9378f1cdd94a1a5608dc57e05f;
wire  [MAX_SUM_WDTH_L-1:0]       I4160ab1aa18e8151c0a5c23b9edeb907;
wire  [MAX_SUM_WDTH_L-1:0]       Ia1f183f2d904d006e46399424e06c614;
wire  [MAX_SUM_WDTH_L-1:0]       If979702738671323995e56108bc9376c;
reg  [ 0:0]                      sgnprod_00078;
reg  [MAX_SUM_WDTH_L-1:0]        I086402c82ec67ae09a9e6360c58904b4;
wire  [MAX_SUM_WDTH_L-1:0]       Ibc96fe0a6bf1f95036f97c7d44fab575;
wire  [MAX_SUM_WDTH_L-1:0]       I755a38220a693ba43701d30e7e9508ad;
wire  [MAX_SUM_WDTH_L-1:0]       I896fb82baa9647a14f4b5b1ecfa70a15;
wire  [MAX_SUM_WDTH_L-1:0]       I23d1c973d7a2048353fbb68e4a294c08;
reg  [ 0:0]                      sgnprod_00079;
reg  [MAX_SUM_WDTH_L-1:0]        I1cefdc831c146187c77f861b3e2d1af0;
wire  [MAX_SUM_WDTH_L-1:0]       If9fd1e08af14f2fd4ca363383f48580a;
wire  [MAX_SUM_WDTH_L-1:0]       I8f3782f78d88a5c3bc93709564999b30;
wire  [MAX_SUM_WDTH_L-1:0]       I986d61d79ce31f4677f3293339db6ad2;
wire  [MAX_SUM_WDTH_L-1:0]       Ica4d93d9fad21316002008ade5106a9d;
reg  [ 0:0]                      sgnprod_00080;
reg  [MAX_SUM_WDTH_L-1:0]        Ida9c16ae57d17b6faee8a54838860447;
wire  [MAX_SUM_WDTH_L-1:0]       If77592d5d8bed32477fd690341e543d0;
wire  [MAX_SUM_WDTH_L-1:0]       I25b70c6b830cbfe1b41d8f289c751924;
wire  [MAX_SUM_WDTH_L-1:0]       I2a5d65eeffa18dd9af9fe36463dafd7c;
wire  [MAX_SUM_WDTH_L-1:0]       Ibafa6e10bd4edf5d224fdeb2f9adbf98;
reg  [ 0:0]                      sgnprod_00081;
reg  [MAX_SUM_WDTH_L-1:0]        Ia3b9fb112f39dd0ccbf7555659369efb;
wire  [MAX_SUM_WDTH_L-1:0]       Ifc25402bd879bc5c43b4945b60cd4540;
wire  [MAX_SUM_WDTH_L-1:0]       Iec48da6882325d8a33e0e0e845eb18a0;
wire  [MAX_SUM_WDTH_L-1:0]       I0fd05e46862fdf8e614afaa3fd478602;
wire  [MAX_SUM_WDTH_L-1:0]       I6253a59dca81842d9ab6e58cf204abbf;
reg  [ 0:0]                      sgnprod_00082;
reg  [MAX_SUM_WDTH_L-1:0]        Ib1bfcdc0c972aafc99116ed8c0511445;
wire  [MAX_SUM_WDTH_L-1:0]       Ib18d64bc58b354358ee6ac16785880e2;
wire  [MAX_SUM_WDTH_L-1:0]       I28689b693a7a5f761a1f252aa3ef3b67;
wire  [MAX_SUM_WDTH_L-1:0]       I1a4e6d12f9776d5e61094e0b5edf71d9;
wire  [MAX_SUM_WDTH_L-1:0]       I8e1ad23b7ac662bb827a83d3709f0adb;
reg  [ 0:0]                      sgnprod_00083;
reg  [MAX_SUM_WDTH_L-1:0]        I7adff505c50450a04f1717cac1adebe7;
wire  [MAX_SUM_WDTH_L-1:0]       I000ad2287813072cc18dad933758f2ab;
wire  [MAX_SUM_WDTH_L-1:0]       I7bc3698b51b89ac38ba5f4b5428a0c96;
wire  [MAX_SUM_WDTH_L-1:0]       I78aea1705621e2845a331c3e61a8055b;
wire  [MAX_SUM_WDTH_L-1:0]       I0a31314c3580f5f9e61e79c133e5d794;
reg  [ 0:0]                      sgnprod_00084;
reg  [MAX_SUM_WDTH_L-1:0]        I699feb4382974a02b21cb387c13f7f3f;
wire  [MAX_SUM_WDTH_L-1:0]       I0e274fd7bfc0388fef95a8ceb939ee91;
wire  [MAX_SUM_WDTH_L-1:0]       Id6f39ddcb73d3f4ec081a365d11d1ef4;
wire  [MAX_SUM_WDTH_L-1:0]       I807770bfa86d160459d6ec3c0f4d6a0b;
wire  [MAX_SUM_WDTH_L-1:0]       I31c89b8a11a3090bfd74b112cbc474bb;
reg  [ 0:0]                      sgnprod_00085;
reg  [MAX_SUM_WDTH_L-1:0]        Idc99c3b23e49aca3c98f0685ea34441c;
wire  [MAX_SUM_WDTH_L-1:0]       I79b82cb1bfc72bd5a9d313b9e9c9203c;
wire  [MAX_SUM_WDTH_L-1:0]       Ib1046ae03c9a77fd2c0b3e9838e9af87;
wire  [MAX_SUM_WDTH_L-1:0]       Ic63723fd43cbbbde51c233a3cca15d3f;
wire  [MAX_SUM_WDTH_L-1:0]       I3abbb59abada1aec6941185f95f738bd;
reg  [ 0:0]                      sgnprod_00086;
reg  [MAX_SUM_WDTH_L-1:0]        Ib67318fa6954ec8f3247927d34e74f8c;
wire  [MAX_SUM_WDTH_L-1:0]       I8d5bd7039a77ce82ce0f6cbba9c2a076;
wire  [MAX_SUM_WDTH_L-1:0]       I527ad0b9382dd7b6e657dc1a32d8e472;
wire  [MAX_SUM_WDTH_L-1:0]       I8de02f32e14e719f4930d99743c04a20;
wire  [MAX_SUM_WDTH_L-1:0]       I7614dd5e9628c761dd9b2a512cb1da98;
reg  [ 0:0]                      sgnprod_00087;
reg  [MAX_SUM_WDTH_L-1:0]        I8774ce3f11362915c4331d1026e452dd;
wire  [MAX_SUM_WDTH_L-1:0]       Icae7efa4742dd0ad943ee1f67b0c9b14;
wire  [MAX_SUM_WDTH_L-1:0]       Ieb1854b79e9a2bc6cf5aa1c319e8e753;
wire  [MAX_SUM_WDTH_L-1:0]       Iff50b77f300183ca59a67ccbcc9573c4;
wire  [MAX_SUM_WDTH_L-1:0]       I4868604f8178663de759d4c63dc6c4bd;
reg  [ 0:0]                      sgnprod_00088;
reg  [MAX_SUM_WDTH_L-1:0]        I2392b2d17ffed6073875fbe8e92534cf;
wire  [MAX_SUM_WDTH_L-1:0]       Ife992a151986c58df4cba79b6bc4ac0a;
wire  [MAX_SUM_WDTH_L-1:0]       I9ab973fb74d9fac5d78eb8fc2c7ecf36;
wire  [MAX_SUM_WDTH_L-1:0]       I5ee7916e859b86a98538659401685016;
reg  [ 0:0]                      sgnprod_00089;
reg  [MAX_SUM_WDTH_L-1:0]        I3a4f0d3e32596ef05477f494768d4266;
wire  [MAX_SUM_WDTH_L-1:0]       I48c284cefb8cfb5a938a8f23ce4d7f03;
wire  [MAX_SUM_WDTH_L-1:0]       I5c1fc666b77a689478654dd29519f458;
wire  [MAX_SUM_WDTH_L-1:0]       I38bba98b59184c75ba3b27e1dcf52182;
reg  [ 0:0]                      sgnprod_00090;
reg  [MAX_SUM_WDTH_L-1:0]        Icd08ff59cf6be3ba97698dd55703339e;
wire  [MAX_SUM_WDTH_L-1:0]       I6905b65403c16b0211643227ece536f6;
wire  [MAX_SUM_WDTH_L-1:0]       I3ed34401bba9d5f229bc98480aedd9a5;
wire  [MAX_SUM_WDTH_L-1:0]       Ib4d05804277cddc7f00ac17ac14f5325;
reg  [ 0:0]                      sgnprod_00091;
reg  [MAX_SUM_WDTH_L-1:0]        I985fb7ed22a8476ea322c9e3c2b3851c;
wire  [MAX_SUM_WDTH_L-1:0]       I41babdca6d3fa462849592d37b0a7998;
wire  [MAX_SUM_WDTH_L-1:0]       I58cfec706dc929ebfdeaca6e01b00c0a;
wire  [MAX_SUM_WDTH_L-1:0]       I7efe3c5b2fc69840a79545e0399ce749;
reg  [ 0:0]                      sgnprod_00092;
reg  [MAX_SUM_WDTH_L-1:0]        Ib985709316b1b0a9d3fa3c1eaf6c641f;
wire  [MAX_SUM_WDTH_L-1:0]       I70e3eeb2b3966676d16a6aa4c85753ab;
wire  [MAX_SUM_WDTH_L-1:0]       I2a32d545d1e7beecc7531174c7e8dfbc;
wire  [MAX_SUM_WDTH_L-1:0]       Ib8fb40e4ba0ba1f5e9f5a99d1271ed06;
wire  [MAX_SUM_WDTH_L-1:0]       Ica792cb9850a61fa4a8bd8a4b6c6ca05;
reg  [ 0:0]                      sgnprod_00093;
reg  [MAX_SUM_WDTH_L-1:0]        I4be898887dff6e2cebe53f135ece131b;
wire  [MAX_SUM_WDTH_L-1:0]       I779e5997c66649d6d54fd7f0514c47bd;
wire  [MAX_SUM_WDTH_L-1:0]       I5aa578b0c2831453683fa44af1878cb8;
wire  [MAX_SUM_WDTH_L-1:0]       I735d6229ef1a4ecda0a1f1dbdfb53fc1;
wire  [MAX_SUM_WDTH_L-1:0]       I62affd47512c5e8f0979244115624d97;
reg  [ 0:0]                      sgnprod_00094;
reg  [MAX_SUM_WDTH_L-1:0]        I004db04f61fb57aba81e15cc015442b3;
wire  [MAX_SUM_WDTH_L-1:0]       I14fe27afb3df5531b18dc9604e8dbe65;
wire  [MAX_SUM_WDTH_L-1:0]       Ib1b1626c84dad8ad13c058f921ffd57d;
wire  [MAX_SUM_WDTH_L-1:0]       Idf4a4bdddb88c21c5afe10a02373a6eb;
wire  [MAX_SUM_WDTH_L-1:0]       Iadefc2a3d07ed4b2c3c46b2ab5dec252;
reg  [ 0:0]                      sgnprod_00095;
reg  [MAX_SUM_WDTH_L-1:0]        I8f7e3dfb2f728d4cd1e79b82b62b0406;
wire  [MAX_SUM_WDTH_L-1:0]       I19315957077b037ffc6415dbb06ef789;
wire  [MAX_SUM_WDTH_L-1:0]       I1f9be09334407fc86c83a7c127e17bbe;
wire  [MAX_SUM_WDTH_L-1:0]       I28e17a5af7a7286a2643100d6d058dc0;
wire  [MAX_SUM_WDTH_L-1:0]       Icb2297c397bfe56be251ffb6b249a020;
reg  [ 0:0]                      sgnprod_00096;
reg  [MAX_SUM_WDTH_L-1:0]        I991054370345e61638ddaf81785505bd;
wire  [MAX_SUM_WDTH_L-1:0]       I64a48984527d660002f1f82c376c7a84;
wire  [MAX_SUM_WDTH_L-1:0]       I238b5fc70ce9f05b6322a2691b3a0207;
wire  [MAX_SUM_WDTH_L-1:0]       I00c16e7ad3821981032a42d5baa767b3;
wire  [MAX_SUM_WDTH_L-1:0]       I42fd5b094da200b33036e6cb8c7d0286;
reg  [ 0:0]                      sgnprod_00097;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa1f503965270d10e7a5c9a15576069b;
wire  [MAX_SUM_WDTH_L-1:0]       I98b7e26a0e9ec9ad750ff87cc0641a73;
wire  [MAX_SUM_WDTH_L-1:0]       I3ec904916870171bf837e162d1030052;
wire  [MAX_SUM_WDTH_L-1:0]       Iedb11b97900b7dd769d31f8a89521975;
wire  [MAX_SUM_WDTH_L-1:0]       Id0dceec6497c9f13ada07138986d4145;
reg  [ 0:0]                      sgnprod_00098;
reg  [MAX_SUM_WDTH_L-1:0]        I24f773842a4742fb58d09cae45717b2f;
wire  [MAX_SUM_WDTH_L-1:0]       Ibfe7d9bac29b8838f20cdcfe8ef7da0c;
wire  [MAX_SUM_WDTH_L-1:0]       I4d6c95605595942a34573d6ed55eb326;
wire  [MAX_SUM_WDTH_L-1:0]       Id6d8f32958dfa1a98958a84e7f1aed02;
wire  [MAX_SUM_WDTH_L-1:0]       I971cdf9ddd1bfff5664eec35f22da335;
reg  [ 0:0]                      sgnprod_00099;
reg  [MAX_SUM_WDTH_L-1:0]        I5bac7e0d778a547a0ae764fe259b6f7a;
wire  [MAX_SUM_WDTH_L-1:0]       Idd8bc1412a0dc5f489ef253a6164ceea;
wire  [MAX_SUM_WDTH_L-1:0]       Idbeec36de0128e5924e214877c82bf11;
wire  [MAX_SUM_WDTH_L-1:0]       I50a9cd240979bc56421bf85011ae99ed;
wire  [MAX_SUM_WDTH_L-1:0]       I6437095f6bad2d4fb2fbe0361f60bba1;
reg  [ 0:0]                      sgnprod_00100;
reg  [MAX_SUM_WDTH_L-1:0]        I255577ebee6768871df0224fc1db2db3;
wire  [MAX_SUM_WDTH_L-1:0]       Ie9b6eb3bbac26635aa00c38110958d46;
wire  [MAX_SUM_WDTH_L-1:0]       I9f34e81e3ffb85539a6273babc2a732e;
wire  [MAX_SUM_WDTH_L-1:0]       Id0a1ab8472d704001e0eba0317b117d6;
reg  [ 0:0]                      sgnprod_00101;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7fb4af3d3529a32f902a52cf5598474;
wire  [MAX_SUM_WDTH_L-1:0]       I9e632217cd0561d8faa28e4b8850d995;
wire  [MAX_SUM_WDTH_L-1:0]       Iedeb5b7b2fa8acf1ea083102678710ea;
wire  [MAX_SUM_WDTH_L-1:0]       I972431d1f5af0bdf4828e4f85591e358;
reg  [ 0:0]                      sgnprod_00102;
reg  [MAX_SUM_WDTH_L-1:0]        I2c98806141f064c9e92935b23a84ede1;
wire  [MAX_SUM_WDTH_L-1:0]       I1f41024b715d8312944ccbf70e95bb40;
wire  [MAX_SUM_WDTH_L-1:0]       Ia6bb5ca05f5d0af452c994dd50004e1d;
wire  [MAX_SUM_WDTH_L-1:0]       I9a1d1d1c862808f9a769cbdb3bc634e1;
reg  [ 0:0]                      sgnprod_00103;
reg  [MAX_SUM_WDTH_L-1:0]        I5680847bc8d224fa4ed93b2fc0d841e1;
wire  [MAX_SUM_WDTH_L-1:0]       I9734eb86f4e73ba217739baf5cb1b13c;
wire  [MAX_SUM_WDTH_L-1:0]       Ifc0fe00f86569956df72d8a960337e8c;
wire  [MAX_SUM_WDTH_L-1:0]       I223341a807a1d555f759632f67815159;
reg  [ 0:0]                      sgnprod_00104;
reg  [MAX_SUM_WDTH_L-1:0]        I365254279ebb10dd7ba0b3482d5e34cd;
wire  [MAX_SUM_WDTH_L-1:0]       I6c1f5cdf5f2917118941f4af14d67fef;
wire  [MAX_SUM_WDTH_L-1:0]       Ie84e88fd1aa2a0b90aa1715fcd27a329;
wire  [MAX_SUM_WDTH_L-1:0]       I558f70d7039a8bb58d8ea3f72e43dac0;
wire  [MAX_SUM_WDTH_L-1:0]       I9924269ed3de12f1f2a28893c7f95292;
wire  [MAX_SUM_WDTH_L-1:0]       If1153befd1396be2798cc14535ddeb8a;
reg  [ 0:0]                      sgnprod_00105;
reg  [MAX_SUM_WDTH_L-1:0]        I57bf4ad773cc058ae1bb7b1911dc3174;
wire  [MAX_SUM_WDTH_L-1:0]       I9bc447b20687fb3e7eff45792bd4dc3a;
wire  [MAX_SUM_WDTH_L-1:0]       If590520f01e452db9867a8d6d5dab29b;
wire  [MAX_SUM_WDTH_L-1:0]       Id93ee7d283016ab9b0aaa21237237c54;
wire  [MAX_SUM_WDTH_L-1:0]       Ic1cf03baabaed466fe532e4db3a9ea78;
wire  [MAX_SUM_WDTH_L-1:0]       If3031f9aa8f6eba90eac12db7839fefd;
reg  [ 0:0]                      sgnprod_00106;
reg  [MAX_SUM_WDTH_L-1:0]        I57072dfb29c4a3d2e2b40e46e62f0d95;
wire  [MAX_SUM_WDTH_L-1:0]       I0dc2708970ca2b6c092273b6626bacd6;
wire  [MAX_SUM_WDTH_L-1:0]       Ia58944aebf0b4f0a7d76a1444fced9de;
wire  [MAX_SUM_WDTH_L-1:0]       Iedd8e69679d10e05f2889f1d71cf0e7b;
wire  [MAX_SUM_WDTH_L-1:0]       I90f0d471914a2333b9dc14d6d01cf927;
wire  [MAX_SUM_WDTH_L-1:0]       Idceeb22013af64b6bb9f0d773e9ffe9a;
reg  [ 0:0]                      sgnprod_00107;
reg  [MAX_SUM_WDTH_L-1:0]        Id8cafb6f76321bdaba9711133be7be99;
wire  [MAX_SUM_WDTH_L-1:0]       If43574342e60a625fb6bee5a495e88f3;
wire  [MAX_SUM_WDTH_L-1:0]       Id285f055275014d9f23d35f91879afa1;
wire  [MAX_SUM_WDTH_L-1:0]       I8c803ab08db372802117de4fa4e2a187;
wire  [MAX_SUM_WDTH_L-1:0]       I13ba48a6b360f3cff5f37ce60cb735c6;
wire  [MAX_SUM_WDTH_L-1:0]       I4547cd1dad45dfd01e335e8cf20eadd6;
reg  [ 0:0]                      sgnprod_00108;
reg  [MAX_SUM_WDTH_L-1:0]        I6344e71ca2b0fd39d36caedd889c3085;
wire  [MAX_SUM_WDTH_L-1:0]       I0a305655b815b0cc159ac1c5f4ce30f8;
wire  [MAX_SUM_WDTH_L-1:0]       I3633737da6b74284b0ea9a06c3f5875f;
wire  [MAX_SUM_WDTH_L-1:0]       Ia949c1b338d1cba07cf6bb6572c3e322;
reg  [ 0:0]                      sgnprod_00109;
reg  [MAX_SUM_WDTH_L-1:0]        I0c99a68e0bed90afce18807acf7d55bb;
wire  [MAX_SUM_WDTH_L-1:0]       I9a0185f8400159415bc0ad6c38284041;
wire  [MAX_SUM_WDTH_L-1:0]       I3eeffe43e7deed7ee77a7f5a3bce3cd2;
wire  [MAX_SUM_WDTH_L-1:0]       I85af0c31ca7002ae569d9f5ce39943f7;
reg  [ 0:0]                      sgnprod_00110;
reg  [MAX_SUM_WDTH_L-1:0]        I1c95650979c86310ae2a949961c9db11;
wire  [MAX_SUM_WDTH_L-1:0]       I3dfb8d2fad83fbd807fbfc6330c5b857;
wire  [MAX_SUM_WDTH_L-1:0]       Ic12be21bcba5fa49437cc44dd8a7f064;
wire  [MAX_SUM_WDTH_L-1:0]       I713a384d022d3012e3d0019f5c4ac077;
reg  [ 0:0]                      sgnprod_00111;
reg  [MAX_SUM_WDTH_L-1:0]        I04eaefa5d133e53494fc270b07be7043;
wire  [MAX_SUM_WDTH_L-1:0]       I80550019479d0323d0dd7e7d0f767d83;
wire  [MAX_SUM_WDTH_L-1:0]       Ib8a866f080dd997e0b6c93b6c844d1bc;
wire  [MAX_SUM_WDTH_L-1:0]       Id542de206d736ee3769ea0bd037cb627;
reg  [ 0:0]                      sgnprod_00112;
reg  [MAX_SUM_WDTH_L-1:0]        I4a64fa2412eb8058c2dfd9351d7b297d;
wire  [MAX_SUM_WDTH_L-1:0]       I77e6cdb09c92492c3303d0213de9c291;
wire  [MAX_SUM_WDTH_L-1:0]       I788c33a9f94b26f4ce0f515891d06f90;
wire  [MAX_SUM_WDTH_L-1:0]       Iaf7074c2b570a296fe2ea8a5a7097ca0;
wire  [MAX_SUM_WDTH_L-1:0]       I8964c6d3f8e02866a6ad86553ab05d99;
reg  [ 0:0]                      sgnprod_00113;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8bb2fcb752c6a33254963d1ebb4130d;
wire  [MAX_SUM_WDTH_L-1:0]       I2aa25edaca90c9dae8ed63b48d333c17;
wire  [MAX_SUM_WDTH_L-1:0]       I51a440917c7ae23339bec6f8a745c103;
wire  [MAX_SUM_WDTH_L-1:0]       I56ce875e4619d4d8d6ca2fa0ddee91b1;
wire  [MAX_SUM_WDTH_L-1:0]       I80607da8f92f5a5d2e4798a62a7b1c5c;
reg  [ 0:0]                      sgnprod_00114;
reg  [MAX_SUM_WDTH_L-1:0]        Iac05b7e3ae18f948b72c356ccfb8000f;
wire  [MAX_SUM_WDTH_L-1:0]       Ic4dcaa520e26bac40b3876f02074f856;
wire  [MAX_SUM_WDTH_L-1:0]       I3b2714d34081a3b6cccc47fa1638e72e;
wire  [MAX_SUM_WDTH_L-1:0]       I2db1d1ee8f546c00e512875ce2e13cee;
wire  [MAX_SUM_WDTH_L-1:0]       If80a6bb104ff3b2020e909103c104063;
reg  [ 0:0]                      sgnprod_00115;
reg  [MAX_SUM_WDTH_L-1:0]        I27da3f75cca6c49e55db90306aa68e94;
wire  [MAX_SUM_WDTH_L-1:0]       Iadb72cc5444816fbd132256493930bb4;
wire  [MAX_SUM_WDTH_L-1:0]       I3a8ec1ad07bfada3d2c6ffca88b8b678;
wire  [MAX_SUM_WDTH_L-1:0]       I0aa042b86d9f68d22a49b4eb480a9088;
wire  [MAX_SUM_WDTH_L-1:0]       I89a387374771b68d87d7ff2dcc810829;
reg  [ 0:0]                      sgnprod_00116;
reg  [MAX_SUM_WDTH_L-1:0]        Idc7fed723190098341225fe01ba65ced;
wire  [MAX_SUM_WDTH_L-1:0]       I2935b3d5c3bba4dddfc7ae03fa77b229;
wire  [MAX_SUM_WDTH_L-1:0]       I4e0c0248f4aa97d263d64dfec36e3aa2;
wire  [MAX_SUM_WDTH_L-1:0]       Ia2871d7493b2727d2cb2fbab596b7e6a;
reg  [ 0:0]                      sgnprod_00117;
reg  [MAX_SUM_WDTH_L-1:0]        Ife9065805598960919ee4f14c3cc6fd4;
wire  [MAX_SUM_WDTH_L-1:0]       Ie57adae8873946d6c706074b52a49786;
wire  [MAX_SUM_WDTH_L-1:0]       If5ac85646e4b339a19af658f01d0a17f;
wire  [MAX_SUM_WDTH_L-1:0]       I1c092426f34be030b3e020f40517b0e1;
reg  [ 0:0]                      sgnprod_00118;
reg  [MAX_SUM_WDTH_L-1:0]        I717c5c2d6a2be61593492ae5f17a112f;
wire  [MAX_SUM_WDTH_L-1:0]       Ic719b72ad271bc7c077067518e6bbb98;
wire  [MAX_SUM_WDTH_L-1:0]       Ib87362230682c88d68a0ba70e25f3c20;
wire  [MAX_SUM_WDTH_L-1:0]       Ifcf097a102f8dc1f912022fed893d222;
reg  [ 0:0]                      sgnprod_00119;
reg  [MAX_SUM_WDTH_L-1:0]        I4c31fa8e6eb648439cdae1de1afe0d6f;
wire  [MAX_SUM_WDTH_L-1:0]       I56483ca3fa550dc59bfa347780cfef7b;
wire  [MAX_SUM_WDTH_L-1:0]       I4aa9f61be376458185c3235442c8fda0;
wire  [MAX_SUM_WDTH_L-1:0]       Id91fde1007d47258273299de80721390;
reg  [ 0:0]                      sgnprod_00120;
reg  [MAX_SUM_WDTH_L-1:0]        Iead549a9af27f1fced7d9c36e7b5c3f5;
wire  [MAX_SUM_WDTH_L-1:0]       Id58498c34aff2e1216c189b9df88822c;
wire  [MAX_SUM_WDTH_L-1:0]       Ib52e0c68caadcf4dd9636a84f5460e53;
wire  [MAX_SUM_WDTH_L-1:0]       Ie19679053b289bb5a0aad570cc81bd14;
wire  [MAX_SUM_WDTH_L-1:0]       I8862c5ef45b723c9abf5d0ab6854a900;
wire  [MAX_SUM_WDTH_L-1:0]       I30db951a07af96a8ddf59360141b9a6a;
reg  [ 0:0]                      sgnprod_00121;
reg  [MAX_SUM_WDTH_L-1:0]        I10422eb79364e7d0e21e1643d9060331;
wire  [MAX_SUM_WDTH_L-1:0]       I4855a0a0c6426d33014ce6a4c96965ce;
wire  [MAX_SUM_WDTH_L-1:0]       I362e8db1791718290bd33a79b4fc0855;
wire  [MAX_SUM_WDTH_L-1:0]       I773f0508440fb71d73fd82a372cc0a00;
wire  [MAX_SUM_WDTH_L-1:0]       I792891cecae468d7a87e12f2da62a718;
wire  [MAX_SUM_WDTH_L-1:0]       I33303820ad094d7a0ab53bca722fc609;
reg  [ 0:0]                      sgnprod_00122;
reg  [MAX_SUM_WDTH_L-1:0]        I914cb87eba8baa40cd515334e59f26b2;
wire  [MAX_SUM_WDTH_L-1:0]       Iff98739de575e25104c0dc30f08912a5;
wire  [MAX_SUM_WDTH_L-1:0]       I1952614b64ea451e9d0646dcce5dd1cd;
wire  [MAX_SUM_WDTH_L-1:0]       I49c1a7d1c20a25496821ad80c7eff790;
wire  [MAX_SUM_WDTH_L-1:0]       Ie2be17a55e79ca76350e033f227800de;
wire  [MAX_SUM_WDTH_L-1:0]       I737a5b06f848cacf0c8da4985c73c66b;
reg  [ 0:0]                      sgnprod_00123;
reg  [MAX_SUM_WDTH_L-1:0]        I32ed679af4ab759901aee43c9d93eb67;
wire  [MAX_SUM_WDTH_L-1:0]       Iab160609bb21501aa55b662d2010357b;
wire  [MAX_SUM_WDTH_L-1:0]       Ief74f1a9d4a43ee5c9def7b83369bb21;
wire  [MAX_SUM_WDTH_L-1:0]       Id144423f50751e661db3860a8487d004;
wire  [MAX_SUM_WDTH_L-1:0]       I623352a4f6705b21d461d6b32e85c12b;
wire  [MAX_SUM_WDTH_L-1:0]       I28d1dc8dc594977b5058b5bb9f6bfc66;
reg  [ 0:0]                      sgnprod_00124;
reg  [MAX_SUM_WDTH_L-1:0]        Id376dfa5141402f4d41a8858180ed87e;
wire  [MAX_SUM_WDTH_L-1:0]       I5371a83bf9d6f334cf8d1c5b082527e9;
wire  [MAX_SUM_WDTH_L-1:0]       If1605d6646fd267e701668a7245b3b44;
wire  [MAX_SUM_WDTH_L-1:0]       Idf5eb1ac2c5bd92fa08ed935ae298255;
reg  [ 0:0]                      sgnprod_00125;
reg  [MAX_SUM_WDTH_L-1:0]        I98a384bc62ee03f5ad7df20ef2d9af95;
wire  [MAX_SUM_WDTH_L-1:0]       I44ce30330c4d2d6033a0a970dd2bdd68;
wire  [MAX_SUM_WDTH_L-1:0]       Ic101b8f56ea1e25c6b752583a1b01242;
wire  [MAX_SUM_WDTH_L-1:0]       Ib7cf44e681881e55d2d353280a6319d6;
reg  [ 0:0]                      sgnprod_00126;
reg  [MAX_SUM_WDTH_L-1:0]        Icfed259ca2bb2732d8e0c26ef67cd4cf;
wire  [MAX_SUM_WDTH_L-1:0]       I35690f724e964248dbb1e80fb1ea49f8;
wire  [MAX_SUM_WDTH_L-1:0]       I5affa2759148a6baf5b9f0cd3122348c;
wire  [MAX_SUM_WDTH_L-1:0]       Iaeea1f06ff0c6e9cfa43ba14420c3adc;
reg  [ 0:0]                      sgnprod_00127;
reg  [MAX_SUM_WDTH_L-1:0]        I20861535c450d6e6bf11c45dac120454;
wire  [MAX_SUM_WDTH_L-1:0]       Iac5a23266c3b038b4b54a916dccdf3a8;
wire  [MAX_SUM_WDTH_L-1:0]       Icdfb7f52cc27b1cfcde90a100d29af13;
wire  [MAX_SUM_WDTH_L-1:0]       I71484d7e00efa02a08b54a1405f2902c;
reg  [ 0:0]                      sgnprod_00128;
reg  [MAX_SUM_WDTH_L-1:0]        I013929385ad819ddfcfcc59c22902ee3;
wire  [MAX_SUM_WDTH_L-1:0]       I68a9b0607e69e8b3dae64689eb288a33;
wire  [MAX_SUM_WDTH_L-1:0]       I2598c48aad48072a7f216b2ab56ee532;
wire  [MAX_SUM_WDTH_L-1:0]       I796e3a193b1b66fa9a04ca60aee11ea1;
wire  [MAX_SUM_WDTH_L-1:0]       Ic96be7e69faf0f43b92618131cf0c98a;
reg  [ 0:0]                      sgnprod_00129;
reg  [MAX_SUM_WDTH_L-1:0]        I34fffcb07fe82f11fe142f7c37f39155;
wire  [MAX_SUM_WDTH_L-1:0]       I648afe4114ce435bf1d13e0ad54425cf;
wire  [MAX_SUM_WDTH_L-1:0]       If05d7e30b4717e0a1bfd20b90d0539bd;
wire  [MAX_SUM_WDTH_L-1:0]       I5fc356af8a62a1d739cb375fb851e90f;
wire  [MAX_SUM_WDTH_L-1:0]       I22f4c5403fbe33d18f97cf21786cdd80;
reg  [ 0:0]                      sgnprod_00130;
reg  [MAX_SUM_WDTH_L-1:0]        I61ca60fde05ed88cce714dcd8c13b827;
wire  [MAX_SUM_WDTH_L-1:0]       I9a1b2b9f924099f1e57fa501ba2e33ba;
wire  [MAX_SUM_WDTH_L-1:0]       If6253af4ebc430e4937269a5f4989b29;
wire  [MAX_SUM_WDTH_L-1:0]       I0427d17423548dbb33cf792883b4be8c;
wire  [MAX_SUM_WDTH_L-1:0]       Ie539faf01ae85253e399308fef98afd6;
reg  [ 0:0]                      sgnprod_00131;
reg  [MAX_SUM_WDTH_L-1:0]        I4907dd45c158dc7e0041c64f1fb388f6;
wire  [MAX_SUM_WDTH_L-1:0]       Iae6e7c42f250cd9223f18f8830fb177d;
wire  [MAX_SUM_WDTH_L-1:0]       Iff47ec1743b59d7f90e9042af7ce44cb;
wire  [MAX_SUM_WDTH_L-1:0]       I1cf4a55ebab332defa32d2922b885285;
wire  [MAX_SUM_WDTH_L-1:0]       I284913858691ad5724073b73a820047a;
reg  [ 0:0]                      sgnprod_00132;
reg  [MAX_SUM_WDTH_L-1:0]        I2c8f6a9b9f655b317bb0af4d60fdbc4b;
wire  [MAX_SUM_WDTH_L-1:0]       I35626ca53adbbf0a3a71cc6fcf43bcb1;
wire  [MAX_SUM_WDTH_L-1:0]       I0d74ef22d31abcec73c7c582310b1e6d;
wire  [MAX_SUM_WDTH_L-1:0]       I15f4cf1aa0ad5ce2bda52df338e677e3;
wire  [MAX_SUM_WDTH_L-1:0]       I6c5ca5e68c8844bb1617a2288b5bbc37;
reg  [ 0:0]                      sgnprod_00133;
reg  [MAX_SUM_WDTH_L-1:0]        Ic7dff631559304ec59f0696c66436d62;
wire  [MAX_SUM_WDTH_L-1:0]       I44343a9491069c3c8ea4fbd6255a5a6c;
wire  [MAX_SUM_WDTH_L-1:0]       I1d8318b94d86e1fd28323a5e5684a37b;
wire  [MAX_SUM_WDTH_L-1:0]       I825e83bd88575868f4fcc9a8b8729663;
wire  [MAX_SUM_WDTH_L-1:0]       I3184a16c71cff80c8c90b40e45f114b8;
reg  [ 0:0]                      sgnprod_00134;
reg  [MAX_SUM_WDTH_L-1:0]        I6a239d3e55b4a9a3be9989a85bbec545;
wire  [MAX_SUM_WDTH_L-1:0]       Iae133550f8bad8357a73e7de1372faa3;
wire  [MAX_SUM_WDTH_L-1:0]       Ibccb4a43c410f698e0fff68553326a77;
wire  [MAX_SUM_WDTH_L-1:0]       I72dc7aa294a3af89101ea62a4223170e;
wire  [MAX_SUM_WDTH_L-1:0]       I91eb3e70921e0b141a344bc57dfbc934;
reg  [ 0:0]                      sgnprod_00135;
reg  [MAX_SUM_WDTH_L-1:0]        I630f905e55f08e7d1569a08e937ad216;
wire  [MAX_SUM_WDTH_L-1:0]       I1986f22f2269cc135c6ed28d35fb0bd1;
wire  [MAX_SUM_WDTH_L-1:0]       Ibef24017bc71de9c002aafa7ce9a784c;
wire  [MAX_SUM_WDTH_L-1:0]       Ieae3ed78fa2c45507066f4e20d96e956;
wire  [MAX_SUM_WDTH_L-1:0]       I730fd25ffc7778fd4bb02d33cb3870d6;
reg  [ 0:0]                      sgnprod_00136;
reg  [MAX_SUM_WDTH_L-1:0]        I8d13eb3669785c4279c685763d4f3fad;
wire  [MAX_SUM_WDTH_L-1:0]       I9a32313f2911b797fb0848f7d97e62b9;
wire  [MAX_SUM_WDTH_L-1:0]       I6373e2d64fdb5dd77733b3e4bb405121;
wire  [MAX_SUM_WDTH_L-1:0]       Ib437aa67ab7c13b45d7a4d56ce9e79b8;
wire  [MAX_SUM_WDTH_L-1:0]       I0cb5c7a759f4c75d4a675f9777f15c5f;
reg  [ 0:0]                      sgnprod_00137;
reg  [MAX_SUM_WDTH_L-1:0]        I25a6f3de9a9a01cbbdd32ed848561aa4;
wire  [MAX_SUM_WDTH_L-1:0]       I0ca91c1426ba14a7b47a081cb3becd19;
wire  [MAX_SUM_WDTH_L-1:0]       I0737e0cc7453e328efab2277bb712ea8;
wire  [MAX_SUM_WDTH_L-1:0]       I456af863661122cc303fccb235f3c7a1;
wire  [MAX_SUM_WDTH_L-1:0]       Idc5916c4800e9f647d51c52444ab6fff;
reg  [ 0:0]                      sgnprod_00138;
reg  [MAX_SUM_WDTH_L-1:0]        Iba3dd4b2c2c85c4cfe770d9b52ef4634;
wire  [MAX_SUM_WDTH_L-1:0]       I57aca70e2b8d126c120736b2606ed333;
wire  [MAX_SUM_WDTH_L-1:0]       Ic6650a6d092b749b4498c08d69cf815e;
wire  [MAX_SUM_WDTH_L-1:0]       Ic2e3b8f91eb218650c7b9c515c7efe97;
wire  [MAX_SUM_WDTH_L-1:0]       I93a084aa1e6881ab8dc905dcdcdfd7ee;
reg  [ 0:0]                      sgnprod_00139;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1b744387b5200a504e4874e14d2f282;
wire  [MAX_SUM_WDTH_L-1:0]       I8cba172573be52c5a90bd40e6f40a508;
wire  [MAX_SUM_WDTH_L-1:0]       I1cccfd1516af59265731121dde878116;
wire  [MAX_SUM_WDTH_L-1:0]       Ia171bbefe2d20b4c058126c33ef28eb8;
wire  [MAX_SUM_WDTH_L-1:0]       I84bc44a5d53a8f66b985b70c7ec1ae7c;
reg  [ 0:0]                      sgnprod_00140;
reg  [MAX_SUM_WDTH_L-1:0]        Icf76cb69aedf4db01cd3444f4c4ba471;
wire  [MAX_SUM_WDTH_L-1:0]       I321b104ca3c818018d4b03adfe1110b9;
wire  [MAX_SUM_WDTH_L-1:0]       Ia79b8994da536c86634bf6f54a21145d;
wire  [MAX_SUM_WDTH_L-1:0]       I4df55ce80eec5fee295b5a0ae92bd6c8;
wire  [MAX_SUM_WDTH_L-1:0]       I46593a7956590d870fe680228081a6d2;
reg  [ 0:0]                      sgnprod_00141;
reg  [MAX_SUM_WDTH_L-1:0]        I4857b5b50556c8e7fff4b2d3e08e4b28;
wire  [MAX_SUM_WDTH_L-1:0]       I906e9da31de73ae45579607a014e8b54;
wire  [MAX_SUM_WDTH_L-1:0]       If5dd1a1b9e3fc0e67a85da3183480aed;
wire  [MAX_SUM_WDTH_L-1:0]       Iadfb1571c78c3f0c05e4ef498267df24;
wire  [MAX_SUM_WDTH_L-1:0]       Icebb43b184c2745cc9da9d01b06bc62f;
reg  [ 0:0]                      sgnprod_00142;
reg  [MAX_SUM_WDTH_L-1:0]        I0a1e9cf99f1d4725327615f50fcc3ad0;
wire  [MAX_SUM_WDTH_L-1:0]       I6e4b0489ec7333abf2245a1b72a8923d;
wire  [MAX_SUM_WDTH_L-1:0]       I24ac5dd30526c1d3bc7b941103a66804;
wire  [MAX_SUM_WDTH_L-1:0]       I33681b2292c086fe536dae2aec70903a;
wire  [MAX_SUM_WDTH_L-1:0]       Ia373ca76c3b15a4148532b3822f82ba5;
reg  [ 0:0]                      sgnprod_00143;
reg  [MAX_SUM_WDTH_L-1:0]        Ie844f4c446983ce381b0bc4c0e8ef7d7;
wire  [MAX_SUM_WDTH_L-1:0]       I7d08adbaf66cea04be4891db610bca3f;
wire  [MAX_SUM_WDTH_L-1:0]       Ic09ed51b20f411683a801eaad61657a3;
wire  [MAX_SUM_WDTH_L-1:0]       I6a9af8c9009b5de47ebe9ee8b79d3831;
wire  [MAX_SUM_WDTH_L-1:0]       Ife18e8a16d4437161b75a93e3dff1b5b;
reg  [ 0:0]                      sgnprod_00144;
reg  [MAX_SUM_WDTH_L-1:0]        I6067f47cccceea96ac46ff0d457b25f2;
wire  [MAX_SUM_WDTH_L-1:0]       I0cde86532c8db1a32d9fbe38a40b91b8;
wire  [MAX_SUM_WDTH_L-1:0]       I49c8ec4cd33e6caed8ed7dab779e7ebb;
wire  [MAX_SUM_WDTH_L-1:0]       Idb86f95570587a0711d796aac7004c25;
wire  [MAX_SUM_WDTH_L-1:0]       I2d1373d0b18992fa46a9607a86d21520;
reg  [ 0:0]                      sgnprod_00145;
reg  [MAX_SUM_WDTH_L-1:0]        Ifd6fd1f3cbf8884ca7f64bc42278e4fa;
wire  [MAX_SUM_WDTH_L-1:0]       I30f26e090ab14551cbac41883ad8a152;
wire  [MAX_SUM_WDTH_L-1:0]       Ib1b4e41ab25733d1d6dd54e1fe81a419;
wire  [MAX_SUM_WDTH_L-1:0]       I146c0d5154a6de44c0536de873904ccf;
wire  [MAX_SUM_WDTH_L-1:0]       I8eb9d4839a478a4e28b45a549b5682a4;
reg  [ 0:0]                      sgnprod_00146;
reg  [MAX_SUM_WDTH_L-1:0]        Iaec9fd9e79371676bfa8ff14b4feae52;
wire  [MAX_SUM_WDTH_L-1:0]       I2501ef991a59512c43693ba9d7db8571;
wire  [MAX_SUM_WDTH_L-1:0]       I38213f78fd4dc52f9d2c9b7b22136c1c;
wire  [MAX_SUM_WDTH_L-1:0]       I49ce91ac152279af421bbc6c4d9b8087;
wire  [MAX_SUM_WDTH_L-1:0]       I6a2b7bb2cb3ca2ab932c211a68dded55;
reg  [ 0:0]                      sgnprod_00147;
reg  [MAX_SUM_WDTH_L-1:0]        I500757c4eda5d3d899aee47b87da585b;
wire  [MAX_SUM_WDTH_L-1:0]       Idaae6ba9da8754615a2c34ef859492db;
wire  [MAX_SUM_WDTH_L-1:0]       Icaca9fc70a3ec6c48c0e41f8168e2bb9;
wire  [MAX_SUM_WDTH_L-1:0]       I4f69b8ff834c7ab3194bc9390ce0f5f6;
wire  [MAX_SUM_WDTH_L-1:0]       I037cb596cd48c5533ed22bc32518d992;
reg  [ 0:0]                      sgnprod_00148;
reg  [MAX_SUM_WDTH_L-1:0]        I47bf091b0fa74ad511a760bad9d2506c;
wire  [MAX_SUM_WDTH_L-1:0]       I94a89577951de90edc4f73b281ad7364;
wire  [MAX_SUM_WDTH_L-1:0]       Ib7493a1a384aebaa7999ff1fb867fc6b;
wire  [MAX_SUM_WDTH_L-1:0]       I2ceb9e423696539135c5bae5cc2d8d98;
reg  [ 0:0]                      sgnprod_00149;
reg  [MAX_SUM_WDTH_L-1:0]        Ia4c3d0cd9957f678880de5775de76e0d;
wire  [MAX_SUM_WDTH_L-1:0]       Ia6bbf236436b2ed22bbaae3b8849de6d;
wire  [MAX_SUM_WDTH_L-1:0]       I33cdaee4676d546dd5507df4704ea1f8;
wire  [MAX_SUM_WDTH_L-1:0]       Ia44daa9ddc3e4d377267333813d4675f;
reg  [ 0:0]                      sgnprod_00150;
reg  [MAX_SUM_WDTH_L-1:0]        If5f957fa2f055b1c2c28e8d7cfe3e9ad;
wire  [MAX_SUM_WDTH_L-1:0]       Ie1f8fff3f43426d6bc39e45322a532ca;
wire  [MAX_SUM_WDTH_L-1:0]       I4ee181895efc22862b6e85802a944095;
wire  [MAX_SUM_WDTH_L-1:0]       I5c24ea83cabbb6be089ac084732cb9d6;
reg  [ 0:0]                      sgnprod_00151;
reg  [MAX_SUM_WDTH_L-1:0]        I3608378a5da8c66bef58528d56192530;
wire  [MAX_SUM_WDTH_L-1:0]       Ifee2342449a3b3d0036ce2ecbc9ae189;
wire  [MAX_SUM_WDTH_L-1:0]       I70a9a9b8f25066612a50e411ad68e6c4;
wire  [MAX_SUM_WDTH_L-1:0]       I1870059af857c79d444bef948bb536ef;
reg  [ 0:0]                      sgnprod_00152;
reg  [MAX_SUM_WDTH_L-1:0]        Ie6dead855e00ea0a8e6a9b7503aaebb8;
wire  [MAX_SUM_WDTH_L-1:0]       Iafe61ab12e232a1090123a0f16eefaca;
wire  [MAX_SUM_WDTH_L-1:0]       I10ca809fe9a04eaf5d7784ba69314178;
wire  [MAX_SUM_WDTH_L-1:0]       I7a1bd0a115b3a1f85cb9c54840f5bf9b;
wire  [MAX_SUM_WDTH_L-1:0]       I986a564393d944d7d202414431c6d165;
reg  [ 0:0]                      sgnprod_00153;
reg  [MAX_SUM_WDTH_L-1:0]        I3bae5e6862e003a8b9a476f72cc6858b;
wire  [MAX_SUM_WDTH_L-1:0]       I464042aaa60a41c7e1faf3d16eeb121d;
wire  [MAX_SUM_WDTH_L-1:0]       I34b9a0bf2b6b562fb36291022ddf5179;
wire  [MAX_SUM_WDTH_L-1:0]       I17dd8612b5c7f9dcc90f17e584aab2d3;
wire  [MAX_SUM_WDTH_L-1:0]       Id77cf7c05844d83e808a694971145261;
reg  [ 0:0]                      sgnprod_00154;
reg  [MAX_SUM_WDTH_L-1:0]        I4431adecba8be9e5f21bc6b3e1f8cb10;
wire  [MAX_SUM_WDTH_L-1:0]       I276c1155d766437253f12b25066b84e4;
wire  [MAX_SUM_WDTH_L-1:0]       Id75b386d8076893cb73baca69c3eff59;
wire  [MAX_SUM_WDTH_L-1:0]       If62ddbe87274965cfd83189c6666401e;
wire  [MAX_SUM_WDTH_L-1:0]       I4f73a07452638a610b31e3ee52cb5639;
reg  [ 0:0]                      sgnprod_00155;
reg  [MAX_SUM_WDTH_L-1:0]        I21c7a2885126d532d00484376588a469;
wire  [MAX_SUM_WDTH_L-1:0]       I2a4faf3344d9bf4ee71da0be8994788a;
wire  [MAX_SUM_WDTH_L-1:0]       I7d7ad0cbb962a47e229fe9d8406e6fe1;
wire  [MAX_SUM_WDTH_L-1:0]       I82988dc2dc83ac61380d2a5cb6551768;
wire  [MAX_SUM_WDTH_L-1:0]       I058c3a9848fd30010e4742d8682081ac;
reg  [ 0:0]                      sgnprod_00156;
reg  [MAX_SUM_WDTH_L-1:0]        I2c4d7339ff2fe68d060dd8d961dcab8c;
wire  [MAX_SUM_WDTH_L-1:0]       I368121c2534820a7147858c06e58b3fc;
wire  [MAX_SUM_WDTH_L-1:0]       I03d4541eeb1440aa72ee490c49977e32;
wire  [MAX_SUM_WDTH_L-1:0]       I75fdf5a355949a87b768b1e67db674e4;
wire  [MAX_SUM_WDTH_L-1:0]       I088f4a0af0239602d422324549cb9799;
reg  [ 0:0]                      sgnprod_00157;
reg  [MAX_SUM_WDTH_L-1:0]        Iee518b15b067eec58cccfa37f7432ea5;
wire  [MAX_SUM_WDTH_L-1:0]       I787fe66b38237caf805ec14970d154c7;
wire  [MAX_SUM_WDTH_L-1:0]       Icef176cff3ae503dbbe2af9ecfc4c859;
wire  [MAX_SUM_WDTH_L-1:0]       Ie0a66e4871bfe94f6716279ecc9ef21c;
wire  [MAX_SUM_WDTH_L-1:0]       I474adf7a975b405c288058139a08be38;
reg  [ 0:0]                      sgnprod_00158;
reg  [MAX_SUM_WDTH_L-1:0]        I42145be9c2a80288ba4a2edd91f661a3;
wire  [MAX_SUM_WDTH_L-1:0]       Iebeadb39658f41dcf8719ed413e46144;
wire  [MAX_SUM_WDTH_L-1:0]       Ie018b0d9f05a86207ae09ca2efac54e2;
wire  [MAX_SUM_WDTH_L-1:0]       I51ee69807609fca0f332c8bc31afd632;
wire  [MAX_SUM_WDTH_L-1:0]       Iee1cb471704b2a8718a68ef93fd2e356;
reg  [ 0:0]                      sgnprod_00159;
reg  [MAX_SUM_WDTH_L-1:0]        I9dc297ad41fafcda77f5347f331cfc25;
wire  [MAX_SUM_WDTH_L-1:0]       I1731c0e3be86eec142c3732ee836e4d5;
wire  [MAX_SUM_WDTH_L-1:0]       Id3b8c0ca32331f94fd98c8dae72bb15d;
wire  [MAX_SUM_WDTH_L-1:0]       I6a86b0a82441c6c14436a3e0af6b0fb7;
wire  [MAX_SUM_WDTH_L-1:0]       I8c92ff598084da7a50f7c68da96620b3;
reg  [ 0:0]                      sgnprod_00160;
reg  [MAX_SUM_WDTH_L-1:0]        I846700c79f30ca954cc2933fc94d355b;
wire  [MAX_SUM_WDTH_L-1:0]       I8bd1862e7bc2e83e9863389d532e6623;
wire  [MAX_SUM_WDTH_L-1:0]       I8053269f8bd78a931878c8350693e1d6;
wire  [MAX_SUM_WDTH_L-1:0]       I2ff66cdd7314276232715ef2361ad184;
wire  [MAX_SUM_WDTH_L-1:0]       Icf541c76bfaf37fe6111de037d205f15;
reg  [ 0:0]                      sgnprod_00161;
reg  [MAX_SUM_WDTH_L-1:0]        I8af96a91457316e49e3f7dd5e57c82da;
wire  [MAX_SUM_WDTH_L-1:0]       I68319c8b9febef9f564832429c91b85a;
wire  [MAX_SUM_WDTH_L-1:0]       I127772614218dd7c50d3136b4f174d7a;
wire  [MAX_SUM_WDTH_L-1:0]       Ib8d1aea4ad24c6ceb44f2cc672e1ff90;
wire  [MAX_SUM_WDTH_L-1:0]       I9ca26c8104bf15f48b19dc3256914544;
reg  [ 0:0]                      sgnprod_00162;
reg  [MAX_SUM_WDTH_L-1:0]        I7d1c247500d7d32e406b2a5f7e2b745b;
wire  [MAX_SUM_WDTH_L-1:0]       Icc76d9ffc3f3d7b410205eeb8232a33b;
wire  [MAX_SUM_WDTH_L-1:0]       I7fc4551d8a0445f79b87b4ba5f2ffeaa;
wire  [MAX_SUM_WDTH_L-1:0]       I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8;
wire  [MAX_SUM_WDTH_L-1:0]       Ie34c07af9f6adb9e4b636dce3d0682c0;
reg  [ 0:0]                      sgnprod_00163;
reg  [MAX_SUM_WDTH_L-1:0]        I66d85c030a8864505298919046056305;
wire  [MAX_SUM_WDTH_L-1:0]       Ib869a349250a765d2f8660e0dbdcf312;
wire  [MAX_SUM_WDTH_L-1:0]       I1a4fb631fdc7b5454c266589962ff5f0;
wire  [MAX_SUM_WDTH_L-1:0]       I9de4e0e86e9edcf948d9eddf0401b94a;
wire  [MAX_SUM_WDTH_L-1:0]       Iee7b4838986c962969c00a0bbe53ce0b;
reg  [ 0:0]                      sgnprod_00164;
reg  [MAX_SUM_WDTH_L-1:0]        I4841257ae596d9d3e4eb1e6f886956b0;
wire  [MAX_SUM_WDTH_L-1:0]       Id81b11a8ca1dd8989e36cef637ae6aab;
wire  [MAX_SUM_WDTH_L-1:0]       Ibe96deab015b799fe7f69bae8432952c;
wire  [MAX_SUM_WDTH_L-1:0]       I986b52155cc1470299321a4933241ed7;
wire  [MAX_SUM_WDTH_L-1:0]       I04be63a04f3942ce749cc9bd7540e055;
reg  [ 0:0]                      sgnprod_00165;
reg  [MAX_SUM_WDTH_L-1:0]        Icd6f7ec117f9ab4eda8c5eba41386ffa;
wire  [MAX_SUM_WDTH_L-1:0]       Ia7adea5b0ec86e9fcd427a5468d72b64;
wire  [MAX_SUM_WDTH_L-1:0]       Ie8990d8abd23f8f9f79d7fe38c57fa8c;
wire  [MAX_SUM_WDTH_L-1:0]       I9d2f90ddddbdbb525d5f070f32546b64;
wire  [MAX_SUM_WDTH_L-1:0]       I905256d73bdb63bf860e15687350795f;
reg  [ 0:0]                      sgnprod_00166;
reg  [MAX_SUM_WDTH_L-1:0]        Ibc0498839d1d9b6dc853b8e5d7a88fa3;
wire  [MAX_SUM_WDTH_L-1:0]       I9adcfc18e4471209edbe9a379e996067;
wire  [MAX_SUM_WDTH_L-1:0]       I3d7d048348bf833f744a9f73889b7802;
wire  [MAX_SUM_WDTH_L-1:0]       Id619e8d4040014d0e415ff71c5e0591f;
wire  [MAX_SUM_WDTH_L-1:0]       Iaf3de2ef283e03dd72002026e1299224;
reg  [ 0:0]                      sgnprod_00167;
reg  [MAX_SUM_WDTH_L-1:0]        I142ebca7f155e287e38ddf45423ab0fd;
wire  [MAX_SUM_WDTH_L-1:0]       I64551529c0028ec145407be7f5dfef71;
wire  [MAX_SUM_WDTH_L-1:0]       I5ebe580a943b65fb16ea722ba101fd05;
wire  [MAX_SUM_WDTH_L-1:0]       I0921901599c43b27e701758026dd3ee1;
wire  [MAX_SUM_WDTH_L-1:0]       I6033532f27c26b2d42bb3ea128f80dfa;

reg  [MAX_SUM_WDTH_L-1:0]        I5deafec6e5f32da1bcf8f7018cf794d8;
reg  [MAX_SUM_WDTH_L-1:0]        I35b3fb2670f3a60d165c1fd10f02c00c;
reg  [MAX_SUM_WDTH_L-1:0]        I68925439e233444a4da44871f31de94a;
reg  [MAX_SUM_WDTH_L-1:0]        I3108702b5ca506422c1ba6174619f193;
reg  [MAX_SUM_WDTH_L-1:0]        Icc8e8f6446ac64350a05f5e1e0541bb9;
reg  [MAX_SUM_WDTH_L-1:0]        Iadebaf3f6cca1ba78feab50ce70c8aef;
reg  [MAX_SUM_WDTH_L-1:0]        I8681cf376dbeceab29279a7637249e7d;
reg  [MAX_SUM_WDTH_L-1:0]        Ie850a07565bed90389bb125ddcd39658;
reg  [MAX_SUM_WDTH_L-1:0]        I97b77743c2311ec629ea24c933b60053;
reg  [MAX_SUM_WDTH_L-1:0]        I07a0a8d41ed8176e92380f2c89c2afdd;
reg  [MAX_SUM_WDTH_L-1:0]        I021842328f948a94159b32903c8bcb68;
reg  [MAX_SUM_WDTH_L-1:0]        Icaf3bd685005a05c8fb334266ea4e4b9;
reg  [MAX_SUM_WDTH_L-1:0]        I92d9e1d7dcf45a4d738c546e959687c3;
reg  [MAX_SUM_WDTH_L-1:0]        I39ca3a8ca714a9726114326ae6bfab0a;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9ae20ed5b2a0cad2c37c5bb2ea05ff4;
reg  [MAX_SUM_WDTH_L-1:0]        I8f131eb6138c23fdcb35195703131e64;
reg  [MAX_SUM_WDTH_L-1:0]        Iff77e08da4bcbb85b95fa277b69653a9;
reg  [MAX_SUM_WDTH_L-1:0]        I703e0a4879a39b3b8b0a49de86ca4ff4;
reg  [MAX_SUM_WDTH_L-1:0]        I3da217f6f2d0f515bb9036673d753a88;
reg  [MAX_SUM_WDTH_L-1:0]        Ifcc06d5a010e01a781ae8a9e9e2b31a0;
reg  [MAX_SUM_WDTH_L-1:0]        I42fd611fec087113ba6e35f281bced9c;
reg  [MAX_SUM_WDTH_L-1:0]        I5bb626e7347bb9ae4219cc72244b38f8;
reg  [MAX_SUM_WDTH_L-1:0]        I47e2dac0068652338f94ddffd2dbe88a;
reg  [MAX_SUM_WDTH_L-1:0]        I59a3f06de2984078a4d4c430a2980fe3;
reg  [MAX_SUM_WDTH_L-1:0]        I857b7fd58279b1063a06a4f33b880ba6;
reg  [MAX_SUM_WDTH_L-1:0]        I3901bbda029cd0a41640001c1efd400f;
reg  [MAX_SUM_WDTH_L-1:0]        Ifceeccf10f1d85a32f70c04654a1a1b4;
reg  [MAX_SUM_WDTH_L-1:0]        I2d810c1d1304658edff74921e8d0f388;
reg  [MAX_SUM_WDTH_L-1:0]        I575b0201be445388607ab83465eab8d6;
reg  [MAX_SUM_WDTH_L-1:0]        I7928c5ce0f821df1cb6271d15e19fa22;
reg  [MAX_SUM_WDTH_L-1:0]        I12695a21c942d02a432cf6382d7d7452;
reg  [MAX_SUM_WDTH_L-1:0]        I00d03f0f71b008dad8035bbf251f41bf;
reg  [MAX_SUM_WDTH_L-1:0]        I41afedcbc0f492e3243436cbefdaf609;
reg  [MAX_SUM_WDTH_L-1:0]        I638c4c2708e437a050ed7cbbac516a59;
reg  [MAX_SUM_WDTH_L-1:0]        I6877d3306b1f08c236b5d1b59f0de259;
reg  [MAX_SUM_WDTH_L-1:0]        Ib3e66aa460f39d32110ea6f115785b3d;
reg  [MAX_SUM_WDTH_L-1:0]        I5e603e8392a5322951b3225b65b19446;
reg  [MAX_SUM_WDTH_L-1:0]        If5da7fa1a615e1122445460e33487772;
reg  [MAX_SUM_WDTH_L-1:0]        Ic4153dafafaf7d047478c5d81109437f;
reg  [MAX_SUM_WDTH_L-1:0]        I7b5476007f04e81afc0125e6a8930303;
reg  [MAX_SUM_WDTH_L-1:0]        I3521a18022925249caddb8e37d2c1262;
reg  [MAX_SUM_WDTH_L-1:0]        Ifd0f52d4f814e2bb4c3bd34c1e09bda7;
reg  [MAX_SUM_WDTH_L-1:0]        I8945f6d420c8b373225451defcd2c805;
reg  [MAX_SUM_WDTH_L-1:0]        Ieec6cb6518cc0d9300de0c4f2d32487d;
reg  [MAX_SUM_WDTH_L-1:0]        Ic62eb7e90d703ef994e68587345a4293;
reg  [MAX_SUM_WDTH_L-1:0]        Id3efd8419da986aa89b8ad8e75848cfa;
reg  [MAX_SUM_WDTH_L-1:0]        I40803f10b7c4dc9ae4969739349b0265;
reg  [MAX_SUM_WDTH_L-1:0]        I7d961743fdeaf1e72e4b25c12a1d4c46;
reg  [MAX_SUM_WDTH_L-1:0]        Ifea156f33eb61fece272efe379327f6e;
reg  [MAX_SUM_WDTH_L-1:0]        Ifc99169b3399f3d14121c1a9bce3fc21;
reg  [MAX_SUM_WDTH_L-1:0]        I6536144383cbda6f3b3c564391866906;
reg  [MAX_SUM_WDTH_L-1:0]        Ic21bf9a8a4cd85ec123d7fe142ed49c0;
reg  [MAX_SUM_WDTH_L-1:0]        I1f31fe6a0ca8510bcadbc2069403150b;
reg  [MAX_SUM_WDTH_L-1:0]        I0e40933d00f4a7d9b53b2764aa0da700;
reg  [MAX_SUM_WDTH_L-1:0]        Ic41a6e00bc84bfc1b8194d15bb899c93;
reg  [MAX_SUM_WDTH_L-1:0]        I2832571f2b0a7fbb41d2e8ca7f64e003;
reg  [MAX_SUM_WDTH_L-1:0]        I9593c853e41952e408a809cb24efa4fd;
reg  [MAX_SUM_WDTH_L-1:0]        I6edffbf4136e193dca0fcec3a74e8e9c;
reg  [MAX_SUM_WDTH_L-1:0]        Ibaed50cc2e36ae58945887d11a6ec9e4;
reg  [MAX_SUM_WDTH_L-1:0]        Ie4570cac44f59e6ff46f73a703026479;
reg  [MAX_SUM_WDTH_L-1:0]        Ibaa136d37936687e9dbe4222749d19c3;
reg  [MAX_SUM_WDTH_L-1:0]        If85de3225f45478827b43b89089cd29e;
reg  [MAX_SUM_WDTH_L-1:0]        I0344b86a6e9c036e103a9c1f3651175f;
reg  [MAX_SUM_WDTH_L-1:0]        I5463d13575e0b9fb8a0f6cc8b35d0ce9;
reg  [MAX_SUM_WDTH_L-1:0]        I8a3c63ef122001a29e5abe93c4e1a48f;
reg  [MAX_SUM_WDTH_L-1:0]        I6a79108484fcb192f6d93bfb98e271c4;
reg  [MAX_SUM_WDTH_L-1:0]        I9001e95b71457a2bd09a9846af370b16;
reg  [MAX_SUM_WDTH_L-1:0]        I51620de618db6327358a5cac97e1e97f;
reg  [MAX_SUM_WDTH_L-1:0]        Ib9c58818059af5c5a03e77a5dcef4654;
reg  [MAX_SUM_WDTH_L-1:0]        I8081c71aa01a8d575bfea6ea7f2f595f;
reg  [MAX_SUM_WDTH_L-1:0]        Iad999607ad8d7da0f3b341f83ea030a6;
reg  [MAX_SUM_WDTH_L-1:0]        Ie7291c914d2cb66f547b0a7717f71311;
reg  [MAX_SUM_WDTH_L-1:0]        Ic01018a5f1bc392bbd267016f6612a83;
reg  [MAX_SUM_WDTH_L-1:0]        Ib11dff839e7e532657b32f29fd9b1651;
reg  [MAX_SUM_WDTH_L-1:0]        I251d7ea16dd5407d22a6846ddcfe12d8;
reg  [MAX_SUM_WDTH_L-1:0]        I773797f81f73b9b6e844441142a1bb48;
reg  [MAX_SUM_WDTH_L-1:0]        I853ecadf30fc10a13dd1ffb1f2dfb5d6;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb8b3c91e1d3b890cfe58f32f8ec3ae3;
reg  [MAX_SUM_WDTH_L-1:0]        I3485d69de942d64e56925da522175b51;
reg  [MAX_SUM_WDTH_L-1:0]        Iae42f12bc0475c8b58341d80027a57cb;
reg  [MAX_SUM_WDTH_L-1:0]        I22fe2af25463f87ee7315a9aac32854e;
reg  [MAX_SUM_WDTH_L-1:0]        Idf44ad78c338c39699721ce511691dfd;
reg  [MAX_SUM_WDTH_L-1:0]        I984a657f9265d41318c0290e249e9712;
reg  [MAX_SUM_WDTH_L-1:0]        I915fccfb1d1ada9aa7c8e24c2eebd04c;
reg  [MAX_SUM_WDTH_L-1:0]        I2bdf58ecd0974720631be830efb48dc8;
reg  [MAX_SUM_WDTH_L-1:0]        Ibaedf6246fa43acc8accb5a24d49cc2f;
reg  [MAX_SUM_WDTH_L-1:0]        I904d13524dcdf55478a5266d50e53ff7;
reg  [MAX_SUM_WDTH_L-1:0]        I22d8e5d57c1bc082169437a654d22bba;
reg  [MAX_SUM_WDTH_L-1:0]        I719cdaa2a2e61a0df7f1fd5efe517426;
reg  [MAX_SUM_WDTH_L-1:0]        I8e92a61eb73c41680652936cfcc614ff;
reg  [MAX_SUM_WDTH_L-1:0]        I7ad5af8319f6da469858300f0777b580;
reg  [MAX_SUM_WDTH_L-1:0]        I32be72eaf04e79120a57ea94296a4e56;
reg  [MAX_SUM_WDTH_L-1:0]        Ie756f6a87d85adb40479ce7cf3545556;
reg  [MAX_SUM_WDTH_L-1:0]        I8794c6ce0a3f2e6697372e2c911ba420;
reg  [MAX_SUM_WDTH_L-1:0]        Ic82b1a29b5e63bcc3686a0d4bf1f5c24;
reg  [MAX_SUM_WDTH_L-1:0]        I253ef976058080beab79646af18e2d5b;
reg  [MAX_SUM_WDTH_L-1:0]        I930dd54c36540d75dc870eef89960163;
reg  [MAX_SUM_WDTH_L-1:0]        Iaf7554cd4e8b5ea6155ec61a8d589b86;
reg  [MAX_SUM_WDTH_L-1:0]        I50907c7d1efa0038d81efed82b192891;
reg  [MAX_SUM_WDTH_L-1:0]        If3e9486d2960d164d94641d4f1917416;
reg  [MAX_SUM_WDTH_L-1:0]        I2bec61db45dd79b98d6ebff6c5a4899e;
reg  [MAX_SUM_WDTH_L-1:0]        I7f31647f3ea6ce7bbd211c25cf4828fb;
reg  [MAX_SUM_WDTH_L-1:0]        Ice65387e606faf9c7b884475b489abba;
reg  [MAX_SUM_WDTH_L-1:0]        I63f914927dcf49552e9f3fe0180a30e8;
reg  [MAX_SUM_WDTH_L-1:0]        I742ff5725e3a18acd03454cf9f313f4b;
reg  [MAX_SUM_WDTH_L-1:0]        I84e4b3bc63ec0b0bff7f98f433c1fd67;
reg  [MAX_SUM_WDTH_L-1:0]        I78c6a1428a1f211c5e89b8c76b3dc033;
reg  [MAX_SUM_WDTH_L-1:0]        I9897cbf9d7cab759f99f5f8f4bc125d0;
reg  [MAX_SUM_WDTH_L-1:0]        I9a6c1ff6dde5141849e4aa925140ebb8;
reg  [MAX_SUM_WDTH_L-1:0]        Icc1c25b229393361f1245c40f573b423;
reg  [MAX_SUM_WDTH_L-1:0]        I53b5a72e41ee53037ee3ae040799f401;
reg  [MAX_SUM_WDTH_L-1:0]        I3cc25fb583118f45babf457fe78d5434;
reg  [MAX_SUM_WDTH_L-1:0]        I20c046dd8a1265e12e902275b73417da;
reg  [MAX_SUM_WDTH_L-1:0]        I1b184c9a34aeb6eda813d86556e235d9;
reg  [MAX_SUM_WDTH_L-1:0]        I70e03db993e1d26d5814ff5fcd38ada1;
reg  [MAX_SUM_WDTH_L-1:0]        I119dc168a44950d215af877eb81152fe;
reg  [MAX_SUM_WDTH_L-1:0]        Id717ed42457eb1d3f4e3edbf0dd72c41;
reg  [MAX_SUM_WDTH_L-1:0]        I79d1f852a03bcc11d6121a12d8c5b86d;
reg  [MAX_SUM_WDTH_L-1:0]        I769e650e49f152c0803b06232740691c;
reg  [MAX_SUM_WDTH_L-1:0]        I1ef3c09b8481f14c3526224430a5f4b9;
reg  [MAX_SUM_WDTH_L-1:0]        I2a38d43a7e25050aa672cbf84a409aa8;
reg  [MAX_SUM_WDTH_L-1:0]        I1c2be5e13c462a8a6b07bca311582ce4;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8fd61caf16aa0e504cc7dc8cec6f0b8;
reg  [MAX_SUM_WDTH_L-1:0]        Icd0fe98ca873ad6dacdf80dfdfc450ec;
reg  [MAX_SUM_WDTH_L-1:0]        I94e1ab698dc93ff0764dc5c1e62179fe;
reg  [MAX_SUM_WDTH_L-1:0]        Ifd48363af9abb390a72991fbdd6f7877;
reg  [MAX_SUM_WDTH_L-1:0]        I44f79397a010088e4ecdcb9669f2efbd;
reg  [MAX_SUM_WDTH_L-1:0]        I124b0b7d91cfb42b0d9722f3229c2d53;
reg  [MAX_SUM_WDTH_L-1:0]        Iadf1875c584adc34f7586a146184a763;
reg  [MAX_SUM_WDTH_L-1:0]        I02d3f9982f02ea85f996bf5b5975b930;
reg  [MAX_SUM_WDTH_L-1:0]        Ia6e1b39d83ddce053518c5ae9a5ca33e;
reg  [MAX_SUM_WDTH_L-1:0]        I3308663053f4307d43ac66f43266f706;
reg  [MAX_SUM_WDTH_L-1:0]        I87ad25dff6c0c9ac46b7a129cb575537;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf5d40b7c46b50866f58f6fa23e1861b;
reg  [MAX_SUM_WDTH_L-1:0]        I0e3a9a3b38875156d15f697adaf95410;
reg  [MAX_SUM_WDTH_L-1:0]        Ie3f87d094e71e4a82f60e8d91cdd768b;
reg  [MAX_SUM_WDTH_L-1:0]        I793f52d174cd09fe000e8d0351753592;
reg  [MAX_SUM_WDTH_L-1:0]        I89ea3da7db40e7e6705020462b2d1df1;
reg  [MAX_SUM_WDTH_L-1:0]        Ib2af2f1a928dd824f25b99f0b602753f;
reg  [MAX_SUM_WDTH_L-1:0]        Ie3e887f5f1a64c37a10404d636212b45;
reg  [MAX_SUM_WDTH_L-1:0]        I5c6a004278f155d33d0cc1b576c3b25f;
reg  [MAX_SUM_WDTH_L-1:0]        I6a03a4a548a0906d1a3e9ce47f3454c6;
reg  [MAX_SUM_WDTH_L-1:0]        I542e525074d049197ac3904e6102f0bd;
reg  [MAX_SUM_WDTH_L-1:0]        Ie0307a43ce71ba73d4c8e5ad556bd341;
reg  [MAX_SUM_WDTH_L-1:0]        Ib03e1d3a1f27721e4ea32629c2e86f85;
reg  [MAX_SUM_WDTH_L-1:0]        I782f4ab4666c9f550a2cfc943cedbe77;
reg  [MAX_SUM_WDTH_L-1:0]        Ib991e16161d5c8b3b655e3c7c08b93c4;
reg  [MAX_SUM_WDTH_L-1:0]        I72f8c6bad4bff3b00055aa8824479931;
reg  [MAX_SUM_WDTH_L-1:0]        I58e5100cc1e9b809e93125fe5d08a9d8;
reg  [MAX_SUM_WDTH_L-1:0]        I0aa7056fdacd6022f328a3be49048856;
reg  [MAX_SUM_WDTH_L-1:0]        Ia2f40b5c49a2284fb6a234bf7472130f;
reg  [MAX_SUM_WDTH_L-1:0]        I8da184aee7953890f2c89e40744402f4;
reg  [MAX_SUM_WDTH_L-1:0]        I613ccfc7dad5627cde02fa1720244d01;
reg  [MAX_SUM_WDTH_L-1:0]        I080fc6c99e506e569b97433f3fdc3e60;
reg  [MAX_SUM_WDTH_L-1:0]        I79aa118ef8ac0d9b13723fb1f5a7e4ad;
reg  [MAX_SUM_WDTH_L-1:0]        I7e6e7601245ca5b3a58b91848e25a6d3;
reg  [MAX_SUM_WDTH_L-1:0]        I2792edda66743635b837aa3bec0c58b9;
reg  [MAX_SUM_WDTH_L-1:0]        I085cc29465c945957d00cbcf804e3ae4;
reg  [MAX_SUM_WDTH_L-1:0]        I74a8e879666bb216a331fd2ab723e37c;
reg  [MAX_SUM_WDTH_L-1:0]        I7a90a43ed71e82862457d9fa40bd005c;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1e7b4bd6201baa02b8d59cb0f6ffb8e;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7b7cdc22b22f276b1c021abaa8fb443;
reg  [MAX_SUM_WDTH_L-1:0]        Ib58e33f31be36b28997ba05ef1004573;
reg  [MAX_SUM_WDTH_L-1:0]        Ibec394e82f499e8d2d5a9524f943d6ac;
reg  [MAX_SUM_WDTH_L-1:0]        Ie06ad127e475dc131859992bb5f350a0;
reg  [MAX_SUM_WDTH_L-1:0]        Ic494a58468b6a7dda76923a9475bf173;
reg  [MAX_SUM_WDTH_L-1:0]        Ib82a2db86d03fe8538fa19d06e501dae;
reg  [MAX_SUM_WDTH_L-1:0]        I5b64727fee9d0825a4ea83261992e489;
reg  [MAX_SUM_WDTH_L-1:0]        Ice7e502b9c2b797719448fde8376087a;
reg  [MAX_SUM_WDTH_L-1:0]        I792b4f73ed7139b8761443cbc0833e39;
reg  [MAX_SUM_WDTH_L-1:0]        I278d57d1964cbf3339db450926ef4782;
reg  [MAX_SUM_WDTH_L-1:0]        I9c1a08b61782ef6c72545504693ac54e;
reg  [MAX_SUM_WDTH_L-1:0]        I363594fb91d01abca7a2b7402e352fd0;
reg  [MAX_SUM_WDTH_L-1:0]        Idd284c75a230f4b97d5acb98a8e38b2d;
reg  [MAX_SUM_WDTH_L-1:0]        If040df53a6410b263f5b3dc3090631c4;
reg  [MAX_SUM_WDTH_L-1:0]        I31df60ffcaea9cee63b920478cb058f1;
reg  [MAX_SUM_WDTH_L-1:0]        Icdd2f6ce69b389fbf712e45bdc0a0257;
reg  [MAX_SUM_WDTH_L-1:0]        I8971b250393b397b94db38b9fd0fe501;
reg  [MAX_SUM_WDTH_L-1:0]        I9199e5e8fdc0e2c62ad1d62fc4d873cb;
reg  [MAX_SUM_WDTH_L-1:0]        I6e03f71fdf20db836c5772658a050e9c;
reg  [MAX_SUM_WDTH_L-1:0]        I2ef49f893dbc8581725ca0f6d1c3305c;
reg  [MAX_SUM_WDTH_L-1:0]        I8796f168c892ac60c38a0a7f1e18035e;
reg  [MAX_SUM_WDTH_L-1:0]        I64a26e5117c8f3ab95bf0dfa97427243;
reg  [MAX_SUM_WDTH_L-1:0]        Id7946a0299ced3ba00f6c3e6e664931f;
reg  [MAX_SUM_WDTH_L-1:0]        I5243b90640ea4680de83021601c85c39;
reg  [MAX_SUM_WDTH_L-1:0]        Ic8301fceed328cc031640ecc4ff34803;
reg  [MAX_SUM_WDTH_L-1:0]        I6e852c94b6105af62ee85f8adf77fa55;
reg  [MAX_SUM_WDTH_L-1:0]        I7d98c5c2a54832b6368ce60009208eb0;
reg  [MAX_SUM_WDTH_L-1:0]        I7e42f2281518bead81a6d18d2dcbd1a3;
reg  [MAX_SUM_WDTH_L-1:0]        I63c126c978154f2d68b11f08a938dcb4;
reg  [MAX_SUM_WDTH_L-1:0]        I2ff7719c35578b47720cacd9ddfd92eb;
reg  [MAX_SUM_WDTH_L-1:0]        I480599aef36967a670155dd77120a37d;
reg  [MAX_SUM_WDTH_L-1:0]        Ic000b2c844de484b8f30b7b84dd6234d;
reg  [MAX_SUM_WDTH_L-1:0]        If0e25df151db991185f992eab5d5be99;
reg  [MAX_SUM_WDTH_L-1:0]        I2f533699abb7a997160bf4ee4cda3efb;
reg  [MAX_SUM_WDTH_L-1:0]        If6b33cfc6d34e33fbb18e08fb4d8a5ed;
reg  [MAX_SUM_WDTH_L-1:0]        I2ea5423dc8726fc0217899e0f406a1e9;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf3f4f8a04cbacc9624ca5cc73bf7069;
reg  [MAX_SUM_WDTH_L-1:0]        I9ba53c36934ab1c7f498241a79cfbae8;
reg  [MAX_SUM_WDTH_L-1:0]        I106a25f18536f96782927bf3bc2ccd72;
reg  [MAX_SUM_WDTH_L-1:0]        Ie5cdad65e918679607cc5f816987b736;
reg  [MAX_SUM_WDTH_L-1:0]        Ica6dc9ded8756fd6f82eec4271e246c3;
reg  [MAX_SUM_WDTH_L-1:0]        Ica42ac6ca5813d0d1a67f14d1248437a;
reg  [MAX_SUM_WDTH_L-1:0]        I13dc6cfc75ef846c30e5dc1dc5305d59;
reg  [MAX_SUM_WDTH_L-1:0]        I33e784182dfb4af39715788b1ae98af6;
reg  [MAX_SUM_WDTH_L-1:0]        I9e1a66805348d2e5bbf5e2316187444b;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9619916a96d218cf5eb5f3a4995d0e7;
reg  [MAX_SUM_WDTH_L-1:0]        I02ce7969c51ad141df227ed7d18e74b1;
reg  [MAX_SUM_WDTH_L-1:0]        Idd73461af0d75c4d820f7f8f0f419e0f;
reg  [MAX_SUM_WDTH_L-1:0]        I3df6c2cdccb2a82c58c1d81b00af7786;
reg  [MAX_SUM_WDTH_L-1:0]        I97f441fc5ffb88efeb5ed66b60f07a7c;
reg  [MAX_SUM_WDTH_L-1:0]        I3194a235eb652c8d0e4307cd056e5e72;
reg  [MAX_SUM_WDTH_L-1:0]        Ibc315f6c79ba2bf336ee57f2e5f7d776;
reg  [MAX_SUM_WDTH_L-1:0]        I937a54f5cda99a7079c7fa46b4ea26f6;
reg  [MAX_SUM_WDTH_L-1:0]        I49c99afecc613656cd1469d8c1e98936;
reg  [MAX_SUM_WDTH_L-1:0]        Id76ce0333f43bf7bccf1ce48e25ca69c;
reg  [MAX_SUM_WDTH_L-1:0]        I2c77f9644145219005751f7a4eb71aaa;
reg  [MAX_SUM_WDTH_L-1:0]        I5cecc266272eef88cda88c1df9bcc37e;
reg  [MAX_SUM_WDTH_L-1:0]        I776a0b1b5c14afa21b7fda3c2cacafed;
reg  [MAX_SUM_WDTH_L-1:0]        I84860b1f933339e0f90beeb3d666393b;
reg  [MAX_SUM_WDTH_L-1:0]        Id24581713f1ecb767db39d5154c2f5f4;
reg  [MAX_SUM_WDTH_L-1:0]        Idb0eae2f0e1dae1d56251d64e2c51f9f;
reg  [MAX_SUM_WDTH_L-1:0]        I2e3ca4b130e6d3d92385928a28644452;
reg  [MAX_SUM_WDTH_L-1:0]        I7922d80ae333dcfafde31d294f0eb4d8;
reg  [MAX_SUM_WDTH_L-1:0]        I82de04cd2dfef5616efca4af26d7c561;
reg  [MAX_SUM_WDTH_L-1:0]        I7ce384520525b15d24c2ef6f161213a5;
reg  [MAX_SUM_WDTH_L-1:0]        I56aeea71c7bd19d47620cf36adf3f115;
reg  [MAX_SUM_WDTH_L-1:0]        I138e1a6db0c6649bc023cc36d81d5b47;
reg  [MAX_SUM_WDTH_L-1:0]        Ib5e8b1c4dd9b5dad56b59cc11c87a258;
reg  [MAX_SUM_WDTH_L-1:0]        I86f785e2d5e8d6c08fad1d334c7d244e;
reg  [MAX_SUM_WDTH_L-1:0]        I9a6c8efca218c724da4ee4c1087d58bc;
reg  [MAX_SUM_WDTH_L-1:0]        Ia30e8dbc6974ea94b763842e8dffa633;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa60f45f4d8848eb0b89f5644ec69668;
reg  [MAX_SUM_WDTH_L-1:0]        I0aeb4b93cfa6d62ec41b7e6dd0287dd0;
reg  [MAX_SUM_WDTH_L-1:0]        Ifce1fc978fb5b0187593f46f53c3b469;
reg  [MAX_SUM_WDTH_L-1:0]        If3b6de7c919c5d53a0e191a75bd7e574;
reg  [MAX_SUM_WDTH_L-1:0]        Iecce594e6e99b0c05fc845144a664b07;
reg  [MAX_SUM_WDTH_L-1:0]        I2c8431500ecb25619d2884a2fb4260c0;
reg  [MAX_SUM_WDTH_L-1:0]        I217c710f7ef39035546efcbb043f63f3;
reg  [MAX_SUM_WDTH_L-1:0]        I1b4236130cb1879d885653fdd9eeab4e;
reg  [MAX_SUM_WDTH_L-1:0]        Iae0f7c13f1564d63b4bfdc152ddf4111;
reg  [MAX_SUM_WDTH_L-1:0]        I010592496030d138a3a4245d00069957;
reg  [MAX_SUM_WDTH_L-1:0]        I9d7f47a6289a16448221d61f301586aa;
reg  [MAX_SUM_WDTH_L-1:0]        I7b8ed2953170c4deadaeb33a6ba165d4;
reg  [MAX_SUM_WDTH_L-1:0]        I4efe9eef6a48aeb0a9ba4e0ffd9906c3;
reg  [MAX_SUM_WDTH_L-1:0]        I5a8466bbd83c39dfbeaa6399e3fb3337;
reg  [MAX_SUM_WDTH_L-1:0]        I1ab96ffa948dd09bcc4f748c6c2575d2;
reg  [MAX_SUM_WDTH_L-1:0]        I016f57568eaf00b26f8a22100858c158;
reg  [MAX_SUM_WDTH_L-1:0]        I1fb995e302f4f1ba493ff85f39938175;
reg  [MAX_SUM_WDTH_L-1:0]        Ie643ad235307c60f1ee96dfdcbc8c2a8;
reg  [MAX_SUM_WDTH_L-1:0]        I8dafdf2c780082d8dfc2961b3447f104;
reg  [MAX_SUM_WDTH_L-1:0]        I3a2841a0f5e1b42556f384231ab0717b;
reg  [MAX_SUM_WDTH_L-1:0]        I2b00d0e6facf01274c0c3446bb0e1599;
reg  [MAX_SUM_WDTH_L-1:0]        I2c645d25871b70dae5b2c283695d5130;
reg  [MAX_SUM_WDTH_L-1:0]        I540a0e8968a6a82aca775a81ef82b520;
reg  [MAX_SUM_WDTH_L-1:0]        I5b95bbc82e6d8d87421efe3f17b97ea5;
reg  [MAX_SUM_WDTH_L-1:0]        Iad81f5e5e728ffdec6296b2aff668d75;
reg  [MAX_SUM_WDTH_L-1:0]        I960a618f63372da74581b8c352f3e618;
reg  [MAX_SUM_WDTH_L-1:0]        I4f5325f1601acde10018d1fd0aff4d35;
reg  [MAX_SUM_WDTH_L-1:0]        Ib297101fe456520e72cd9d208af44eea;
reg  [MAX_SUM_WDTH_L-1:0]        I73a21342321a9d81a0fa5308149d72b0;
reg  [MAX_SUM_WDTH_L-1:0]        I2a486524f4f53b3454ee02a8892d4fa3;
reg  [MAX_SUM_WDTH_L-1:0]        Ic6c4e4e6a9ba43a3354f9f3192ab069e;
reg  [MAX_SUM_WDTH_L-1:0]        Ie3cdee3560bd06aed84dac5fcd2a259a;
reg  [MAX_SUM_WDTH_L-1:0]        I584febaa4c440fd9353108af36d3a5c6;
reg  [MAX_SUM_WDTH_L-1:0]        I515e78507d7419ca14d77b6d52f75a78;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9578453a57d2b3b9c3b98844044b5f0;
reg  [MAX_SUM_WDTH_L-1:0]        I1e58b3062097a46d8d590232b40278cf;
reg  [MAX_SUM_WDTH_L-1:0]        I3af126eb28c67797ce625b0d82943833;
reg  [MAX_SUM_WDTH_L-1:0]        I130ee1a8acacf4cae8818cd8320d050d;
reg  [MAX_SUM_WDTH_L-1:0]        Idf92dd09c29ce8e921b2b34089550586;
reg  [MAX_SUM_WDTH_L-1:0]        Iba74a64cc1d2ec3c83a4061db298ad37;
reg  [MAX_SUM_WDTH_L-1:0]        I01364c233ca541914d790354515aa5c1;
reg  [MAX_SUM_WDTH_L-1:0]        Ic6a8297308a63ed3113008a3cdc76358;
reg  [MAX_SUM_WDTH_L-1:0]        I6c7ee9d0bd684a7f54bed3d52452219d;
reg  [MAX_SUM_WDTH_L-1:0]        I985ea87550ec8a222e6af621589e186d;
reg  [MAX_SUM_WDTH_L-1:0]        I6836a7d1e006d7f7556edf8b31aea32e;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7a356a18af18ec131b9df46019f3e58;
reg  [MAX_SUM_WDTH_L-1:0]        If3a7e111247232c47ceccb5e05338312;
reg  [MAX_SUM_WDTH_L-1:0]        I5f38d1665294b2d3c18f9cd888ff60f1;
reg  [MAX_SUM_WDTH_L-1:0]        I10290b9576bf3d8caf90583a388226b7;
reg  [MAX_SUM_WDTH_L-1:0]        Ief36236305fc1521c5bb4c60753a676a;
reg  [MAX_SUM_WDTH_L-1:0]        Ibaa0539fbf5ccc979511c09c061cf494;
reg  [MAX_SUM_WDTH_L-1:0]        I95664ffd0ff13c2893421032149f24d2;
reg  [MAX_SUM_WDTH_L-1:0]        Ie390153b3b7985dc63d65913de215377;
reg  [MAX_SUM_WDTH_L-1:0]        I704147dda658f4a03627dacc1c91dd48;
reg  [MAX_SUM_WDTH_L-1:0]        Ifb09672d505898f081aa13c95fcb88b5;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb5cb89097dd11bf292d5b5a2422175b;
reg  [MAX_SUM_WDTH_L-1:0]        I4a305956b18d6ad6901d2c17e99f2bab;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf5bb3b9eb1812383db9634fa9a27ad3;
reg  [MAX_SUM_WDTH_L-1:0]        I66b37d055c3735f011095ee4b1ad02ed;
reg  [MAX_SUM_WDTH_L-1:0]        I43e71dd694d97217e242f267248cd594;
reg  [MAX_SUM_WDTH_L-1:0]        I4baa925db1ec733bd4bd25d9dc873e23;
reg  [MAX_SUM_WDTH_L-1:0]        I547928c9db7acc531af251264d576ffb;
reg  [MAX_SUM_WDTH_L-1:0]        Ie4ce634b2fb62a20781f8a2e8fddc762;
reg  [MAX_SUM_WDTH_L-1:0]        I0e90e96ffa64c2874d79110b622994bf;
reg  [MAX_SUM_WDTH_L-1:0]        I767e37e3c6f4224eb07adeda480ce253;
reg  [MAX_SUM_WDTH_L-1:0]        I75fcaf2c65b7e63adac834054850c6d6;
reg  [MAX_SUM_WDTH_L-1:0]        I5f1de2dfbd79204ab2db9b686d6a6862;
reg  [MAX_SUM_WDTH_L-1:0]        I8d01de6be4091dca2589cef625c05229;
reg  [MAX_SUM_WDTH_L-1:0]        Ic09e773899fdd208c0fdd874933b2cec;
reg  [MAX_SUM_WDTH_L-1:0]        I24a3f9fd851c4af70ef66bfcee44af65;
reg  [MAX_SUM_WDTH_L-1:0]        Idd31807ecd603db8c719349a2be1be40;
reg  [MAX_SUM_WDTH_L-1:0]        Iaf680cae40d1adf7649da12b31a2be0d;
reg  [MAX_SUM_WDTH_L-1:0]        I22d948171c1a66f7a28d5e51007700ea;
reg  [MAX_SUM_WDTH_L-1:0]        I3954318b2392a82f2da71a0ca1504497;
reg  [MAX_SUM_WDTH_L-1:0]        I15c78b909cbd04fe25820d777655d829;
reg  [MAX_SUM_WDTH_L-1:0]        Ia529c5ec88a9f6c14ceda5cad56b346d;
reg  [MAX_SUM_WDTH_L-1:0]        I5b73c81f28901705f6ee26d63847db0a;
reg  [MAX_SUM_WDTH_L-1:0]        I1a9bd3f728db23b679639e5657ced179;
reg  [MAX_SUM_WDTH_L-1:0]        I57ca72784a7c91cecbd694ddd08bcb98;
reg  [MAX_SUM_WDTH_L-1:0]        I50f31ecd3f2b498cc7b759efa057f12f;
reg  [MAX_SUM_WDTH_L-1:0]        I8ccaf29848defdd264f522642968fa29;
reg  [MAX_SUM_WDTH_L-1:0]        I808ea92ee1340876cf1d2c47255dc2fe;
reg  [MAX_SUM_WDTH_L-1:0]        I3da806790125328b626be1949f71267a;
reg  [MAX_SUM_WDTH_L-1:0]        I55e59bc1daeb8b2be3d7a1e4b272df93;
reg  [MAX_SUM_WDTH_L-1:0]        Ib0ffadc6a0091ceff91ad1fa435413a6;
reg  [MAX_SUM_WDTH_L-1:0]        Ic863f139e6bed2d06789a07c6dedf6f8;
reg  [MAX_SUM_WDTH_L-1:0]        Id0e8f6ada5060a911090f76cfaa3c6bf;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb8c9b8fc9b58f5f8a6ad342934804a8;
reg  [MAX_SUM_WDTH_L-1:0]        I9323a188737ca54c2dd553cd99bd416c;
reg  [MAX_SUM_WDTH_L-1:0]        I2694cef38855f496e7ca12f42dfdb9fc;
reg  [MAX_SUM_WDTH_L-1:0]        I75790b4c0b1f6c7935f5cfbea26407d1;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8b366c47e56a49fc53ea4a9e1ebbd99;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1c86256df2bc6c4dad41237eca41986;
reg  [MAX_SUM_WDTH_L-1:0]        I7c9e3f97a94f9a078c209a1b84ff916d;
reg  [MAX_SUM_WDTH_L-1:0]        Idde839d34403fdbba62671b83801ea8d;
reg  [MAX_SUM_WDTH_L-1:0]        I824e23c3e43434e0a7bf8c8b8e0de597;
reg  [MAX_SUM_WDTH_L-1:0]        I0f83a2c488c229e971030fc66ce212f5;
reg  [MAX_SUM_WDTH_L-1:0]        I8fdda3dea7a63fd6e57f70365d7b6571;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa2fc30c14c549339edc65c3670d90a0;
reg  [MAX_SUM_WDTH_L-1:0]        If69bb1bfa10ca7dd37ba57485c3429e7;
reg  [MAX_SUM_WDTH_L-1:0]        I2ab0738fa2d5916d77a81b9da2315376;
reg  [MAX_SUM_WDTH_L-1:0]        I50a9ce776ad2ccd8048b56ce101c80d2;
reg  [MAX_SUM_WDTH_L-1:0]        I9c9d0332ee7ad6a3488b7e39bcb06ca2;
reg  [MAX_SUM_WDTH_L-1:0]        Idc155814976f0aef9b56b2bb3d52b3a5;
reg  [MAX_SUM_WDTH_L-1:0]        I2e02fbd496d08acb3ad3359b49b9f680;
reg  [MAX_SUM_WDTH_L-1:0]        If0f8b3dfce99a5a75c2105d45ccad985;
reg  [MAX_SUM_WDTH_L-1:0]        I6790223e6a7cf136a7e2b261ba4fdb0a;
reg  [MAX_SUM_WDTH_L-1:0]        I6a9643afea7a6cc9b94806ccc8e84c0f;
reg  [MAX_SUM_WDTH_L-1:0]        Id3d19d7c2b941930478a7ab01049e390;
reg  [MAX_SUM_WDTH_L-1:0]        Ib0a25312d51cb6aa1741f7e425bc5cd8;
reg  [MAX_SUM_WDTH_L-1:0]        I44dd1b66f5a9a6b0b976d3d61d6c5cbe;
reg  [MAX_SUM_WDTH_L-1:0]        I3ee456f2f0e7f447ae92b7523136adb5;
reg  [MAX_SUM_WDTH_L-1:0]        Ic110e2a08b550acd3c8bda4a1bc2bbae;
reg  [MAX_SUM_WDTH_L-1:0]        I3f87162d2874effd66a82f821aa6c73a;
reg  [MAX_SUM_WDTH_L-1:0]        I660ea6d341fcb38f108270c08d82473b;
reg  [MAX_SUM_WDTH_L-1:0]        Ic128d603fc08affd2f3d0ab3425710e5;
reg  [MAX_SUM_WDTH_L-1:0]        Id5372641727970383a59e08f550814b4;
reg  [MAX_SUM_WDTH_L-1:0]        Ie99ad992d66880542dcd330ef6ccee04;
reg  [MAX_SUM_WDTH_L-1:0]        I9ed0b194f7d210d57c54b289e01c75e6;
reg  [MAX_SUM_WDTH_L-1:0]        I227828831c4ad21b06ed00fb5781b0e3;
reg  [MAX_SUM_WDTH_L-1:0]        I09d5ad12cb836adfbb4833ee80fad2c9;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa9c94ee94e4beb2e7c8d2d57150df41;
reg  [MAX_SUM_WDTH_L-1:0]        Icb88e59e194db215382e8e949603a9be;
reg  [MAX_SUM_WDTH_L-1:0]        Id4ebd28aaf1076acec266666f88a02ad;
reg  [MAX_SUM_WDTH_L-1:0]        Idf0a0bd862167392357501b3233a8d8c;
reg  [MAX_SUM_WDTH_L-1:0]        If94cdb867ea0fc2c5578b16aacb1acfc;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8c066b0700941a4fa739820ff12b948;
reg  [MAX_SUM_WDTH_L-1:0]        I11e0f8dc46b286bafb05f901f968e1ad;
reg  [MAX_SUM_WDTH_L-1:0]        I608537f5639d5e0cd3e80453e21f6f85;
reg  [MAX_SUM_WDTH_L-1:0]        I0e9d8db1bb6347c9507b645132308b3a;
reg  [MAX_SUM_WDTH_L-1:0]        I17033b417fa383a2db41d157df33d9de;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7f45dbcad513b4dafee60f33622b0c3;
reg  [MAX_SUM_WDTH_L-1:0]        Ibfbd8e00e00272f32428c7b4a3c53050;
reg  [MAX_SUM_WDTH_L-1:0]        I27973d1d4e07eaa49608d6f6975d0a93;
reg  [MAX_SUM_WDTH_L-1:0]        If77fcedbcf99f89045de87e5cae45d8a;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8f8691820e7a560db8116f38dae5d49;
reg  [MAX_SUM_WDTH_L-1:0]        If0b19af59ad851aded19970494514034;
reg  [MAX_SUM_WDTH_L-1:0]        I98b8e05818925a4b65082fa57affde83;
reg  [MAX_SUM_WDTH_L-1:0]        I69317e8c556ed67630829c990f8b74db;
reg  [MAX_SUM_WDTH_L-1:0]        I9147d103cf235310393f9339f1cbb376;
reg  [MAX_SUM_WDTH_L-1:0]        Ibe0b2cab6e2d3f3cc8baf3623ff50988;
reg  [MAX_SUM_WDTH_L-1:0]        Idc64f1443dd2497dfaa223cda3fbd682;
reg  [MAX_SUM_WDTH_L-1:0]        I6e37e92b812099985436851da8a6ccb2;
reg  [MAX_SUM_WDTH_L-1:0]        I057df2bf67d5580275654bdc28b40027;
reg  [MAX_SUM_WDTH_L-1:0]        Ie87a151c8b90942a899b8167bcb34afb;
reg  [MAX_SUM_WDTH_L-1:0]        I735752035af159b48f53d8302bb33c21;
reg  [MAX_SUM_WDTH_L-1:0]        I1f26bc7cb30a9659a638e2ab65e1f187;
reg  [MAX_SUM_WDTH_L-1:0]        If39a50e88c4a7c43428c1d15b0bfbbcc;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf966c12f049d603361ad32f55b0a2c8;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1b3ed6d3fdae47669d3c4cb8af8d969;
reg  [MAX_SUM_WDTH_L-1:0]        I4ec6c8d9e87224ecbe7c69d92f9419c8;
reg  [MAX_SUM_WDTH_L-1:0]        I2acb34de8c3fc53117a7ea4f9ce7dd2b;
reg  [MAX_SUM_WDTH_L-1:0]        I7fa4009267e80ea7eb71194843c3b22b;
reg  [MAX_SUM_WDTH_L-1:0]        I6854329daadea2734e52180a41f56bcc;
reg  [MAX_SUM_WDTH_L-1:0]        Ifca16aebaf75b2990188de201e4536fd;
reg  [MAX_SUM_WDTH_L-1:0]        I46cc26afc8475f2fb290eefc95a542eb;
reg  [MAX_SUM_WDTH_L-1:0]        Id746d6515cec9e60e7478898a09787e5;
reg  [MAX_SUM_WDTH_L-1:0]        I09a3ad636db96e00adac78c3c94bdaaa;
reg  [MAX_SUM_WDTH_L-1:0]        I28b3baa225a5fd602c9fee9c948ae58b;
reg  [MAX_SUM_WDTH_L-1:0]        Ibe12ef0f56d875c7a44030882deb0e29;
reg  [MAX_SUM_WDTH_L-1:0]        I9bd9979e4acc4944227a4bd62b910c1d;
reg  [MAX_SUM_WDTH_L-1:0]        Idcfa802f458499150055dbe4b1ce8146;
reg  [MAX_SUM_WDTH_L-1:0]        Iee010958cc3e9389cb8ecacff84fccee;
reg  [MAX_SUM_WDTH_L-1:0]        I3d74b31096917c53757c829a67cf06df;
reg  [MAX_SUM_WDTH_L-1:0]        Ic27031a9654db9459815fe0ca35408db;
reg  [MAX_SUM_WDTH_L-1:0]        Idf6ead2c37f75f3cde1d4b40cd73db00;
reg  [MAX_SUM_WDTH_L-1:0]        I66a56161cd0ed67f65834b9eb0e94d17;
reg  [MAX_SUM_WDTH_L-1:0]        If6de990e26ca9e8efc009188f8a5a4d9;
reg  [MAX_SUM_WDTH_L-1:0]        I8d866786bb2dea06f5b30f6ea80cff17;
reg  [MAX_SUM_WDTH_L-1:0]        I01ca9a1d4901ec9b2a64300617ce4cd1;
reg  [MAX_SUM_WDTH_L-1:0]        I2dbead35e15afb9affaa6ad4edd3829e;
reg  [MAX_SUM_WDTH_L-1:0]        I83c57653e24cc09214075b04b06bad83;
reg  [MAX_SUM_WDTH_L-1:0]        I56b9c1f555b24c2dc197168decfdb8d1;
reg  [MAX_SUM_WDTH_L-1:0]        Id5c48111f1b93de2cfe89f92fd182b43;
reg  [MAX_SUM_WDTH_L-1:0]        I32908c3c90ed6488357ce4869e8a1721;
reg  [MAX_SUM_WDTH_L-1:0]        I16b4601f2e07e6cecdb5a030178e75c0;
reg  [MAX_SUM_WDTH_L-1:0]        I0ae08a41ebd0e6b402a4980478087bb5;
reg  [MAX_SUM_WDTH_L-1:0]        Icb57267a66f117943e964dd6420d7a58;
reg  [MAX_SUM_WDTH_L-1:0]        Icfa47fb87b74106cd3814adfce909424;
reg  [MAX_SUM_WDTH_L-1:0]        I63067cef0e1a348a3e6d8cd9bd88b907;
reg  [MAX_SUM_WDTH_L-1:0]        I10aa5ba0f53632578c0e1cefa4bf4fde;
reg  [MAX_SUM_WDTH_L-1:0]        I427c0215d0ac047e8402c20610676752;
reg  [MAX_SUM_WDTH_L-1:0]        Icf4efa87688bd1b80437686eb0126057;
reg  [MAX_SUM_WDTH_L-1:0]        Ic373f785ddd1bf8eccce263df5a82c87;
reg  [MAX_SUM_WDTH_L-1:0]        I56f8e8d2d7052af26528530d389b6dc1;
reg  [MAX_SUM_WDTH_L-1:0]        Ifb145bc18d435fb66779e7415417bc0f;
reg  [MAX_SUM_WDTH_L-1:0]        I62a6e0c9952d6c6e6095e2364df93078;
reg  [MAX_SUM_WDTH_L-1:0]        Id6405c2b2b9aea6bc457f1064d5f3ffa;
reg  [MAX_SUM_WDTH_L-1:0]        I079df9611bd81f672f2ae028bf267995;
reg  [MAX_SUM_WDTH_L-1:0]        I096b226cc511363946a39307a7d97867;
reg  [MAX_SUM_WDTH_L-1:0]        I4cc42c5a75ef339510ee0e86fb44e16a;
reg  [MAX_SUM_WDTH_L-1:0]        I680c01c3327cb9372a42c1ec5b4193e3;
reg  [MAX_SUM_WDTH_L-1:0]        I83451a072082194ecb3f9419edd728b3;
reg  [MAX_SUM_WDTH_L-1:0]        I52ad85b6a1c822ca8c2459bde8fbd510;
reg  [MAX_SUM_WDTH_L-1:0]        I1c44d2ef638825862061a8ee1a0a2f95;
reg  [MAX_SUM_WDTH_L-1:0]        I8fa1fd425809cc39cd8e2785773c1d7a;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa22335f04d35680eb8cfec8f862f357;
reg  [MAX_SUM_WDTH_L-1:0]        I6aff673c27811b81530453906312aa9c;
reg  [MAX_SUM_WDTH_L-1:0]        If674ac0540f457a21235664c213d4923;
reg  [MAX_SUM_WDTH_L-1:0]        Iac223ac498bdcf2cb2514582aeaf76f3;
reg  [MAX_SUM_WDTH_L-1:0]        I7f40931ab78ededfcb52ccaac9b81282;
reg  [MAX_SUM_WDTH_L-1:0]        Iab7c8dad0ca20eb0988fbd99f25591a8;
reg  [MAX_SUM_WDTH_L-1:0]        I3cb5f890a5bd3daaae34c8dfb6ecfc49;
reg  [MAX_SUM_WDTH_L-1:0]        Id80e145586d7e539a6514dd67ebabf6a;
reg  [MAX_SUM_WDTH_L-1:0]        I01e09bc554768f30dc490041d19b4da2;
reg  [MAX_SUM_WDTH_L-1:0]        I0196f7df6f834ae20c4fdd127e66104d;
reg  [MAX_SUM_WDTH_L-1:0]        I4669c4f256c123a0fcceb55c1e72193a;
reg  [MAX_SUM_WDTH_L-1:0]        I4a02ffa2a79df824f406909aa189a404;
reg  [MAX_SUM_WDTH_L-1:0]        I3117e5029119e70846dff61d746699e7;
reg  [MAX_SUM_WDTH_L-1:0]        I1e4e705b3bda1451fc384cd934c0bb52;
reg  [MAX_SUM_WDTH_L-1:0]        Ib5bea8e0072de3de2c8431ea6a35dd51;
reg  [MAX_SUM_WDTH_L-1:0]        I7d9d94022ea95ea01cddc237f3df8cb8;
reg  [MAX_SUM_WDTH_L-1:0]        I3f0f9aab07427fa81fc3096c6b6d3d6d;
reg  [MAX_SUM_WDTH_L-1:0]        I12a7983041f9c298d533bad58f41d24b;
reg  [MAX_SUM_WDTH_L-1:0]        I78503880e5c96ec0a03c75266b1226e8;
reg  [MAX_SUM_WDTH_L-1:0]        I8adeae445b33f634977957bb1a2259aa;
reg  [MAX_SUM_WDTH_L-1:0]        I73bd13f381d15e0b0198b60cee44bb42;
reg  [MAX_SUM_WDTH_L-1:0]        Ic8b651c2b043a4a6e4cd259774322230;
reg  [MAX_SUM_WDTH_L-1:0]        I76979d7df582f9306e796a03cb540963;
reg  [MAX_SUM_WDTH_L-1:0]        If61d4585986757a525c54589ec93d8c6;
reg  [MAX_SUM_WDTH_L-1:0]        I1bc5766a4a3cc2b468ab8ef62eab691c;
reg  [MAX_SUM_WDTH_L-1:0]        I21585169e5fceda643bd03fddf8153be;
reg  [MAX_SUM_WDTH_L-1:0]        Idb2990946f60939136b3bfddbc7b1671;
reg  [MAX_SUM_WDTH_L-1:0]        Icfbf703890f684bfc96decc429deaa04;
reg  [MAX_SUM_WDTH_L-1:0]        Id5bb42639a1c1c1d67df1c89a14a2bfc;
reg  [MAX_SUM_WDTH_L-1:0]        I55b8ef91d667c1c1d9e58dbc86a2288a;
reg  [MAX_SUM_WDTH_L-1:0]        I17ff683da41b469c8c8b82ee32a7378a;
reg  [MAX_SUM_WDTH_L-1:0]        I51f10296c38872338ec7df35ccd520d8;
reg  [MAX_SUM_WDTH_L-1:0]        Ia59ff33765ddf4aeb17f90a70c01d76c;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf97abffb1ec40f2f0e099a814e04ab2;
reg  [MAX_SUM_WDTH_L-1:0]        I3efc3271e18a1e350473dcf3375088aa;
reg  [MAX_SUM_WDTH_L-1:0]        I1efd1220ea9100f2fb4f169ceaf462a5;
reg  [MAX_SUM_WDTH_L-1:0]        I9af399f27c8e2b62b7f3fc6481ef9318;
reg  [MAX_SUM_WDTH_L-1:0]        I171bb4ee9be2f92e4d82997108572426;
reg  [MAX_SUM_WDTH_L-1:0]        Ib13cd76c20fcaf95f26f4914380c4fcf;
reg  [MAX_SUM_WDTH_L-1:0]        Iafb219f1c8c6883e01fbfb4c887c8d6a;
reg  [MAX_SUM_WDTH_L-1:0]        I94fc9b0bdd2b0a89a9f6351f1fdd4ff5;
reg  [MAX_SUM_WDTH_L-1:0]        Ia9ceb45f33402293c162cef4037ba007;
reg  [MAX_SUM_WDTH_L-1:0]        I0fa4e12e62e8a30b3b8045143b344b4f;
reg  [MAX_SUM_WDTH_L-1:0]        Icec1c637d24ca277bb2e488257e92a40;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9aca08b988fad20904545fe070defd5;
reg  [MAX_SUM_WDTH_L-1:0]        Ie82304b2c8583f967649475e309e68fa;
reg  [MAX_SUM_WDTH_L-1:0]        I60da0fb8a2c0669d5f9037ae99b23565;
reg  [MAX_SUM_WDTH_L-1:0]        Id8c19a3547c17ed513d2d857adc66885;
reg  [MAX_SUM_WDTH_L-1:0]        Id74984743844e9495ea0f528a391f4b8;
reg  [MAX_SUM_WDTH_L-1:0]        I9edcdd5b927b3f6b3a4c7cacebeb4a82;
reg  [MAX_SUM_WDTH_L-1:0]        Ic89597a95f50382cd3a2730896735d55;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb7d203dfc75bf6211b09ab94877f93d;
reg  [MAX_SUM_WDTH_L-1:0]        Id2f2e6837c83973cb2173454433acb88;
reg  [MAX_SUM_WDTH_L-1:0]        I1259d5918f8d65b4b22ccfef22fe3afa;
reg  [MAX_SUM_WDTH_L-1:0]        Ib84e8c6e7fd9d7762e6e7e508d5ee40a;
reg  [MAX_SUM_WDTH_L-1:0]        Ia032017912715abde99ffdf5ba732c5f;
reg  [MAX_SUM_WDTH_L-1:0]        I55c310bfefb635448ef9c25c5d15987e;
reg  [MAX_SUM_WDTH_L-1:0]        I92c0f229cf7fdb2cc0fe4d84f4d9b11d;
reg  [MAX_SUM_WDTH_L-1:0]        I5570eb486d238fd96f9a59b174f5a22a;
reg  [MAX_SUM_WDTH_L-1:0]        If6f01d24acf4a8b38bdbb1b366cd9a47;
reg  [MAX_SUM_WDTH_L-1:0]        Iff29fff36064aa4f9d339d4c62956e61;
reg  [MAX_SUM_WDTH_L-1:0]        I818d7cae6f1b80ac452dbfc073ccfe7a;
reg  [MAX_SUM_WDTH_L-1:0]        I77ecfe991c6ec778495d7d5e5e442eca;
reg  [MAX_SUM_WDTH_L-1:0]        Ie7c6a56e8b6f7756bb5a24bdfd6a855e;
reg  [MAX_SUM_WDTH_L-1:0]        I9f9bc8eb8b2978a3dc529c34516fdf75;
reg  [MAX_SUM_WDTH_L-1:0]        Ie3c0e5a4b00a92357a5d37e527d59b61;
reg  [MAX_SUM_WDTH_L-1:0]        I9b9a9486420e7d4aa105c48dd50aa74d;
reg  [MAX_SUM_WDTH_L-1:0]        Id12199a504f7aa298fffaaedd1aacc99;
reg  [MAX_SUM_WDTH_L-1:0]        I813691fd8ea36626d32c8d2562163f32;
reg  [MAX_SUM_WDTH_L-1:0]        I5fd3aaddc3eb8afeb82768b45e2d53d7;
reg  [MAX_SUM_WDTH_L-1:0]        I1ac281eab6c7459e835fe992142b7857;
reg  [MAX_SUM_WDTH_L-1:0]        I49e5078c9161e8bee00fb76bc00b5288;
reg  [MAX_SUM_WDTH_L-1:0]        Ia697adf14616bf50d6e8178596b9fa7e;
reg  [MAX_SUM_WDTH_L-1:0]        Iff3128a26dabe63b015dc6afc98a85a9;
reg  [MAX_SUM_WDTH_L-1:0]        Ifc04708ee5a7cc2b3f1850db778fa42e;
reg  [MAX_SUM_WDTH_L-1:0]        Ia405859c9dff67905b2e91bcbc06259e;
reg  [MAX_SUM_WDTH_L-1:0]        I2fec8f62b28575e8f3af756db66fa232;
reg  [MAX_SUM_WDTH_L-1:0]        I98e97c02477032ead66dc50f3f274e5a;
reg  [MAX_SUM_WDTH_L-1:0]        I9f2dc5add3a4d1e6eb3116c741cd2f82;
reg  [MAX_SUM_WDTH_L-1:0]        Ie122f7d8a48d7ad29d998b6a14b8e70f;
reg  [MAX_SUM_WDTH_L-1:0]        Ib5576c996062391f44066d893dd5cb91;
reg  [MAX_SUM_WDTH_L-1:0]        If931597aab866a74c3a3ffb1cd429583;
reg  [MAX_SUM_WDTH_L-1:0]        I79878bd69ed53785b8a5f025a2a00a4f;
reg  [MAX_SUM_WDTH_L-1:0]        Iefb0a20652954fc2002154ea874c120a;
reg  [MAX_SUM_WDTH_L-1:0]        I646ca66e4e9f24b4fb75b38bf293b4cc;
reg  [MAX_SUM_WDTH_L-1:0]        I051f0d4c44123e3637b84a32c9a00a75;
reg  [MAX_SUM_WDTH_L-1:0]        I1876f9ec3f6f637ee40cdad7cc347f6f;
reg  [MAX_SUM_WDTH_L-1:0]        Ic3d6b8dbec6cf92a9b6a17fb2f75dcd4;
reg  [MAX_SUM_WDTH_L-1:0]        I7d89f1db7b1015d34363ad781374de58;
reg  [MAX_SUM_WDTH_L-1:0]        Ife217ec4da1f1477bce034cb3545160f;
reg  [MAX_SUM_WDTH_L-1:0]        Idc5e5e98508c94b87a760f8eb36fad41;
reg  [MAX_SUM_WDTH_L-1:0]        I9e72b0c823f297535f13a1b3072c2776;
reg  [MAX_SUM_WDTH_L-1:0]        Ia81da7c58d6636ab70e0cf3e263a12c0;
reg  [MAX_SUM_WDTH_L-1:0]        Ibfc69ef08382c79e30cfafd89bfeff69;
reg  [MAX_SUM_WDTH_L-1:0]        I2d2afa9165b7121dc8289e9e6cdab5de;
reg  [MAX_SUM_WDTH_L-1:0]        I065052693fd8ca87614feb60f7ef37c3;
reg  [MAX_SUM_WDTH_L-1:0]        I13344a81551374f665cbc17c7e94296a;
reg  [MAX_SUM_WDTH_L-1:0]        If5a1d2de0715fa87d191ee5f48171676;
reg  [MAX_SUM_WDTH_L-1:0]        I02b256f74ee86b42ff1eba5e3d242737;
reg  [MAX_SUM_WDTH_L-1:0]        Ic113fc051eefaef846f440e98f2f8913;
reg  [MAX_SUM_WDTH_L-1:0]        Iabeab9bdd0bd82dd145218b563b5dac1;
reg  [MAX_SUM_WDTH_L-1:0]        If9ce0a09e3a4e816dda002a24319ac0b;
reg  [MAX_SUM_WDTH_L-1:0]        Ib5a7d72c36e41754033a64fbe0718784;
reg  [MAX_SUM_WDTH_L-1:0]        I41df12c7dee8526abf92b8e98965fa06;
reg  [MAX_SUM_WDTH_L-1:0]        I83dfbd224e7465a6fd769e407182829a;
reg  [MAX_SUM_WDTH_L-1:0]        Ie57bba5092ec318456365b81b36aaa65;
reg  [MAX_SUM_WDTH_L-1:0]        Ibcf043d24474ab8c1002d15fde2d7da2;
reg  [MAX_SUM_WDTH_L-1:0]        I2e3385871c6ed8cf9519f273c8a19fda;
reg  [MAX_SUM_WDTH_L-1:0]        I664917b9f44515bf556d69ade4ca408c;
reg  [MAX_SUM_WDTH_L-1:0]        I28deacdec0fbd0bce49b654c2620ac38;
reg  [MAX_SUM_WDTH_L-1:0]        Ibdfc4852c620f573f929584e6b816f35;
reg  [MAX_SUM_WDTH_L-1:0]        I5a69b2bbb63ab919ea2270503cd326f1;
reg  [MAX_SUM_WDTH_L-1:0]        I2eccd8d60a19481fa595566f51c7aa4e;
reg  [MAX_SUM_WDTH_L-1:0]        I49eb4bba42440657fe04b711eedfa67f;
reg  [MAX_SUM_WDTH_L-1:0]        I9ed8323951af0de78ae89153cbf9e9eb;
reg  [MAX_SUM_WDTH_L-1:0]        I1d00816529836546b514f54b1275d39e;
reg  [MAX_SUM_WDTH_L-1:0]        Icc58b9a24fb9ef7e8fa5f13a2cc0a0cb;
reg  [MAX_SUM_WDTH_L-1:0]        I9339aef608b029175b488e82f5b3f1bb;
reg  [MAX_SUM_WDTH_L-1:0]        Ibd2f24860b701ab46e0c436d774e43f9;
reg  [MAX_SUM_WDTH_L-1:0]        I37fe66ec8927f27f646b304500400ccf;
reg  [MAX_SUM_WDTH_L-1:0]        I4bd6a48f494cf633a857b8ccbd67af68;
reg  [MAX_SUM_WDTH_L-1:0]        Icd7a7566438dc67e77f138ac814844f0;
reg  [MAX_SUM_WDTH_L-1:0]        Ic3d4239413333883dd926c7a42c0a87f;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8298d1ead61bc00eb31599b3087d769;
reg  [MAX_SUM_WDTH_L-1:0]        I23dbe33ce46f94d3dff1e6d391305609;
reg  [MAX_SUM_WDTH_L-1:0]        I138286817f424c76e8a4f30540b0530b;
reg  [MAX_SUM_WDTH_L-1:0]        I30c645a78b900306864a1ab23e923bde;
reg  [MAX_SUM_WDTH_L-1:0]        Id88681d0fe3ea62530166938503db05a;
reg  [MAX_SUM_WDTH_L-1:0]        I808008402174fa4edf42783135c0c3a9;
reg  [MAX_SUM_WDTH_L-1:0]        I3ad4d02ea2e52a49b6fa4f1da9b58149;
reg  [MAX_SUM_WDTH_L-1:0]        I39486eecb7bbfecf26573a7a5876feb9;
reg  [MAX_SUM_WDTH_L-1:0]        I21e8ea20029fb2cb62103405b81b21b0;
reg  [MAX_SUM_WDTH_L-1:0]        Id0b67fa451e276889e02779ddb667904;
reg  [MAX_SUM_WDTH_L-1:0]        Ic328d25a58ec4559b753da3bcff938de;
reg  [MAX_SUM_WDTH_L-1:0]        I49c44c2f2522e086c2db8a00647ba35c;
reg  [MAX_SUM_WDTH_L-1:0]        Id4152a04385391294f4b8a18df2cb9ee;
reg  [MAX_SUM_WDTH_L-1:0]        I5b0213a3df61e94fd0b744a8141f7502;
reg  [MAX_SUM_WDTH_L-1:0]        If0ad11ed403cbbed68614b01e2a3793e;
reg  [MAX_SUM_WDTH_L-1:0]        Icfa1170bc73534bee13778bc3b88a2f7;
reg  [MAX_SUM_WDTH_L-1:0]        Ife1bd938a0dd06d8d3cf30ff41a303b2;
reg  [MAX_SUM_WDTH_L-1:0]        I4a09cb1b99b476fa6fae0bc44c41a041;
reg  [MAX_SUM_WDTH_L-1:0]        Ie08cf323944813e4b9e2d59a680ffe8d;
reg  [MAX_SUM_WDTH_L-1:0]        I85fc307fb52d58550eeecd33bc4207a4;
reg  [MAX_SUM_WDTH_L-1:0]        Id00dd13741fe621d0a240bdc92318f55;
reg  [MAX_SUM_WDTH_L-1:0]        Idc8e891fd432df75a4eb133ce35ecec4;
reg  [MAX_SUM_WDTH_L-1:0]        I2a51cada20cbd14f7d5a289599e68b53;
reg  [MAX_SUM_WDTH_L-1:0]        I65a701d1e083e501544bb0fce24f0c4e;
reg  [MAX_SUM_WDTH_L-1:0]        If3020a9109ac83274b5bafac18d176de;
reg  [MAX_SUM_WDTH_L-1:0]        Iaa6bd55038c2ae911e4df08f707c55f5;
reg  [MAX_SUM_WDTH_L-1:0]        Id49065cedf20e13abac8971534bb8b0e;
reg  [MAX_SUM_WDTH_L-1:0]        I0bb64952d77b59803a561e14b950b9b1;
reg  [MAX_SUM_WDTH_L-1:0]        I01e295a6ab88c6f34b44efcc32a23233;
reg  [MAX_SUM_WDTH_L-1:0]        I2acf864d587b7681ca0fb6e2e2bea617;
reg  [MAX_SUM_WDTH_L-1:0]        Idfd0410b37713e8808f8bea81e2af881;
reg  [MAX_SUM_WDTH_L-1:0]        I02861f333b5adfd4962356cdf5a11f23;
reg  [MAX_SUM_WDTH_L-1:0]        I4ddbc3daa65b111cb0d45e13d62cc292;
reg  [MAX_SUM_WDTH_L-1:0]        Id363d158feb8fec19b5f3d73d84f0068;
reg  [MAX_SUM_WDTH_L-1:0]        I8ec9b7a6e65e727abbed336ce240a4cf;
reg  [MAX_SUM_WDTH_L-1:0]        I128fa1e99b7eb9b6905c2cfd26b95ab4;
reg  [MAX_SUM_WDTH_L-1:0]        I93d459b6da42a205c91c48622f0c5032;
reg  [MAX_SUM_WDTH_L-1:0]        I1243cc8d5dddf7dd65b40c0b3b958b9e;
reg  [MAX_SUM_WDTH_L-1:0]        I238df7e09d42bc93a972da349a00f511;
reg  [MAX_SUM_WDTH_L-1:0]        Ic658b2afdc7331653fc84d6372d47418;
reg  [MAX_SUM_WDTH_L-1:0]        If39be111eb101c9c983fe0baa9a1cb18;
reg  [MAX_SUM_WDTH_L-1:0]        I9d19d5b7d8b256c1707de97a4549c458;
reg  [MAX_SUM_WDTH_L-1:0]        I6c2fffe204091f7f64aea16b0ac98769;
reg  [MAX_SUM_WDTH_L-1:0]        Ic4ba4d2e5c12d9f1dd233d64929f1072;
reg  [MAX_SUM_WDTH_L-1:0]        Ia9dec5831998d472d11429e5a7e60ed8;
reg  [MAX_SUM_WDTH_L-1:0]        Ieaaf52c1e663f260292bc1529718d681;
reg  [MAX_SUM_WDTH_L-1:0]        I37061896a09588a73445deed73d3746c;
reg  [MAX_SUM_WDTH_L-1:0]        I02f25b80945b6f58193fb37add3da2d8;
reg  [MAX_SUM_WDTH_L-1:0]        I19045602bb77f12666ebd44f813db2c5;
reg  [MAX_SUM_WDTH_L-1:0]        I4abdc8d5318d2922696a8aaee46ffa59;
reg  [MAX_SUM_WDTH_L-1:0]        Ie139f2048f346d82623c8fc6d40c9acc;
reg  [MAX_SUM_WDTH_L-1:0]        I8d99c96e203fafc81d13ce5aee925d75;
reg  [MAX_SUM_WDTH_L-1:0]        I37b0bdeb3cc54d6a97720c4912c67832;
reg  [MAX_SUM_WDTH_L-1:0]        I08257e9e6c74c60448e22fb9855f0825;
reg  [MAX_SUM_WDTH_L-1:0]        I32188cca2fc715698fc05b0fc6506434;
reg  [MAX_SUM_WDTH_L-1:0]        I88f1cbab9b8fa3802345f745d024931c;
reg  [MAX_SUM_WDTH_L-1:0]        Idf548c0e78bd221bf9f612f27002fae0;
reg  [MAX_SUM_WDTH_L-1:0]        Iedfd2e04f5740d283388639dde3ecdb5;
reg  [MAX_SUM_WDTH_L-1:0]        I7088c83eacff6f1dfb134f79d469c8f1;
reg  [MAX_SUM_WDTH_L-1:0]        I6f8431671331f4ca7ea19656e0677cd4;
reg  [MAX_SUM_WDTH_L-1:0]        I1e31259e267e04920cbbd16bd7aa18bc;
reg  [MAX_SUM_WDTH_L-1:0]        If54d9f8088e67e44cfa3026f5a520fd7;
reg  [MAX_SUM_WDTH_L-1:0]        I6fd2c0746407b23aec5dff1e083f5fca;
reg  [MAX_SUM_WDTH_L-1:0]        Ib2147a19b44d361da628a628fbfaa988;
reg  [MAX_SUM_WDTH_L-1:0]        Ie804d1f4b241a2de3e9d9c7c876d914a;
reg  [MAX_SUM_WDTH_L-1:0]        I6cd1e6db57e06d8f5e60a31f48ae4809;
reg  [MAX_SUM_WDTH_L-1:0]        I3e0e8832d5338423284ac4b2a0c5f3f5;
reg  [MAX_SUM_WDTH_L-1:0]        I6ac006d79e95e222cdc66754b67a08ed;
reg  [MAX_SUM_WDTH_L-1:0]        I29087dda1a527842aeb3d35d66c853cb;
reg  [MAX_SUM_WDTH_L-1:0]        Ia67e5920bbac700dfee52cd96b15963e;
reg  [MAX_SUM_WDTH_L-1:0]        I1f6ecd894d90547f661e7a3888d048bb;
reg  [MAX_SUM_WDTH_L-1:0]        I3112e793c6e79e1f5da2776e69a34e3c;
reg  [MAX_SUM_WDTH_L-1:0]        I79152f32b45ed5b4a5302f6460707b01;
reg  [MAX_SUM_WDTH_L-1:0]        I3d16e7d6b190639b88a217f19ac63233;
reg  [MAX_SUM_WDTH_L-1:0]        Ia1be780c686163cea54b62d6ede72dc6;
reg  [MAX_SUM_WDTH_L-1:0]        Ic398c31a2a6ca89d0236534589a5919b;
reg  [MAX_SUM_WDTH_L-1:0]        Ie91c3202bc957b350d1915000564392f;
reg  [MAX_SUM_WDTH_L-1:0]        I687957f5300b0d4f50d6893cc556bf25;
reg  [MAX_SUM_WDTH_L-1:0]        I7816b368e8e8b8dd69383b2c9327120d;
reg  [MAX_SUM_WDTH_L-1:0]        I5f021f4a664205afbe0761af4c8914f1;
reg  [MAX_SUM_WDTH_L-1:0]        I69728004b59b5206a03a8e2087834f7d;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbe1d623f8f5f3aa7fc70197acc6df5e;
reg  [MAX_SUM_WDTH_L-1:0]        I4cb9f74288811592fd97fdff52bd6fe7;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb471dbccd39d41e951e98348812e343;
reg  [MAX_SUM_WDTH_L-1:0]        I7f37d68f8ddcf8b4d5e99fb51eada873;
reg  [MAX_SUM_WDTH_L-1:0]        I72ded7153883418a712ef967439d2159;
reg  [MAX_SUM_WDTH_L-1:0]        Ie071e08299bff6bbdbe1f84703aaec08;
reg  [MAX_SUM_WDTH_L-1:0]        I1b79aa38a39ccfc839260af89aa78e7a;
reg  [MAX_SUM_WDTH_L-1:0]        I7384296e4190d83fb9d9a92cf965125b;
reg  [MAX_SUM_WDTH_L-1:0]        Ie03034ce6233ca24effe53a2c0c8f6f3;
reg  [MAX_SUM_WDTH_L-1:0]        Ic298f77f42fc1d41cce684790036ecfe;
reg  [MAX_SUM_WDTH_L-1:0]        I805269f95afbeb6b93182f68868d08eb;
reg  [MAX_SUM_WDTH_L-1:0]        I881328804c45b06767af51e11182b27b;
reg  [MAX_SUM_WDTH_L-1:0]        I958993626e6e44e12f7c1e8026914680;
reg  [MAX_SUM_WDTH_L-1:0]        If31528d1fc3a083ebc364e75cdd9c71f;
reg  [MAX_SUM_WDTH_L-1:0]        I4703b8d5a9033027889bfa8685e09e4f;
reg  [MAX_SUM_WDTH_L-1:0]        I22d8e84d2db4b07111b7fdc6eef34cc8;
reg  [MAX_SUM_WDTH_L-1:0]        I8b7c6df3b5ea575caab7820c95974608;
reg  [MAX_SUM_WDTH_L-1:0]        Ia8aa76bccf7eb310a9356e8b7ea1609d;
reg  [MAX_SUM_WDTH_L-1:0]        If9de547bf469b8424f1625e990f72b04;
reg  [MAX_SUM_WDTH_L-1:0]        I27d51b2015ea9af9bc345adabdb07b6f;
reg  [MAX_SUM_WDTH_L-1:0]        I93dddce2a0dc01ecb3039fac5cf04011;
reg  [MAX_SUM_WDTH_L-1:0]        I746da2c1d5a620eb7e749f72f0f04a06;
reg  [MAX_SUM_WDTH_L-1:0]        I1e15f8d6fdb4ac732768d0cf73af829e;
reg  [MAX_SUM_WDTH_L-1:0]        Ib719e667d7ba857f4f7432a245f4a30f;
reg  [MAX_SUM_WDTH_L-1:0]        I4c6eec4a0c46e4f5d7c9734df48a16bb;
reg  [MAX_SUM_WDTH_L-1:0]        I95623ec1fd5516040a9492aae0fc2b70;
reg  [MAX_SUM_WDTH_L-1:0]        I69017b49c11de463fe6d881e5c96a1aa;
reg  [MAX_SUM_WDTH_L-1:0]        I4fb9ed32471aa614ce6923f6a2279b36;
reg  [MAX_SUM_WDTH_L-1:0]        I2f0bc217c8a39d71adc1fc45c10b81c3;
reg  [MAX_SUM_WDTH_L-1:0]        I0f1c6bb577ea2b8b2ab636e64378544b;
reg  [MAX_SUM_WDTH_L-1:0]        I7a248af9d606c566e03977e985c280e0;
reg  [MAX_SUM_WDTH_L-1:0]        I0bf9d47bff47277de1e72518e8d88362;
reg  [MAX_SUM_WDTH_L-1:0]        I24b6f4f68f291dc50caf03dc902282cf;
reg  [MAX_SUM_WDTH_L-1:0]        I79335b28eea15735f760b7a8b803e93a;
reg  [MAX_SUM_WDTH_L-1:0]        I0b14b34b06cfa90539c2abca5639abec;
reg  [MAX_SUM_WDTH_L-1:0]        I26878777354945712f834740b17dabcb;
reg  [MAX_SUM_WDTH_L-1:0]        I6cc5daed4de5950c02c0a57b993e22fc;
reg  [MAX_SUM_WDTH_L-1:0]        I52c382d5b0c4829127c011fae402ce04;
reg  [MAX_SUM_WDTH_L-1:0]        I46ea9871e867034daa2d0501038f15e0;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb8a202599550e87831647a93a14181a;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb79f2ce0b6028ebb638fc6661444cf1;
reg  [MAX_SUM_WDTH_L-1:0]        I0d0c07d65eda2eee01df9c330c0d6f4a;
reg  [MAX_SUM_WDTH_L-1:0]        Ie6940736944bac9be609b8d58b2cb13c;
reg  [MAX_SUM_WDTH_L-1:0]        I472a71363435cb3ec054e00f9123ae64;
reg  [MAX_SUM_WDTH_L-1:0]        I553223e9166dcbddd1a51d0f92d68f28;
reg  [MAX_SUM_WDTH_L-1:0]        I495309d795905a53b0a3d3daa4f1f9d0;
reg  [MAX_SUM_WDTH_L-1:0]        I21d358fd7673c4392f4e4b3d3a858b2c;
reg  [MAX_SUM_WDTH_L-1:0]        Ia1a60175112362f015c5531f7c48b90b;
reg  [MAX_SUM_WDTH_L-1:0]        I5644ece811bddcec04c9e3559c86109d;
reg  [MAX_SUM_WDTH_L-1:0]        I37d2f9d3f05cb90e2d45bd578299885c;
reg  [MAX_SUM_WDTH_L-1:0]        Ie7d10f3c0f8b0add66d2cdd4435ccc88;
reg  [MAX_SUM_WDTH_L-1:0]        I3c37396a1cef2f9e42b8ccc126db6eda;
reg  [MAX_SUM_WDTH_L-1:0]        I2f82390734079b8d289d48a6682cc624;
reg  [MAX_SUM_WDTH_L-1:0]        I9061728c3163ae684e8c5aec3e807868;
reg  [MAX_SUM_WDTH_L-1:0]        I672d7ecc28a788c2602aff76187aa568;
reg  [MAX_SUM_WDTH_L-1:0]        I660b2fe99cd0bcaac34e9540118b54bc;
reg  [MAX_SUM_WDTH_L-1:0]        I6aa263fc2a061d2c4059b08309f860f4;
reg  [MAX_SUM_WDTH_L-1:0]        If3aef2d755013d195fd44f734365d7dc;
reg  [MAX_SUM_WDTH_L-1:0]        I3ad2e0bbff17683824f575deff82c6bc;
reg  [MAX_SUM_WDTH_L-1:0]        I5087dc4b32d29bfd7bad49026fa58a5d;
reg  [MAX_SUM_WDTH_L-1:0]        I8a7d893f3ef6d6a93ba552320d901599;
reg  [MAX_SUM_WDTH_L-1:0]        Ic057537712e09fa794918e5cde87e084;
reg  [MAX_SUM_WDTH_L-1:0]        I0cbab5173052c450504e3a7d15ffda52;
reg  [MAX_SUM_WDTH_L-1:0]        I81ee40feb7abd0fec3faee653f778f5f;
reg  [MAX_SUM_WDTH_L-1:0]        Ia344347a85d4e6afafa2ee3487e65def;
reg  [MAX_SUM_WDTH_L-1:0]        I038fce1597157a3d95bd9579cc2dcbc6;
reg  [MAX_SUM_WDTH_L-1:0]        I546585b819c289d855cd098818792e90;
reg  [MAX_SUM_WDTH_L-1:0]        Ibc3a6609765818327e79519f3e348494;
reg  [MAX_SUM_WDTH_L-1:0]        Id1c71a2a34f9e6239559d28fe2780907;
reg  [MAX_SUM_WDTH_L-1:0]        I1cd6cf5f8119d5e6b4ca40694399b1c2;
reg  [MAX_SUM_WDTH_L-1:0]        I15e2a1b4356785d73e2ab5d51f1f5ec0;
reg  [MAX_SUM_WDTH_L-1:0]        I803aeb29e66384bfc62744a841bcc83e;
reg  [MAX_SUM_WDTH_L-1:0]        Ib6e220dd4f54410239dd0c791d84a700;
reg  [MAX_SUM_WDTH_L-1:0]        I8a009007fec23f4d492b0da1b6b404fa;
reg  [MAX_SUM_WDTH_L-1:0]        I5f89adcb1ba235a74639eca119fb2655;
reg  [MAX_SUM_WDTH_L-1:0]        I8fd2b001ff154e4760ead2df355c80da;
reg  [MAX_SUM_WDTH_L-1:0]        I581569cc2e63bc68a8466b07ca471b25;
reg  [MAX_SUM_WDTH_L-1:0]        Ia9cfdea21a65b0270de42cef7ebbf822;
reg  [MAX_SUM_WDTH_L-1:0]        Id66a233d2e312aff939549dfa96a8cf0;
reg  [MAX_SUM_WDTH_L-1:0]        Ie479c12c25a1964c3804936d45725bdc;
reg  [MAX_SUM_WDTH_L-1:0]        Ie30d8770ab7e6643fcb67463f6999125;
reg  [MAX_SUM_WDTH_L-1:0]        I4a17ff532c9341e80f7ed0626f728054;
reg  [MAX_SUM_WDTH_L-1:0]        I597bc1ec224007a78c25f7eea24c2c3e;
reg  [MAX_SUM_WDTH_L-1:0]        If198ec15fcf66e97e69f88f718979c2b;
reg  [MAX_SUM_WDTH_L-1:0]        I6aa13ef29cf7e86ec83affca4fa11e42;
reg  [MAX_SUM_WDTH_L-1:0]        Ide136b08f4b6211bca8cccf494a0baa5;
reg  [MAX_SUM_WDTH_L-1:0]        Ieeab247764c23256749776b0a164314d;
reg  [MAX_SUM_WDTH_L-1:0]        I210e9ff7f4588185bd712915954543ce;
reg  [MAX_SUM_WDTH_L-1:0]        I59186d5219833d6dd2e813a2910a61f5;
reg  [MAX_SUM_WDTH_L-1:0]        I0c8b2bb61a9c3a67ac7e03e40be2b98e;
reg  [MAX_SUM_WDTH_L-1:0]        Ide24c1f9033e7057262da1bc4762b840;
reg  [MAX_SUM_WDTH_L-1:0]        I4677558b9faf190e7960cfa9b8ee00fd;
reg  [MAX_SUM_WDTH_L-1:0]        Ie38ab94215851e531d2100b6602d5fa5;
reg  [MAX_SUM_WDTH_L-1:0]        I3f5119e8fac99376aa38e4765b8b0f99;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8040301d224f78c1fd18bfe9e29e5ba;
reg  [MAX_SUM_WDTH_L-1:0]        Ied989966cebf0d730633606c5182a249;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8818bc4ca106ae38cacd5c20083aa08;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf08556fc39044222321912e84a4436b;
reg  [MAX_SUM_WDTH_L-1:0]        I985e2740ac0f656da8f9dd973bca99e6;
reg  [MAX_SUM_WDTH_L-1:0]        I73012d2d9f6f237bc50bbffc199e012b;
reg  [MAX_SUM_WDTH_L-1:0]        Iefd0d59e58623b14437b17297fdbf4ff;
reg  [MAX_SUM_WDTH_L-1:0]        I68d2443e98f2fd3fa3baf96f98e1f4bc;
reg  [MAX_SUM_WDTH_L-1:0]        Ia2d1b6833cd8ed02f05281e508e4d716;
reg  [MAX_SUM_WDTH_L-1:0]        I512e2251bef73108eb0f3e01e79ca3fb;
reg  [MAX_SUM_WDTH_L-1:0]        I9bf64811d14ca8b4c633342ad22669a3;
reg  [MAX_SUM_WDTH_L-1:0]        I45a910acd40d5b9417bdfdc50cddf241;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbcf5c5f4528b03508b506c43e4511c4;
reg  [MAX_SUM_WDTH_L-1:0]        I2b8b54048e164ef2f1c072517fdfe400;
reg  [MAX_SUM_WDTH_L-1:0]        Ia48d8883fe4f685477da6b4b05ecd387;
reg  [MAX_SUM_WDTH_L-1:0]        I276395da1f3f1ae246b082408be2cb80;
reg  [MAX_SUM_WDTH_L-1:0]        I4d0e2e01d9abf9ce839fe650abfaaddd;
reg  [MAX_SUM_WDTH_L-1:0]        I7e4e7909094f762c54137cbee99255e5;
reg  [MAX_SUM_WDTH_L-1:0]        I761255e100d161b25645ca3a5187e82a;
reg  [MAX_SUM_WDTH_L-1:0]        Icc2ce1fa3cde69256378ec3f4a07b0fc;
reg  [MAX_SUM_WDTH_L-1:0]        Idd99afa80ca23644675d3edd60e74fe4;
reg  [MAX_SUM_WDTH_L-1:0]        I486bcb4fb0af80c98c2ea21ac64f7a90;
reg  [MAX_SUM_WDTH_L-1:0]        I759cca2c0003fc2c2af7709c5ebc59f7;
reg  [MAX_SUM_WDTH_L-1:0]        I1d5ce9f132cd1f46e96b511c77234e21;
reg  [MAX_SUM_WDTH_L-1:0]        I032e26ea05e88c6d325a810b67e82306;
reg  [MAX_SUM_WDTH_L-1:0]        I0f72df5225a1fec2f276fd3c9138e8c3;
reg  [MAX_SUM_WDTH_L-1:0]        I0d18cf087b2335f1b9e1a621acd5379f;
reg  [MAX_SUM_WDTH_L-1:0]        I7684fc23c57105e856050a45640f2bfd;
reg  [MAX_SUM_WDTH_L-1:0]        If778767ab80e59e940deeaa8a0dac99a;
reg  [MAX_SUM_WDTH_L-1:0]        Idaf86833beb8c334f99291db9302ed29;
reg  [MAX_SUM_WDTH_L-1:0]        I6610e8d41cea10498d95850440ce388b;
reg  [MAX_SUM_WDTH_L-1:0]        Ibc653e701eb995e828c8180efaa122c9;
reg  [MAX_SUM_WDTH_L-1:0]        I21d36c49c9c766139b4b01df7c00a8f3;
reg  [MAX_SUM_WDTH_L-1:0]        I0e4ffded936d7ccfc32b410aec617df8;
reg  [MAX_SUM_WDTH_L-1:0]        I1a5745021323efb5327d0b893962e852;
reg  [MAX_SUM_WDTH_L-1:0]        I65547afdcd7fedb7b44bd51358eec4d2;
reg  [MAX_SUM_WDTH_L-1:0]        Iada3eb71e94ff6a6f4e5c702e83036ed;
reg  [MAX_SUM_WDTH_L-1:0]        I077404a911da16d707a326f18717dc7a;
reg  [MAX_SUM_WDTH_L-1:0]        I6da1e92759c96aab8b9207a9acb244ab;
reg  [MAX_SUM_WDTH_L-1:0]        If7110182720ffa279b1cec1305cf9889;
reg  [MAX_SUM_WDTH_L-1:0]        If0e20ea1696ff84329b9928d7f9e3381;
reg  [MAX_SUM_WDTH_L-1:0]        I4e69ae6e73a856d4e26203fb9acf3565;
reg  [MAX_SUM_WDTH_L-1:0]        I64c939aa568669b4567c21be09ad0e94;
reg  [MAX_SUM_WDTH_L-1:0]        Ia88eb16f68265e322509d541eb457993;
reg  [MAX_SUM_WDTH_L-1:0]        I916f75e5a3858a420ab5cd4c43b13921;
reg  [MAX_SUM_WDTH_L-1:0]        Id076f99460a8f73a9fd43467216e8f8e;
reg  [MAX_SUM_WDTH_L-1:0]        Ib4d7aeb8544fbdc36575a55b9f67f2dc;
reg  [MAX_SUM_WDTH_L-1:0]        If65d2514892fb7ee64fa4dc37fc0fed3;
reg  [MAX_SUM_WDTH_L-1:0]        Ibef07e48768252e9b41baf067bb1ff5d;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8fb61fa9cb8e92bc57c53a567891895;
reg  [MAX_SUM_WDTH_L-1:0]        Id8f5f32cd0757b4d6861d17fcbd6e8d0;
reg  [MAX_SUM_WDTH_L-1:0]        I8be241f29e7eb258e9b3501430820b0d;
reg  [MAX_SUM_WDTH_L-1:0]        Ica8a188ea43e2f28e70b8ea4e2431dc3;
reg  [MAX_SUM_WDTH_L-1:0]        I83ceb726e57d52698b57dc39ce585897;
reg  [MAX_SUM_WDTH_L-1:0]        Ic88e7e05d83ff800b4a941ae4b424557;
reg  [MAX_SUM_WDTH_L-1:0]        I7de81aaac1e5776dfb60eed2d12d4f6d;
reg  [MAX_SUM_WDTH_L-1:0]        I37058036bd9f4331387ee4a9348541e2;
reg  [MAX_SUM_WDTH_L-1:0]        I570f85838c418d8501c8ccdc38a53f00;
reg  [MAX_SUM_WDTH_L-1:0]        I4aa6f0c0f5163b944f11328888af73e0;
reg  [MAX_SUM_WDTH_L-1:0]        Ic7fc1f38ad4e9b2cb472ae75bc3c100c;
reg  [MAX_SUM_WDTH_L-1:0]        Ibace8d2fba25834c83b1e57195c81086;
reg  [MAX_SUM_WDTH_L-1:0]        Iefc1488e3eb60b99ae08d904a15c5242;



assign I97afe24956b7f87cd431f048202bab67 =  ~I5deafec6e5f32da1bcf8f7018cf794d8+ 1'b1 ;
assign I117235e3ac8e68e4c1ab34db1612aba0 =  ~I35b3fb2670f3a60d165c1fd10f02c00c+ 1'b1 ;
assign Ifd700cc9d18f99b63f1947f3ae631976 =  ~I68925439e233444a4da44871f31de94a+ 1'b1 ;
assign Ifffbe3d1007fb07a20d3b37902b3ec95 =  ~I3108702b5ca506422c1ba6174619f193+ 1'b1 ;
assign If5443777169422ea6e1e3f709b970e05 =  ~Icc8e8f6446ac64350a05f5e1e0541bb9+ 1'b1 ;
assign Ifaf9fc93e4609d818aa46751754c17f1 =  ~Iadebaf3f6cca1ba78feab50ce70c8aef+ 1'b1 ;
assign I419caf964986c655df84d043badc37c9 =  ~I8681cf376dbeceab29279a7637249e7d+ 1'b1 ;
assign I3095214ac0e6c1323e75ee4ec85e6821 =  ~Ie850a07565bed90389bb125ddcd39658+ 1'b1 ;
assign Ided9739bf63937933250a6d0c37535f9 =  ~I97b77743c2311ec629ea24c933b60053+ 1'b1 ;
assign Id0f139b9f3848b45554ac8429230eea2 =  ~I07a0a8d41ed8176e92380f2c89c2afdd+ 1'b1 ;
assign Id9feed58cf9565255abfd0bf7e3ec068 =  ~I021842328f948a94159b32903c8bcb68+ 1'b1 ;
assign I30a3be3b5f6ad1880a917eb35659a1bf =  ~Icaf3bd685005a05c8fb334266ea4e4b9+ 1'b1 ;
assign Ie8148d9aa962a733eb65877b902a187d =  ~I92d9e1d7dcf45a4d738c546e959687c3+ 1'b1 ;
assign I69e98cf3e679183aef6005bb582b18dc =  ~I39ca3a8ca714a9726114326ae6bfab0a+ 1'b1 ;
assign I7f42a504fc61c9548acebdd8b1858eaa =  ~Ie9ae20ed5b2a0cad2c37c5bb2ea05ff4+ 1'b1 ;
assign I08b1b4639b5a9ca509b943b977f6d4bb =  ~I8f131eb6138c23fdcb35195703131e64+ 1'b1 ;
assign I8d7296627d886566783e79c01b9fa423 =  ~Iff77e08da4bcbb85b95fa277b69653a9+ 1'b1 ;
assign I4fc4c97229a8b1f631a3b505941159e4 =  ~I703e0a4879a39b3b8b0a49de86ca4ff4+ 1'b1 ;
assign Ib9b16bf51891c328dba2699eb9bcef95 =  ~I3da217f6f2d0f515bb9036673d753a88+ 1'b1 ;
assign I6c30501ec81fce286817788d614a7824 =  ~Ifcc06d5a010e01a781ae8a9e9e2b31a0+ 1'b1 ;
assign Ia4d4f37baec48121a88808075dd655ef =  ~I42fd611fec087113ba6e35f281bced9c+ 1'b1 ;
assign I385495ea2bf6442a95ab7561456254ac =  ~I5bb626e7347bb9ae4219cc72244b38f8+ 1'b1 ;
assign I5128e03d383c226befa6f7422f3a6f04 =  ~I47e2dac0068652338f94ddffd2dbe88a+ 1'b1 ;
assign Ib208908bab4c20713cd17e20139c8db3 =  ~I59a3f06de2984078a4d4c430a2980fe3+ 1'b1 ;
assign Id939992b99a11c09f4688c10ca1a34d1 =  ~I857b7fd58279b1063a06a4f33b880ba6+ 1'b1 ;
assign I823453ccb90d5b2b2d9dfc6e8358224d =  ~I3901bbda029cd0a41640001c1efd400f+ 1'b1 ;
assign I279c5c00b92eb1b872b5afa168b0306e =  ~Ifceeccf10f1d85a32f70c04654a1a1b4+ 1'b1 ;
assign I66f25b1c3c0eb226295179adcca2c3d2 =  ~I2d810c1d1304658edff74921e8d0f388+ 1'b1 ;
assign I3068627e91b667d14cd3e55a9371931a =  ~I575b0201be445388607ab83465eab8d6+ 1'b1 ;
assign I44c4e0a2d8a7289f8660b81a9ecfa19b =  ~I7928c5ce0f821df1cb6271d15e19fa22+ 1'b1 ;
assign Ibe868e258dc87f0dd1460ba6b8354671 =  ~I12695a21c942d02a432cf6382d7d7452+ 1'b1 ;
assign Idc3083c3021200345e3edd35a9d4725a =  ~I00d03f0f71b008dad8035bbf251f41bf+ 1'b1 ;
assign I320d4f19a5b18c23ff407508d47caa77 =  ~I41afedcbc0f492e3243436cbefdaf609+ 1'b1 ;
assign I16becf3c92615d98d5ec51ee9641cc0a =  ~I638c4c2708e437a050ed7cbbac516a59+ 1'b1 ;
assign Ifbfacc3b3a0128119943bcbf80176612 =  ~I6877d3306b1f08c236b5d1b59f0de259+ 1'b1 ;
assign I6b4f670c9e8e25984e8891f2440322ab =  ~Ib3e66aa460f39d32110ea6f115785b3d+ 1'b1 ;
assign I19bf0990a30c72421f231772b8627e8e =  ~I5e603e8392a5322951b3225b65b19446+ 1'b1 ;
assign I3ec3eb096ebe3ee8a47e1cba6487b997 =  ~If5da7fa1a615e1122445460e33487772+ 1'b1 ;
assign I7379ef16405c461ac44b66c4315df831 =  ~Ic4153dafafaf7d047478c5d81109437f+ 1'b1 ;
assign I79db45b23d21d533a1f9a6e8f94d403d =  ~I7b5476007f04e81afc0125e6a8930303+ 1'b1 ;
assign I0979534730cc2b53547d413dbb6b75f4 =  ~I3521a18022925249caddb8e37d2c1262+ 1'b1 ;
assign I5aa2f9c0667d1a6e871efbd4d2bad3a8 =  ~Ifd0f52d4f814e2bb4c3bd34c1e09bda7+ 1'b1 ;
assign Iadb28dc990ccf2dd3099544de16b8f16 =  ~I8945f6d420c8b373225451defcd2c805+ 1'b1 ;
assign I1f71aebf698788d6ada66891e9ea756f =  ~Ieec6cb6518cc0d9300de0c4f2d32487d+ 1'b1 ;
assign Ib234e9cf7e7616a1ebc6ab99df2a7ccb =  ~Ic62eb7e90d703ef994e68587345a4293+ 1'b1 ;
assign I297d1edcc583ea4d69da780150f0620c =  ~Id3efd8419da986aa89b8ad8e75848cfa+ 1'b1 ;
assign Ib0a717cbb4fe38a3fc85520ca0826fd9 =  ~I40803f10b7c4dc9ae4969739349b0265+ 1'b1 ;
assign I037ecd5945b1f1280b4469d73fe1c7ff =  ~I7d961743fdeaf1e72e4b25c12a1d4c46+ 1'b1 ;
assign I367ff6b11b884e02a3065fc7fe811e15 =  ~Ifea156f33eb61fece272efe379327f6e+ 1'b1 ;
assign I6fab19692b512166fe9c74b5e987788d =  ~Ifc99169b3399f3d14121c1a9bce3fc21+ 1'b1 ;
assign I04dd73af505f618ccdb209b3cf97ceec =  ~I6536144383cbda6f3b3c564391866906+ 1'b1 ;
assign If8c559905d4120488d431719c4e8ce24 =  ~Ic21bf9a8a4cd85ec123d7fe142ed49c0+ 1'b1 ;
assign I20ed4f6f14e20ce3f0e106d1b7782fcd =  ~I1f31fe6a0ca8510bcadbc2069403150b+ 1'b1 ;
assign Ib10626ffa126188c5bf1fc8399107b26 =  ~I0e40933d00f4a7d9b53b2764aa0da700+ 1'b1 ;
assign I29007c52357ac7afbda39d72a5bb60af =  ~Ic41a6e00bc84bfc1b8194d15bb899c93+ 1'b1 ;
assign I66d367c046611f145e607a90911cf499 =  ~I2832571f2b0a7fbb41d2e8ca7f64e003+ 1'b1 ;
assign I9c4c2556f6170a8df61d909855a846ed =  ~I9593c853e41952e408a809cb24efa4fd+ 1'b1 ;
assign I6fadc3e8d995bb4317bf7b4377c3c2c5 =  ~I6edffbf4136e193dca0fcec3a74e8e9c+ 1'b1 ;
assign I99b20e911c189e0616f02376ab736e91 =  ~Ibaed50cc2e36ae58945887d11a6ec9e4+ 1'b1 ;
assign I5793c12f5dbdd8245dbb202d550ca960 =  ~Ie4570cac44f59e6ff46f73a703026479+ 1'b1 ;
assign Id0660e9637cad1ce1a73d37188060154 =  ~Ibaa136d37936687e9dbe4222749d19c3+ 1'b1 ;
assign If5a7af7ca023e1393526e888f4220a44 =  ~If85de3225f45478827b43b89089cd29e+ 1'b1 ;
assign Id043eb50634e803e53adc1168379a5d0 =  ~I0344b86a6e9c036e103a9c1f3651175f+ 1'b1 ;
assign I1f866dd0b129267550aea1a267d9c91e =  ~I5463d13575e0b9fb8a0f6cc8b35d0ce9+ 1'b1 ;
assign I8c4da05c08210fe33139c3d3e5d75d58 =  ~I8a3c63ef122001a29e5abe93c4e1a48f+ 1'b1 ;
assign Ib41f7b823681fdd084b6d8436a407aa8 =  ~I6a79108484fcb192f6d93bfb98e271c4+ 1'b1 ;
assign Ic5b50a785b7acac7e3be4095aa92e50a =  ~I9001e95b71457a2bd09a9846af370b16+ 1'b1 ;
assign I3ffbe03796b66d00d47fd918be60ab89 =  ~I51620de618db6327358a5cac97e1e97f+ 1'b1 ;
assign Ifc92a916da938ef6164db250be635f88 =  ~Ib9c58818059af5c5a03e77a5dcef4654+ 1'b1 ;
assign I8ccd42508ce7d5bd897c2cf0c54caeb3 =  ~I8081c71aa01a8d575bfea6ea7f2f595f+ 1'b1 ;
assign I4920e7e82749cc036b58a7cd0a03e327 =  ~Iad999607ad8d7da0f3b341f83ea030a6+ 1'b1 ;
assign Ie1040b2aa91f272e4449c4b5f9f8f575 =  ~Ie7291c914d2cb66f547b0a7717f71311+ 1'b1 ;
assign I65968fb0f63d52ad96cd8fa270126a1b =  ~Ic01018a5f1bc392bbd267016f6612a83+ 1'b1 ;
assign I839ac8ee59f51d4c3de92ba5cb26e788 =  ~Ib11dff839e7e532657b32f29fd9b1651+ 1'b1 ;
assign I33cd95f1919318a0f3df5df7310d64c6 =  ~I251d7ea16dd5407d22a6846ddcfe12d8+ 1'b1 ;
assign I4933e8d16fba26cd797b25a9ac2a2de8 =  ~I773797f81f73b9b6e844441142a1bb48+ 1'b1 ;
assign I218f7578eb748e31d0002052f30c5842 =  ~I853ecadf30fc10a13dd1ffb1f2dfb5d6+ 1'b1 ;
assign I2a808d1c42ad758ae3baaaee8129dfb2 =  ~Ibb8b3c91e1d3b890cfe58f32f8ec3ae3+ 1'b1 ;
assign I4e851fd3c114af87f5e8c68c02594e3a =  ~I3485d69de942d64e56925da522175b51+ 1'b1 ;
assign I0da40f88adc46e90f616acdcdb8e0e2c =  ~Iae42f12bc0475c8b58341d80027a57cb+ 1'b1 ;
assign I0dee7767e472a5fd71250ae6c57cc8b5 =  ~I22fe2af25463f87ee7315a9aac32854e+ 1'b1 ;
assign I9f40be7552b3dd625e5bce0befc5a548 =  ~Idf44ad78c338c39699721ce511691dfd+ 1'b1 ;
assign I8fdf98ffd757c8845ed6ffa4ddd1a16b =  ~I984a657f9265d41318c0290e249e9712+ 1'b1 ;
assign I8103b777314a4fa471e0898fde9cde08 =  ~I915fccfb1d1ada9aa7c8e24c2eebd04c+ 1'b1 ;
assign If6c3ee8e0d7dea58043d5be0f4630873 =  ~I2bdf58ecd0974720631be830efb48dc8+ 1'b1 ;
assign I711a5171f591f472cdbfc9a0f5e1aa17 =  ~Ibaedf6246fa43acc8accb5a24d49cc2f+ 1'b1 ;
assign Ic30bc38184dfbbd694af52640692709d =  ~I904d13524dcdf55478a5266d50e53ff7+ 1'b1 ;
assign I422f6fd1d273a3834d04b04ab8e2812d =  ~I22d8e5d57c1bc082169437a654d22bba+ 1'b1 ;
assign Ia0fdc60b90ad18b6585ec1ad4e89e80b =  ~I719cdaa2a2e61a0df7f1fd5efe517426+ 1'b1 ;
assign I7809fe7a30d041a7e569ffe890242df8 =  ~I8e92a61eb73c41680652936cfcc614ff+ 1'b1 ;
assign I672b14ec1b3c4797545f266727505a85 =  ~I7ad5af8319f6da469858300f0777b580+ 1'b1 ;
assign If9620d20ebaae6245a2c386d9bf5fdb1 =  ~I32be72eaf04e79120a57ea94296a4e56+ 1'b1 ;
assign Ic74e22bffd88f32eefe499cde0fafa8a =  ~Ie756f6a87d85adb40479ce7cf3545556+ 1'b1 ;
assign I76d38ce67387bd76ab45c9cba7d18b31 =  ~I8794c6ce0a3f2e6697372e2c911ba420+ 1'b1 ;
assign I44413c6f6f6493f8a86abf6eb32604f6 =  ~Ic82b1a29b5e63bcc3686a0d4bf1f5c24+ 1'b1 ;
assign I67f632fca617fe06565ddcaaee8fa8b8 =  ~I253ef976058080beab79646af18e2d5b+ 1'b1 ;
assign I3fd38a71ce6aa3db1d7a5a9f8a991e12 =  ~I930dd54c36540d75dc870eef89960163+ 1'b1 ;
assign I63e5718bf7d8771ef90b91be73d73264 =  ~Iaf7554cd4e8b5ea6155ec61a8d589b86+ 1'b1 ;
assign Ie385e1aeb2b0dcf6d2454be3d7708b27 =  ~I50907c7d1efa0038d81efed82b192891+ 1'b1 ;
assign Ib2d1b7e105b25b492b45da72536d7578 =  ~If3e9486d2960d164d94641d4f1917416+ 1'b1 ;
assign I588abf5ef4c583f0fec422736a0ce6a0 =  ~I2bec61db45dd79b98d6ebff6c5a4899e+ 1'b1 ;
assign I58bb95c56c7be17c263a2161210d7d8d =  ~I7f31647f3ea6ce7bbd211c25cf4828fb+ 1'b1 ;
assign Ifaf0e1f21b3bd7393c475b5126540a72 =  ~Ice65387e606faf9c7b884475b489abba+ 1'b1 ;
assign I7027db9e0450724a6d417d708f1043f2 =  ~I63f914927dcf49552e9f3fe0180a30e8+ 1'b1 ;
assign Iebcb7206d8860b5094459c5d10b4efed =  ~I742ff5725e3a18acd03454cf9f313f4b+ 1'b1 ;
assign I6bbf2b47a7dc50e66a3d8d258d6e31fb =  ~I84e4b3bc63ec0b0bff7f98f433c1fd67+ 1'b1 ;
assign I8459abaa907f5afcd11884b1ec8c06c5 =  ~I78c6a1428a1f211c5e89b8c76b3dc033+ 1'b1 ;
assign Ia16ae2f6ef5000d47b6b84ed058252aa =  ~I9897cbf9d7cab759f99f5f8f4bc125d0+ 1'b1 ;
assign Ica32690dbc9ea110fefdce92260b125c =  ~I9a6c1ff6dde5141849e4aa925140ebb8+ 1'b1 ;
assign Ic431d9383cce30b1889c92e2be4cb9d0 =  ~Icc1c25b229393361f1245c40f573b423+ 1'b1 ;
assign Ib9cca4c0e58373c26d5fd9f51f793898 =  ~I53b5a72e41ee53037ee3ae040799f401+ 1'b1 ;
assign I99bf0bc8ac20832b3724b2753f6ca449 =  ~I3cc25fb583118f45babf457fe78d5434+ 1'b1 ;
assign Ie701008f3c60c51ed72c5f964a8fc36e =  ~I20c046dd8a1265e12e902275b73417da+ 1'b1 ;
assign I3e2d78f8307a1787f8b2eccba94c7557 =  ~I1b184c9a34aeb6eda813d86556e235d9+ 1'b1 ;
assign Ic1b4444ab0df9745d29bf893d9b83168 =  ~I70e03db993e1d26d5814ff5fcd38ada1+ 1'b1 ;
assign I5f52dbf600656a8f5dc6b6b8a45ccebe =  ~I119dc168a44950d215af877eb81152fe+ 1'b1 ;
assign I7f307af79f45ad4b9511e3961c917078 =  ~Id717ed42457eb1d3f4e3edbf0dd72c41+ 1'b1 ;
assign Ie17a5be2a16d2efb98c976d7ee882535 =  ~I79d1f852a03bcc11d6121a12d8c5b86d+ 1'b1 ;
assign I5f19d2adff2f34a4bebe03f929a09c49 =  ~I769e650e49f152c0803b06232740691c+ 1'b1 ;
assign I3cd69aeed9e869a2096d6dced5c209a0 =  ~I1ef3c09b8481f14c3526224430a5f4b9+ 1'b1 ;
assign I359b6a22c9568a13b81670c741281393 =  ~I2a38d43a7e25050aa672cbf84a409aa8+ 1'b1 ;
assign I24ba99614df383c38bbac50ae8b4487e =  ~I1c2be5e13c462a8a6b07bca311582ce4+ 1'b1 ;
assign I7498bee46de6b1c946ce95fdcc89f6e5 =  ~Ie8fd61caf16aa0e504cc7dc8cec6f0b8+ 1'b1 ;
assign I0f644f42cabf871b71e5a82871bc7b5d =  ~Icd0fe98ca873ad6dacdf80dfdfc450ec+ 1'b1 ;
assign I71f9e059726a6cac8bdf0efcc0eadd2b =  ~I94e1ab698dc93ff0764dc5c1e62179fe+ 1'b1 ;
assign I0c9b2c1da30bfab514bbb556ae7bd4c4 =  ~Ifd48363af9abb390a72991fbdd6f7877+ 1'b1 ;
assign I7918b2e37e96aee94fbccca7e0f75fc4 =  ~I44f79397a010088e4ecdcb9669f2efbd+ 1'b1 ;
assign I76eebd77eb77e0abcbc727d2c511370a =  ~I124b0b7d91cfb42b0d9722f3229c2d53+ 1'b1 ;
assign Ibb2288e62110bae5b2d3fe901974e5c7 =  ~Iadf1875c584adc34f7586a146184a763+ 1'b1 ;
assign I080f931dfef9d8adfb1dc1ee073eb64c =  ~I02d3f9982f02ea85f996bf5b5975b930+ 1'b1 ;
assign Ide1106431e3565158bd81ccd6b18f3a1 =  ~Ia6e1b39d83ddce053518c5ae9a5ca33e+ 1'b1 ;
assign I63df19931e8d28666cccd79922cbd418 =  ~I3308663053f4307d43ac66f43266f706+ 1'b1 ;
assign I9a7e4a59447048de90446f877eb06627 =  ~I87ad25dff6c0c9ac46b7a129cb575537+ 1'b1 ;
assign I0917e92ed84363ca92fd2074acd74eba =  ~Ibf5d40b7c46b50866f58f6fa23e1861b+ 1'b1 ;
assign Ie3eefdf7b5561a90a6ddd9e6aa432509 =  ~I0e3a9a3b38875156d15f697adaf95410+ 1'b1 ;
assign I56eeb10d11e886cff629457a640a1c76 =  ~Ie3f87d094e71e4a82f60e8d91cdd768b+ 1'b1 ;
assign I7a9eea89c4e76d856df44b6bdc332840 =  ~I793f52d174cd09fe000e8d0351753592+ 1'b1 ;
assign If8d8f4333e893788fcb9ec54256e5b7a =  ~I89ea3da7db40e7e6705020462b2d1df1+ 1'b1 ;
assign Ie4af0e7e04778d85f5dee73da33376a8 =  ~Ib2af2f1a928dd824f25b99f0b602753f+ 1'b1 ;
assign I019a4e997adf54f5f5ca651f80b7901b =  ~Ie3e887f5f1a64c37a10404d636212b45+ 1'b1 ;
assign I10294667f09abbfd4e2f757c414072fc =  ~I5c6a004278f155d33d0cc1b576c3b25f+ 1'b1 ;
assign Id4e8ab8f15b36bd27d1e4ebc5cbe1495 =  ~I6a03a4a548a0906d1a3e9ce47f3454c6+ 1'b1 ;
assign I6c93588ca9e7c623d75314da39e89a91 =  ~I542e525074d049197ac3904e6102f0bd+ 1'b1 ;
assign I1020412efc78d12a9ebcbaeb83e5dcea =  ~Ie0307a43ce71ba73d4c8e5ad556bd341+ 1'b1 ;
assign Id0b574f35a83dcfd4481a10043cd1884 =  ~Ib03e1d3a1f27721e4ea32629c2e86f85+ 1'b1 ;
assign Ifc577e5c2c7288373a8c5e3969ac1589 =  ~I782f4ab4666c9f550a2cfc943cedbe77+ 1'b1 ;
assign Id18a1a17c1cf6e8a2492aa73b62898f2 =  ~Ib991e16161d5c8b3b655e3c7c08b93c4+ 1'b1 ;
assign Id8ce8f636723b9f119bb86c25017e6b3 =  ~I72f8c6bad4bff3b00055aa8824479931+ 1'b1 ;
assign Ic29a18d8d504a2d5280c1d7771346518 =  ~I58e5100cc1e9b809e93125fe5d08a9d8+ 1'b1 ;
assign I96a79193aa2956b8f901d5fcc9cf65cf =  ~I0aa7056fdacd6022f328a3be49048856+ 1'b1 ;
assign I8c97a246c749fbef029f8b1671c772bd =  ~Ia2f40b5c49a2284fb6a234bf7472130f+ 1'b1 ;
assign If9ba9d221909ce7499725f6fd7d519f8 =  ~I8da184aee7953890f2c89e40744402f4+ 1'b1 ;
assign I53a7878f44253f0f1a82d9d27b1a44c3 =  ~I613ccfc7dad5627cde02fa1720244d01+ 1'b1 ;
assign Ie0e928125f9d3d17d123d97e00f1fc34 =  ~I080fc6c99e506e569b97433f3fdc3e60+ 1'b1 ;
assign I2bd0f77efeca09eebe82ea234e9fe638 =  ~I79aa118ef8ac0d9b13723fb1f5a7e4ad+ 1'b1 ;
assign I94f2e7ef9b3463bd598dc9049f6fb0ef =  ~I7e6e7601245ca5b3a58b91848e25a6d3+ 1'b1 ;
assign I6dc16510af6b61b79b339d0fce77ac24 =  ~I2792edda66743635b837aa3bec0c58b9+ 1'b1 ;
assign Ic655e213ab81f5d61a018d3ed7016b12 =  ~I085cc29465c945957d00cbcf804e3ae4+ 1'b1 ;
assign I2ffc4a604025a2f5c4e273c1d070a725 =  ~I74a8e879666bb216a331fd2ab723e37c+ 1'b1 ;
assign I1c76818a9a3b688ca897aa479f7d807f =  ~I7a90a43ed71e82862457d9fa40bd005c+ 1'b1 ;
assign I3bfee9d3d88f0569010a4e0101200c19 =  ~Ie1e7b4bd6201baa02b8d59cb0f6ffb8e+ 1'b1 ;
assign I5d4738755a26beb6d0f61dd3dec0f804 =  ~Ib7b7cdc22b22f276b1c021abaa8fb443+ 1'b1 ;
assign I2f3c800091275bcb72d1a2a38fba53f3 =  ~Ib58e33f31be36b28997ba05ef1004573+ 1'b1 ;
assign I378e67cca7c4ff6325683f8346963210 =  ~Ibec394e82f499e8d2d5a9524f943d6ac+ 1'b1 ;
assign I04c8915a7f4bbde003f7facc84435c1a =  ~Ie06ad127e475dc131859992bb5f350a0+ 1'b1 ;
assign I3f50b10072f38b6addee6845e6df9118 =  ~Ic494a58468b6a7dda76923a9475bf173+ 1'b1 ;
assign Icc60eb18ba740036d2a17f98f15cfb98 =  ~Ib82a2db86d03fe8538fa19d06e501dae+ 1'b1 ;
assign I1677daa18aa8b226753b1a887b9420d1 =  ~I5b64727fee9d0825a4ea83261992e489+ 1'b1 ;
assign I36bc2d4c9a4480daa9b0944c08b50738 =  ~Ice7e502b9c2b797719448fde8376087a+ 1'b1 ;
assign I38419a6905f50135a6783aacca0384dd =  ~I792b4f73ed7139b8761443cbc0833e39+ 1'b1 ;
assign Ib48892dcb0715987289662a14672611e =  ~I278d57d1964cbf3339db450926ef4782+ 1'b1 ;
assign Icd9c94f929dbc71c9b836fda3019630b =  ~I9c1a08b61782ef6c72545504693ac54e+ 1'b1 ;
assign I5d0249d9a772805b3fba3f3c7f5d35bd =  ~I363594fb91d01abca7a2b7402e352fd0+ 1'b1 ;
assign Ie97341deb6fb24d49eb8b96bd0fd3f35 =  ~Idd284c75a230f4b97d5acb98a8e38b2d+ 1'b1 ;
assign I17dd788f9d8e91307b6b1ab7488f9ce2 =  ~If040df53a6410b263f5b3dc3090631c4+ 1'b1 ;
assign I92ae370022ed107b152b10fd0aa3d2b7 =  ~I31df60ffcaea9cee63b920478cb058f1+ 1'b1 ;
assign Iebb39f0d19ec1208bbfba6cf67a3bfc7 =  ~Icdd2f6ce69b389fbf712e45bdc0a0257+ 1'b1 ;
assign I81861f6bb8bbbab6e93407cfb4a852b8 =  ~I8971b250393b397b94db38b9fd0fe501+ 1'b1 ;
assign I217b2e3ca0a534fc5b1910adf3c1b57d =  ~I9199e5e8fdc0e2c62ad1d62fc4d873cb+ 1'b1 ;
assign I8429b08891dc56af24c72ce1b7725457 =  ~I6e03f71fdf20db836c5772658a050e9c+ 1'b1 ;
assign If96747262303f6c5c6b129e39224bd23 =  ~I2ef49f893dbc8581725ca0f6d1c3305c+ 1'b1 ;
assign If7012457af15c405baeaa1710319b541 =  ~I8796f168c892ac60c38a0a7f1e18035e+ 1'b1 ;
assign Ia0a0229ef71b85195352bb664ea4e4e3 =  ~I64a26e5117c8f3ab95bf0dfa97427243+ 1'b1 ;
assign I42aeb7c23accc2ca874c7f8221c3af93 =  ~Id7946a0299ced3ba00f6c3e6e664931f+ 1'b1 ;
assign I7df6a95bf51f40693c439c6df36510d4 =  ~I5243b90640ea4680de83021601c85c39+ 1'b1 ;
assign I8fe65f9c344d7ec8657f192abefc3fb6 =  ~Ic8301fceed328cc031640ecc4ff34803+ 1'b1 ;
assign I4d75c95d34d8d8aeeb528456bbe136e1 =  ~I6e852c94b6105af62ee85f8adf77fa55+ 1'b1 ;
assign I43746054a38c9521f8da9db9d0e91f99 =  ~I7d98c5c2a54832b6368ce60009208eb0+ 1'b1 ;
assign I0430ac2a4b2b2e2fc7f8154bf946553c =  ~I7e42f2281518bead81a6d18d2dcbd1a3+ 1'b1 ;
assign I25dc807fd55b81c9f24fd0d1edcaa758 =  ~I63c126c978154f2d68b11f08a938dcb4+ 1'b1 ;
assign I7881184f1779b9fd4fdf329c5f7664da =  ~I2ff7719c35578b47720cacd9ddfd92eb+ 1'b1 ;
assign I8e6de2d692a307ee8a5a4b2a9265a633 =  ~I480599aef36967a670155dd77120a37d+ 1'b1 ;
assign I54b2b18ab051b468808a3d0fc4bc893f =  ~Ic000b2c844de484b8f30b7b84dd6234d+ 1'b1 ;
assign I37ee86e2ca32832862cb57efe76bbedf =  ~If0e25df151db991185f992eab5d5be99+ 1'b1 ;
assign Ic95f2fc697574803c0f7fa35c2609f0c =  ~I2f533699abb7a997160bf4ee4cda3efb+ 1'b1 ;
assign I933a30c52c9bec5172530b2d739a3b63 =  ~If6b33cfc6d34e33fbb18e08fb4d8a5ed+ 1'b1 ;
assign I7bbd7df18f85197c22fe8cfe37312af6 =  ~I2ea5423dc8726fc0217899e0f406a1e9+ 1'b1 ;
assign I50d5ada7c91c7af16492c6b41151b68f =  ~Ibf3f4f8a04cbacc9624ca5cc73bf7069+ 1'b1 ;
assign I32c8e7996b3473d4906c40018799a16b =  ~I9ba53c36934ab1c7f498241a79cfbae8+ 1'b1 ;
assign Ic0eacd5a4812ad7ae3fa251ab2db4694 =  ~I106a25f18536f96782927bf3bc2ccd72+ 1'b1 ;
assign Ideecf8ab87d28a840cd93851169ab05b =  ~Ie5cdad65e918679607cc5f816987b736+ 1'b1 ;
assign I1ac6775eb38457b7962241d2e7336b0d =  ~Ica6dc9ded8756fd6f82eec4271e246c3+ 1'b1 ;
assign I2ecaa89698604fddd863d7e28d643a57 =  ~Ica42ac6ca5813d0d1a67f14d1248437a+ 1'b1 ;
assign I273e0fe9c51c8549c8dfff393ca2e4e1 =  ~I13dc6cfc75ef846c30e5dc1dc5305d59+ 1'b1 ;
assign Ifb1fc76002f6920a1f44c7b1bbcd0020 =  ~I33e784182dfb4af39715788b1ae98af6+ 1'b1 ;
assign Idf6d4e3aa753aa396a9bffb27732f851 =  ~I9e1a66805348d2e5bbf5e2316187444b+ 1'b1 ;
assign If14ca1f5d1c2977f9da79eaebaad1bf9 =  ~Ie9619916a96d218cf5eb5f3a4995d0e7+ 1'b1 ;
assign If8f1505d9f10e30bd3320f500d34932f =  ~I02ce7969c51ad141df227ed7d18e74b1+ 1'b1 ;
assign Id32aa77c6406b35a00168bb5452b12fb =  ~Idd73461af0d75c4d820f7f8f0f419e0f+ 1'b1 ;
assign I9a73686acefeb361337511f6943b036b =  ~I3df6c2cdccb2a82c58c1d81b00af7786+ 1'b1 ;
assign Ib6eb7ce5a070f3a87bcf0e18be8c855d =  ~I97f441fc5ffb88efeb5ed66b60f07a7c+ 1'b1 ;
assign If69b0b717c35d33fc8c0e59b07eb9edc =  ~I3194a235eb652c8d0e4307cd056e5e72+ 1'b1 ;
assign Ibb0d73078b779585e6b0e228391ecb96 =  ~Ibc315f6c79ba2bf336ee57f2e5f7d776+ 1'b1 ;
assign I2894546e399fe3e33d7579772a1310df =  ~I937a54f5cda99a7079c7fa46b4ea26f6+ 1'b1 ;
assign I97f99a266267859aed199b278a430417 =  ~I49c99afecc613656cd1469d8c1e98936+ 1'b1 ;
assign Ie18cc792329941a3654322376a937d8d =  ~Id76ce0333f43bf7bccf1ce48e25ca69c+ 1'b1 ;
assign Ie914a99f08d60b74c3c36a632a4ca9b0 =  ~I2c77f9644145219005751f7a4eb71aaa+ 1'b1 ;
assign I82916e9dc3894ad88e12de01a68d6aa5 =  ~I5cecc266272eef88cda88c1df9bcc37e+ 1'b1 ;
assign I6cbf576b3d652e34c0221f8316b5a392 =  ~I776a0b1b5c14afa21b7fda3c2cacafed+ 1'b1 ;
assign I9141b2516d7f855cd186472780af7b67 =  ~I84860b1f933339e0f90beeb3d666393b+ 1'b1 ;
assign I07bf32ed72de9c02abf700c64853af61 =  ~Id24581713f1ecb767db39d5154c2f5f4+ 1'b1 ;
assign I52663a2999fb9571834d517538691b6f =  ~Idb0eae2f0e1dae1d56251d64e2c51f9f+ 1'b1 ;
assign I8dcb88c94506367aabe8d7ed62cc56c2 =  ~I2e3ca4b130e6d3d92385928a28644452+ 1'b1 ;
assign Ie676a4bee61154145391d9cc473fe91d =  ~I7922d80ae333dcfafde31d294f0eb4d8+ 1'b1 ;
assign I9502c8fbf6b48749bf9f84a89a937dfe =  ~I82de04cd2dfef5616efca4af26d7c561+ 1'b1 ;
assign I0c91e540e7106f32ae59491d8ed1853e =  ~I7ce384520525b15d24c2ef6f161213a5+ 1'b1 ;
assign Iddfb8a8e261389eb4a2a10880c19446a =  ~I56aeea71c7bd19d47620cf36adf3f115+ 1'b1 ;
assign If0d55f861d4b3f0970c529024ca142d5 =  ~I138e1a6db0c6649bc023cc36d81d5b47+ 1'b1 ;
assign Ib054f5d3f5cbb29a053d0e50c23cb3a8 =  ~Ib5e8b1c4dd9b5dad56b59cc11c87a258+ 1'b1 ;
assign I1d65e9f97e93de8cc2a5dd532f8e482a =  ~I86f785e2d5e8d6c08fad1d334c7d244e+ 1'b1 ;
assign I3bdeab8c87325d46e45d9e2d44756934 =  ~I9a6c8efca218c724da4ee4c1087d58bc+ 1'b1 ;
assign If9228f7ecf19c41f4bbd8dabd0d5816c =  ~Ia30e8dbc6974ea94b763842e8dffa633+ 1'b1 ;
assign I9e3edee214c4937d2aa462d3cffa624b =  ~Ifa60f45f4d8848eb0b89f5644ec69668+ 1'b1 ;
assign I9fcbbd2e81b006b50e2d35ed2627bf83 =  ~I0aeb4b93cfa6d62ec41b7e6dd0287dd0+ 1'b1 ;
assign Ie16f3d50ad5e5581ca099549db7232d2 =  ~Ifce1fc978fb5b0187593f46f53c3b469+ 1'b1 ;
assign I6345e93f3fa7f5eb2008dd41742afc2d =  ~If3b6de7c919c5d53a0e191a75bd7e574+ 1'b1 ;
assign I698b93e10073b5d29357cde4bcac9dbe =  ~Iecce594e6e99b0c05fc845144a664b07+ 1'b1 ;
assign Ie7ced910d84655790823e6173a5a314a =  ~I2c8431500ecb25619d2884a2fb4260c0+ 1'b1 ;
assign If6e3b6fd1810f6964e9024329d7cb3e3 =  ~I217c710f7ef39035546efcbb043f63f3+ 1'b1 ;
assign If1045908c6d7476bd5507e57d08c406c =  ~I1b4236130cb1879d885653fdd9eeab4e+ 1'b1 ;
assign I4d4f6705ed77a16ff31b34bae0d8b6d9 =  ~Iae0f7c13f1564d63b4bfdc152ddf4111+ 1'b1 ;
assign I70a492396580ac1143d8a2f4b181e873 =  ~I010592496030d138a3a4245d00069957+ 1'b1 ;
assign I2fade32b5bdf245fa15289620dae2670 =  ~I9d7f47a6289a16448221d61f301586aa+ 1'b1 ;
assign Ie0dc166f57fea074496241a32cdb6015 =  ~I7b8ed2953170c4deadaeb33a6ba165d4+ 1'b1 ;
assign If6a2518891412caa6d6d507082501f1e =  ~I4efe9eef6a48aeb0a9ba4e0ffd9906c3+ 1'b1 ;
assign Ic9912e5a838a377b26a19d22148a64df =  ~I5a8466bbd83c39dfbeaa6399e3fb3337+ 1'b1 ;
assign Ibc0fca22d16444bc17877106ca772c31 =  ~I1ab96ffa948dd09bcc4f748c6c2575d2+ 1'b1 ;
assign Ie4291d233597d5d676a80fd62d9bd208 =  ~I016f57568eaf00b26f8a22100858c158+ 1'b1 ;
assign Ifc13b798d76aa70ec1877c275fb31d36 =  ~I1fb995e302f4f1ba493ff85f39938175+ 1'b1 ;
assign I57d6637f0bdab578a790e4a12ccaa16b =  ~Ie643ad235307c60f1ee96dfdcbc8c2a8+ 1'b1 ;
assign If8ea04fe685b4f20cdaf9a84984d56fe =  ~I8dafdf2c780082d8dfc2961b3447f104+ 1'b1 ;
assign Ie0c86f20c28bcbe410b191b90d29bf76 =  ~I3a2841a0f5e1b42556f384231ab0717b+ 1'b1 ;
assign I3dc5d3f66726e15968a70cbf3d3b656a =  ~I2b00d0e6facf01274c0c3446bb0e1599+ 1'b1 ;
assign Id674686e7ac37fd6f63846f9a9cede19 =  ~I2c645d25871b70dae5b2c283695d5130+ 1'b1 ;
assign Ie2ed9668d13d219c60f2e0614488cd42 =  ~I540a0e8968a6a82aca775a81ef82b520+ 1'b1 ;
assign I98abc995ff89934534543be93c6e3ffa =  ~I5b95bbc82e6d8d87421efe3f17b97ea5+ 1'b1 ;
assign I579cf9386ab7b08efa204d735335e462 =  ~Iad81f5e5e728ffdec6296b2aff668d75+ 1'b1 ;
assign I9efa4d729d10a6b7cc335fb765ed032c =  ~I960a618f63372da74581b8c352f3e618+ 1'b1 ;
assign If9191ebc8e88d4e75f0f35897ebb1421 =  ~I4f5325f1601acde10018d1fd0aff4d35+ 1'b1 ;
assign I3511287cfe69d5cedc5a8fbcad708437 =  ~Ib297101fe456520e72cd9d208af44eea+ 1'b1 ;
assign I91812179d44cb675b90d477f33ec48ad =  ~I73a21342321a9d81a0fa5308149d72b0+ 1'b1 ;
assign Idb04a1aae91fdc477ca38ed66789ee88 =  ~I2a486524f4f53b3454ee02a8892d4fa3+ 1'b1 ;
assign I566054aece562960590ee28b157e4a3e =  ~Ic6c4e4e6a9ba43a3354f9f3192ab069e+ 1'b1 ;
assign I7b2ffb762cd9ef7aa8ba224efb75c46c =  ~Ie3cdee3560bd06aed84dac5fcd2a259a+ 1'b1 ;
assign Id90bbb642b0f4434d8a148a28b6b2f65 =  ~I584febaa4c440fd9353108af36d3a5c6+ 1'b1 ;
assign Ia4e297e35d484b15adce7e1d67f582b0 =  ~I515e78507d7419ca14d77b6d52f75a78+ 1'b1 ;
assign I84996b1d03b692f6f736fb04c7f91e83 =  ~Ie9578453a57d2b3b9c3b98844044b5f0+ 1'b1 ;
assign I83078cc7857fc17b30f640854a4d6be5 =  ~I1e58b3062097a46d8d590232b40278cf+ 1'b1 ;
assign I94bb467129904032736fb13dd636c600 =  ~I3af126eb28c67797ce625b0d82943833+ 1'b1 ;
assign Ifa76758b50f439170ecd6d86ff898bc4 =  ~I130ee1a8acacf4cae8818cd8320d050d+ 1'b1 ;
assign I9d831dd976e8cd5d8f6a6818601e6424 =  ~Idf92dd09c29ce8e921b2b34089550586+ 1'b1 ;
assign I474774ae149804412ed4aaf1cdcaba88 =  ~Iba74a64cc1d2ec3c83a4061db298ad37+ 1'b1 ;
assign I964cdcb4e6b49a62d30c2a2540851317 =  ~I01364c233ca541914d790354515aa5c1+ 1'b1 ;
assign I6df268bc9f85ce88674a9165664ea84a =  ~Ic6a8297308a63ed3113008a3cdc76358+ 1'b1 ;
assign I74fdcbe9f49f7bce1f5e31d956c5883c =  ~I6c7ee9d0bd684a7f54bed3d52452219d+ 1'b1 ;
assign I4a1b8453cb7a21745d5f74ad05653ed2 =  ~I985ea87550ec8a222e6af621589e186d+ 1'b1 ;
assign I9c53b478b2011fac0615a152fe60d5b6 =  ~I6836a7d1e006d7f7556edf8b31aea32e+ 1'b1 ;
assign Id75dbed8f1a5befda32c60b994681013 =  ~Ia7a356a18af18ec131b9df46019f3e58+ 1'b1 ;
assign I378a59323b74623c5524f854d6e11226 =  ~If3a7e111247232c47ceccb5e05338312+ 1'b1 ;
assign I080bf885464a0cc948a4450e9f7d1d26 =  ~I5f38d1665294b2d3c18f9cd888ff60f1+ 1'b1 ;
assign If769e73adea227de1fd85c2e89d0ba08 =  ~I10290b9576bf3d8caf90583a388226b7+ 1'b1 ;
assign Ifa6a34b83225e9d9b28b14874c4444e3 =  ~Ief36236305fc1521c5bb4c60753a676a+ 1'b1 ;
assign I584b1d4d6fb7ee4f20ad9c96715cdf90 =  ~Ibaa0539fbf5ccc979511c09c061cf494+ 1'b1 ;
assign I265f9b91fbb62164e589dcf96818c4f5 =  ~I95664ffd0ff13c2893421032149f24d2+ 1'b1 ;
assign I3d59a47c88227734cf6fc0d6fd30db11 =  ~Ie390153b3b7985dc63d65913de215377+ 1'b1 ;
assign I6144b6df2c87ea0948d730343b42129f =  ~I704147dda658f4a03627dacc1c91dd48+ 1'b1 ;
assign Ia7ca7400e36ea572fba8e19bcc81ecbd =  ~Ifb09672d505898f081aa13c95fcb88b5+ 1'b1 ;
assign I302e61b49accf5db556b87517f2341f5 =  ~Ibb5cb89097dd11bf292d5b5a2422175b+ 1'b1 ;
assign I5d9af1abff6efe3a55c6568d936b6ec7 =  ~I4a305956b18d6ad6901d2c17e99f2bab+ 1'b1 ;
assign I8cde0aa611c476b5112edeb8f17f15bf =  ~Ibf5bb3b9eb1812383db9634fa9a27ad3+ 1'b1 ;
assign Icaa40ec40d6d26cdf70bb5ae7d492e47 =  ~I66b37d055c3735f011095ee4b1ad02ed+ 1'b1 ;
assign I8346f15d822cacfeecbe5d75412cb53f =  ~I43e71dd694d97217e242f267248cd594+ 1'b1 ;
assign I5ee364aab320ab40c0f65feda6f53b18 =  ~I4baa925db1ec733bd4bd25d9dc873e23+ 1'b1 ;
assign I1f0ecba054900f96cd7100741191c5f4 =  ~I547928c9db7acc531af251264d576ffb+ 1'b1 ;
assign I4faf2caf62966416118a54015908c889 =  ~Ie4ce634b2fb62a20781f8a2e8fddc762+ 1'b1 ;
assign Idd0329980a36f87859150530ab44b52d =  ~I0e90e96ffa64c2874d79110b622994bf+ 1'b1 ;
assign Ie66bc10dde27f08813d4d347fd7cf6ce =  ~I767e37e3c6f4224eb07adeda480ce253+ 1'b1 ;
assign Ie1d8b3ea7c6603cebf2f9adb776910b7 =  ~I75fcaf2c65b7e63adac834054850c6d6+ 1'b1 ;
assign Ia37488e9a50cf5cc08de74ade676db96 =  ~I5f1de2dfbd79204ab2db9b686d6a6862+ 1'b1 ;
assign I08aa45211cab01d567cd5eb172fd2f0c =  ~I8d01de6be4091dca2589cef625c05229+ 1'b1 ;
assign If4ff0c63ec1deb46412858e496451a01 =  ~Ic09e773899fdd208c0fdd874933b2cec+ 1'b1 ;
assign Ife7bfd15fc4c392b5d2288d9a4e879b3 =  ~I24a3f9fd851c4af70ef66bfcee44af65+ 1'b1 ;
assign I24ac26debafd03c7333d174e8725afd6 =  ~Idd31807ecd603db8c719349a2be1be40+ 1'b1 ;
assign I99d80ad68e2563d0f78a0e3bb82c5328 =  ~Iaf680cae40d1adf7649da12b31a2be0d+ 1'b1 ;
assign I9943733ef305983c629565c881054bbf =  ~I22d948171c1a66f7a28d5e51007700ea+ 1'b1 ;
assign I7cb4420bc55c03a6500f5228d31fe43c =  ~I3954318b2392a82f2da71a0ca1504497+ 1'b1 ;
assign Ic4d19dec464359c0a9fa75148fe90c73 =  ~I15c78b909cbd04fe25820d777655d829+ 1'b1 ;
assign I44993416e1d22613dbd78402c37a934d =  ~Ia529c5ec88a9f6c14ceda5cad56b346d+ 1'b1 ;
assign Ibc9b94a9dea471805cb442ac6904bc97 =  ~I5b73c81f28901705f6ee26d63847db0a+ 1'b1 ;
assign I917d9f9b144d3bffafc77bddae7fba6b =  ~I1a9bd3f728db23b679639e5657ced179+ 1'b1 ;
assign Ibc91c6c3d56bb8a14e22909c43ffec51 =  ~I57ca72784a7c91cecbd694ddd08bcb98+ 1'b1 ;
assign If7c2d3eddd96b47b6c2aea8b27c8c7f4 =  ~I50f31ecd3f2b498cc7b759efa057f12f+ 1'b1 ;
assign I4df093ed94d26b058e97db550e347e3c =  ~I8ccaf29848defdd264f522642968fa29+ 1'b1 ;
assign Ie90303b0326bee4ab203a8cf1e643da9 =  ~I808ea92ee1340876cf1d2c47255dc2fe+ 1'b1 ;
assign I19030d352fd059156ee42c66f9270beb =  ~I3da806790125328b626be1949f71267a+ 1'b1 ;
assign I36767a902c53a384128ae1443cf88963 =  ~I55e59bc1daeb8b2be3d7a1e4b272df93+ 1'b1 ;
assign I868dffa3f07407f7996bb5bc596939b7 =  ~Ib0ffadc6a0091ceff91ad1fa435413a6+ 1'b1 ;
assign I7d928be164d0dce8b1322ff230c053e9 =  ~Ic863f139e6bed2d06789a07c6dedf6f8+ 1'b1 ;
assign I98be4971a8a9a08abb3ebe474d7f0c6d =  ~Id0e8f6ada5060a911090f76cfaa3c6bf+ 1'b1 ;
assign I779e70dea33201e9237f29681ffd5e27 =  ~Ibb8c9b8fc9b58f5f8a6ad342934804a8+ 1'b1 ;
assign Ie2262914042172ab7e08599278f36af5 =  ~I9323a188737ca54c2dd553cd99bd416c+ 1'b1 ;
assign I4001323da8f7956cdd480ac2d56df929 =  ~I2694cef38855f496e7ca12f42dfdb9fc+ 1'b1 ;
assign Ib1cd6731034887a0a55e405c9db3e8de =  ~I75790b4c0b1f6c7935f5cfbea26407d1+ 1'b1 ;
assign I51aa496e8c03944c28a908102514e6f8 =  ~Ib8b366c47e56a49fc53ea4a9e1ebbd99+ 1'b1 ;
assign I6415f3996318472532e161510ccc8ca3 =  ~Ie1c86256df2bc6c4dad41237eca41986+ 1'b1 ;
assign Ia11b671b59240988737979328c472812 =  ~I7c9e3f97a94f9a078c209a1b84ff916d+ 1'b1 ;
assign Id4fabe0165a117a402dc14f2f3ec626a =  ~Idde839d34403fdbba62671b83801ea8d+ 1'b1 ;
assign I57238f501ab7278b308d76211ced8cf7 =  ~I824e23c3e43434e0a7bf8c8b8e0de597+ 1'b1 ;
assign I9b257f8556ca4e5402637f01081b78e1 =  ~I0f83a2c488c229e971030fc66ce212f5+ 1'b1 ;
assign I2e093412a9fa3972cea01664389d8c27 =  ~I8fdda3dea7a63fd6e57f70365d7b6571+ 1'b1 ;
assign I17907fd8c6975c8c642535ff929221a6 =  ~Ifa2fc30c14c549339edc65c3670d90a0+ 1'b1 ;
assign I3c6577b04ad56d864bbaa2c048323c11 =  ~If69bb1bfa10ca7dd37ba57485c3429e7+ 1'b1 ;
assign I6f0c341c05eaa8f35bbce4521f6e8f94 =  ~I2ab0738fa2d5916d77a81b9da2315376+ 1'b1 ;
assign Ib72ba950ecf9ae2668374f6633a67ca7 =  ~I50a9ce776ad2ccd8048b56ce101c80d2+ 1'b1 ;
assign I3d7c72d725f4563bb562e2992093cb02 =  ~I9c9d0332ee7ad6a3488b7e39bcb06ca2+ 1'b1 ;
assign I813c881ac61a59041be3be78f6a466c8 =  ~Idc155814976f0aef9b56b2bb3d52b3a5+ 1'b1 ;
assign I866510e7dc721fa5aac312bc5ab5ba0a =  ~I2e02fbd496d08acb3ad3359b49b9f680+ 1'b1 ;
assign Ib4432359f97849dff6ad3e0f044157bd =  ~If0f8b3dfce99a5a75c2105d45ccad985+ 1'b1 ;
assign Ic86aa6eb1b4dcc2520309089b43292e6 =  ~I6790223e6a7cf136a7e2b261ba4fdb0a+ 1'b1 ;
assign I0731115afe5c15bcf131f7ef4f05802b =  ~I6a9643afea7a6cc9b94806ccc8e84c0f+ 1'b1 ;
assign Ib080b8fd34385aa7986dace4afd95267 =  ~Id3d19d7c2b941930478a7ab01049e390+ 1'b1 ;
assign I134890b77451d0b78afc7402a6a28048 =  ~Ib0a25312d51cb6aa1741f7e425bc5cd8+ 1'b1 ;
assign I956da75f13433c1dd7a3cbd3b78922c1 =  ~I44dd1b66f5a9a6b0b976d3d61d6c5cbe+ 1'b1 ;
assign I440b26c9f1b9ccf70f97c9d5f732d38e =  ~I3ee456f2f0e7f447ae92b7523136adb5+ 1'b1 ;
assign I5e3a441faca44bffc4368d96d8fb0bfd =  ~Ic110e2a08b550acd3c8bda4a1bc2bbae+ 1'b1 ;
assign I21d7ba25247a87a1a9c245d0d1f553b0 =  ~I3f87162d2874effd66a82f821aa6c73a+ 1'b1 ;
assign I55aafa8162cfc4fccfae68cf78cd1c2b =  ~I660ea6d341fcb38f108270c08d82473b+ 1'b1 ;
assign Ib99c25f0d8d6493cac4d5c816884c704 =  ~Ic128d603fc08affd2f3d0ab3425710e5+ 1'b1 ;
assign Iee7c9f0a0e8ca127efee008b4874edbd =  ~Id5372641727970383a59e08f550814b4+ 1'b1 ;
assign I17b4a3baae65161387f472037ffc6fc4 =  ~Ie99ad992d66880542dcd330ef6ccee04+ 1'b1 ;
assign Ie7b7b202a968fe73f6b1e02a044414c5 =  ~I9ed0b194f7d210d57c54b289e01c75e6+ 1'b1 ;
assign I479ab5c0e483c36267d8248340006666 =  ~I227828831c4ad21b06ed00fb5781b0e3+ 1'b1 ;
assign I777bfe165e25d7fde4fc950f23db7b84 =  ~I09d5ad12cb836adfbb4833ee80fad2c9+ 1'b1 ;
assign I146d505a34ddb8d65e0a1769f623a7fd =  ~Ifa9c94ee94e4beb2e7c8d2d57150df41+ 1'b1 ;
assign Ia85239bddc04bf50bcf037ed2f76d7ac =  ~Icb88e59e194db215382e8e949603a9be+ 1'b1 ;
assign Ia7306bacf3c2b180d3261a5c1f0f4a30 =  ~Id4ebd28aaf1076acec266666f88a02ad+ 1'b1 ;
assign I2018147b86e47af5842c4f29d047d157 =  ~Idf0a0bd862167392357501b3233a8d8c+ 1'b1 ;
assign Id17a85459845f8a8be694c4bf1fc29c9 =  ~If94cdb867ea0fc2c5578b16aacb1acfc+ 1'b1 ;
assign Ic012b15584d9d25af38f83d0526503da =  ~Ib8c066b0700941a4fa739820ff12b948+ 1'b1 ;
assign I7f09bd4a45143a036ce04af11b9927f9 =  ~I11e0f8dc46b286bafb05f901f968e1ad+ 1'b1 ;
assign Ica32f94af6e6f3eaf2b724a2173fa463 =  ~I608537f5639d5e0cd3e80453e21f6f85+ 1'b1 ;
assign Ib750bb83ddfbbad2a2be8d1c8392b4ff =  ~I0e9d8db1bb6347c9507b645132308b3a+ 1'b1 ;
assign I3906ece39480f96020717c6243e8ba4c =  ~I17033b417fa383a2db41d157df33d9de+ 1'b1 ;
assign Ie68ce21ade07fa53c30ebf27216b03f9 =  ~Ib7f45dbcad513b4dafee60f33622b0c3+ 1'b1 ;
assign I6cc6fa167c0d2b4b62ddbeecea175ed2 =  ~Ibfbd8e00e00272f32428c7b4a3c53050+ 1'b1 ;
assign Ibddf3468ae7c27d5a4b1388e524aa9c2 =  ~I27973d1d4e07eaa49608d6f6975d0a93+ 1'b1 ;
assign Iadcb2b3acaac2e1bb505c65d3cbe4235 =  ~If77fcedbcf99f89045de87e5cae45d8a+ 1'b1 ;
assign I37cd96b8b0a4939d9a70098fd8bcf452 =  ~Ie8f8691820e7a560db8116f38dae5d49+ 1'b1 ;
assign Ib34b169dcc76daee2d1aa2b2a7513af3 =  ~If0b19af59ad851aded19970494514034+ 1'b1 ;
assign If36fc316d6ec7c7e09eae77807b37099 =  ~I98b8e05818925a4b65082fa57affde83+ 1'b1 ;
assign Ifd214c332218ac5c0fe5aded4b952711 =  ~I69317e8c556ed67630829c990f8b74db+ 1'b1 ;
assign Idcd0fc8f86e2b6f03606b818b8346e5a =  ~I9147d103cf235310393f9339f1cbb376+ 1'b1 ;
assign If486aa8ac2cfb46f936714812cc760df =  ~Ibe0b2cab6e2d3f3cc8baf3623ff50988+ 1'b1 ;
assign I2d8e5b5fdbda7d599423c38aaace6658 =  ~Idc64f1443dd2497dfaa223cda3fbd682+ 1'b1 ;
assign I6d0878fb7ec75c0a26be4dbba62f80dc =  ~I6e37e92b812099985436851da8a6ccb2+ 1'b1 ;
assign I16a16ff0e8a6685a09803634da429fd2 =  ~I057df2bf67d5580275654bdc28b40027+ 1'b1 ;
assign Idb211abaa54ac26e7379c64a63f7d07c =  ~Ie87a151c8b90942a899b8167bcb34afb+ 1'b1 ;
assign I351205eb71acb31b59d2b4470f0ba28c =  ~I735752035af159b48f53d8302bb33c21+ 1'b1 ;
assign If5660c495bf7690252783d888d1ad6e8 =  ~I1f26bc7cb30a9659a638e2ab65e1f187+ 1'b1 ;
assign I3a5229cb8e44a15560b5c7bef96e65cc =  ~If39a50e88c4a7c43428c1d15b0bfbbcc+ 1'b1 ;
assign I889b9b0828e97fe44d8366c5ef71a8f2 =  ~Ibf966c12f049d603361ad32f55b0a2c8+ 1'b1 ;
assign Ie23062e00e39ead706f5b6ead233747d =  ~Ie1b3ed6d3fdae47669d3c4cb8af8d969+ 1'b1 ;
assign I8a2589544c75ecfdc31d28912c639695 =  ~I4ec6c8d9e87224ecbe7c69d92f9419c8+ 1'b1 ;
assign I5c21c59147e9c3a74c7cbbb6f2a23919 =  ~I2acb34de8c3fc53117a7ea4f9ce7dd2b+ 1'b1 ;
assign Idacd78e24408e432abbbfb0c447fdde5 =  ~I7fa4009267e80ea7eb71194843c3b22b+ 1'b1 ;
assign I0e8b171fe5080485a7f4fef83f1f1528 =  ~I6854329daadea2734e52180a41f56bcc+ 1'b1 ;
assign Ib22c2bd76e6c29cc2f1440885bf24b7b =  ~Ifca16aebaf75b2990188de201e4536fd+ 1'b1 ;
assign I149559fccd9def4ec1ead1fdcff3c7fd =  ~I46cc26afc8475f2fb290eefc95a542eb+ 1'b1 ;
assign Icfa8fed3239748abca27a5fc17de79c0 =  ~Id746d6515cec9e60e7478898a09787e5+ 1'b1 ;
assign I2ff115fa483f080d93bada49a9566b33 =  ~I09a3ad636db96e00adac78c3c94bdaaa+ 1'b1 ;
assign Ibee4f3cd2f516c29ab68e07a640ab65e =  ~I28b3baa225a5fd602c9fee9c948ae58b+ 1'b1 ;
assign Ie495ab560f59ad038992c573de7d2f5b =  ~Ibe12ef0f56d875c7a44030882deb0e29+ 1'b1 ;
assign Ibd812def78c3a9c02f9ba45cc0413711 =  ~I9bd9979e4acc4944227a4bd62b910c1d+ 1'b1 ;
assign I98166634dc80201b0cefb01d9559c228 =  ~Idcfa802f458499150055dbe4b1ce8146+ 1'b1 ;
assign Ic2f03a980b5f0b042853ca746abab22b =  ~Iee010958cc3e9389cb8ecacff84fccee+ 1'b1 ;
assign I2807a88097d2683ebdb9e0e785e3af02 =  ~I3d74b31096917c53757c829a67cf06df+ 1'b1 ;
assign I8bebbb3a676c8506af0768516abcd740 =  ~Ic27031a9654db9459815fe0ca35408db+ 1'b1 ;
assign I31d380f34691c9fe9022035f233b77e2 =  ~Idf6ead2c37f75f3cde1d4b40cd73db00+ 1'b1 ;
assign I1ffb5675c98ab5b3c62b24eb23441473 =  ~I66a56161cd0ed67f65834b9eb0e94d17+ 1'b1 ;
assign If56424546ec4f3445853538207ea864e =  ~If6de990e26ca9e8efc009188f8a5a4d9+ 1'b1 ;
assign I31a49be4a34d9bac2e0d815097439772 =  ~I8d866786bb2dea06f5b30f6ea80cff17+ 1'b1 ;
assign I6b96a2498078953e87de223aa2236d50 =  ~I01ca9a1d4901ec9b2a64300617ce4cd1+ 1'b1 ;
assign I79bf36e298a85a42c7432f877055f0b4 =  ~I2dbead35e15afb9affaa6ad4edd3829e+ 1'b1 ;
assign I90c070b9bde5da05e8a5d25d2de3ba6b =  ~I83c57653e24cc09214075b04b06bad83+ 1'b1 ;
assign I28d0e4e6d772dd58d845d91952ada300 =  ~I56b9c1f555b24c2dc197168decfdb8d1+ 1'b1 ;
assign I7232b4e277acc6f1acefcb606ca24508 =  ~Id5c48111f1b93de2cfe89f92fd182b43+ 1'b1 ;
assign I32da124c433c55f692ffa4734d0dc8fc =  ~I32908c3c90ed6488357ce4869e8a1721+ 1'b1 ;
assign I56e487db14eeb8d93f494d2f11b57a49 =  ~I16b4601f2e07e6cecdb5a030178e75c0+ 1'b1 ;
assign I94d3c02bd5b8e84926d4b3c2f56efeac =  ~I0ae08a41ebd0e6b402a4980478087bb5+ 1'b1 ;
assign I0c35b2e9176f9a06e26ca67d036411b4 =  ~Icb57267a66f117943e964dd6420d7a58+ 1'b1 ;
assign Ia6ee7b70d0b7fe7c346760b1784e50b9 =  ~Icfa47fb87b74106cd3814adfce909424+ 1'b1 ;
assign I7ce57c278c683ad045526e49bcc47412 =  ~I63067cef0e1a348a3e6d8cd9bd88b907+ 1'b1 ;
assign Ie3d3e681cac0bb919946ac27057409e2 =  ~I10aa5ba0f53632578c0e1cefa4bf4fde+ 1'b1 ;
assign I8ea0a8cdd6506c982ad75f23136bcebe =  ~I427c0215d0ac047e8402c20610676752+ 1'b1 ;
assign Ic812f8bc775c5ee6a83e2b9aeb22b2a4 =  ~Icf4efa87688bd1b80437686eb0126057+ 1'b1 ;
assign I0f0adf7fe957b9a68772bd8a1bc163d4 =  ~Ic373f785ddd1bf8eccce263df5a82c87+ 1'b1 ;
assign If09562f8d82bc1dea7c38ed51523a889 =  ~I56f8e8d2d7052af26528530d389b6dc1+ 1'b1 ;
assign Ib0fd21d66cd89c4e5c95fbc9c7680b62 =  ~Ifb145bc18d435fb66779e7415417bc0f+ 1'b1 ;
assign I5a2b2bfadc638fe3fdc31136a8f09a8d =  ~I62a6e0c9952d6c6e6095e2364df93078+ 1'b1 ;
assign Ica914d8c556285d6b90b35747065a6e5 =  ~Id6405c2b2b9aea6bc457f1064d5f3ffa+ 1'b1 ;
assign I00c5d739bccb0ab6d05da70fe51aafea =  ~I079df9611bd81f672f2ae028bf267995+ 1'b1 ;
assign I18e448761bc014ce490b766183350312 =  ~I096b226cc511363946a39307a7d97867+ 1'b1 ;
assign I1b5920f488e9469bd416a6af3072a30b =  ~I4cc42c5a75ef339510ee0e86fb44e16a+ 1'b1 ;
assign I70b41ffed4b6d88ddff219c567b8e968 =  ~I680c01c3327cb9372a42c1ec5b4193e3+ 1'b1 ;
assign I935e083b4561da7d015e98ca7f02854e =  ~I83451a072082194ecb3f9419edd728b3+ 1'b1 ;
assign Iaca9ef263bf220d786242b88c994fd21 =  ~I52ad85b6a1c822ca8c2459bde8fbd510+ 1'b1 ;
assign I92169291959eb33452b79bfd32618cbc =  ~I1c44d2ef638825862061a8ee1a0a2f95+ 1'b1 ;
assign I126dabc3ebb9c4157adf62b57f217bd0 =  ~I8fa1fd425809cc39cd8e2785773c1d7a+ 1'b1 ;
assign If4433b1ef2eb963cd301946958b69884 =  ~Ifa22335f04d35680eb8cfec8f862f357+ 1'b1 ;
assign I67ac5b9b794787b3c4738c3366689871 =  ~I6aff673c27811b81530453906312aa9c+ 1'b1 ;
assign I4f022d70078c412bdbef158f750d3da3 =  ~If674ac0540f457a21235664c213d4923+ 1'b1 ;
assign I6be6165385f6a77aeedb88f2baaa9cab =  ~Iac223ac498bdcf2cb2514582aeaf76f3+ 1'b1 ;
assign Id1f7fe91547e158e1d39edffb1421ff3 =  ~I7f40931ab78ededfcb52ccaac9b81282+ 1'b1 ;
assign I7a51924134902612db53941390891245 =  ~Iab7c8dad0ca20eb0988fbd99f25591a8+ 1'b1 ;
assign I45128b9e29dd2fdd94a78fc5ffdff2b1 =  ~I3cb5f890a5bd3daaae34c8dfb6ecfc49+ 1'b1 ;
assign I7f1082408c8ebb5be18e8f71ff9510e5 =  ~Id80e145586d7e539a6514dd67ebabf6a+ 1'b1 ;
assign I655ebf19c2f4b3dde716668f9ce12e59 =  ~I01e09bc554768f30dc490041d19b4da2+ 1'b1 ;
assign Ibc9d493a507122d92af42d858cdc4c61 =  ~I0196f7df6f834ae20c4fdd127e66104d+ 1'b1 ;
assign Ib3d3103e5ee4feb160a97c7e26f7102b =  ~I4669c4f256c123a0fcceb55c1e72193a+ 1'b1 ;
assign I6cc56b119e72175df3b7ce64dc3d9305 =  ~I4a02ffa2a79df824f406909aa189a404+ 1'b1 ;
assign I57cf4a9378f1cdd94a1a5608dc57e05f =  ~I3117e5029119e70846dff61d746699e7+ 1'b1 ;
assign I4160ab1aa18e8151c0a5c23b9edeb907 =  ~I1e4e705b3bda1451fc384cd934c0bb52+ 1'b1 ;
assign Ia1f183f2d904d006e46399424e06c614 =  ~Ib5bea8e0072de3de2c8431ea6a35dd51+ 1'b1 ;
assign If979702738671323995e56108bc9376c =  ~I7d9d94022ea95ea01cddc237f3df8cb8+ 1'b1 ;
assign Ibc96fe0a6bf1f95036f97c7d44fab575 =  ~I3f0f9aab07427fa81fc3096c6b6d3d6d+ 1'b1 ;
assign I755a38220a693ba43701d30e7e9508ad =  ~I12a7983041f9c298d533bad58f41d24b+ 1'b1 ;
assign I896fb82baa9647a14f4b5b1ecfa70a15 =  ~I78503880e5c96ec0a03c75266b1226e8+ 1'b1 ;
assign I23d1c973d7a2048353fbb68e4a294c08 =  ~I8adeae445b33f634977957bb1a2259aa+ 1'b1 ;
assign If9fd1e08af14f2fd4ca363383f48580a =  ~I73bd13f381d15e0b0198b60cee44bb42+ 1'b1 ;
assign I8f3782f78d88a5c3bc93709564999b30 =  ~Ic8b651c2b043a4a6e4cd259774322230+ 1'b1 ;
assign I986d61d79ce31f4677f3293339db6ad2 =  ~I76979d7df582f9306e796a03cb540963+ 1'b1 ;
assign Ica4d93d9fad21316002008ade5106a9d =  ~If61d4585986757a525c54589ec93d8c6+ 1'b1 ;
assign If77592d5d8bed32477fd690341e543d0 =  ~I1bc5766a4a3cc2b468ab8ef62eab691c+ 1'b1 ;
assign I25b70c6b830cbfe1b41d8f289c751924 =  ~I21585169e5fceda643bd03fddf8153be+ 1'b1 ;
assign I2a5d65eeffa18dd9af9fe36463dafd7c =  ~Idb2990946f60939136b3bfddbc7b1671+ 1'b1 ;
assign Ibafa6e10bd4edf5d224fdeb2f9adbf98 =  ~Icfbf703890f684bfc96decc429deaa04+ 1'b1 ;
assign Ifc25402bd879bc5c43b4945b60cd4540 =  ~Id5bb42639a1c1c1d67df1c89a14a2bfc+ 1'b1 ;
assign Iec48da6882325d8a33e0e0e845eb18a0 =  ~I55b8ef91d667c1c1d9e58dbc86a2288a+ 1'b1 ;
assign I0fd05e46862fdf8e614afaa3fd478602 =  ~I17ff683da41b469c8c8b82ee32a7378a+ 1'b1 ;
assign I6253a59dca81842d9ab6e58cf204abbf =  ~I51f10296c38872338ec7df35ccd520d8+ 1'b1 ;
assign Ib18d64bc58b354358ee6ac16785880e2 =  ~Ia59ff33765ddf4aeb17f90a70c01d76c+ 1'b1 ;
assign I28689b693a7a5f761a1f252aa3ef3b67 =  ~Ibf97abffb1ec40f2f0e099a814e04ab2+ 1'b1 ;
assign I1a4e6d12f9776d5e61094e0b5edf71d9 =  ~I3efc3271e18a1e350473dcf3375088aa+ 1'b1 ;
assign I8e1ad23b7ac662bb827a83d3709f0adb =  ~I1efd1220ea9100f2fb4f169ceaf462a5+ 1'b1 ;
assign I000ad2287813072cc18dad933758f2ab =  ~I9af399f27c8e2b62b7f3fc6481ef9318+ 1'b1 ;
assign I7bc3698b51b89ac38ba5f4b5428a0c96 =  ~I171bb4ee9be2f92e4d82997108572426+ 1'b1 ;
assign I78aea1705621e2845a331c3e61a8055b =  ~Ib13cd76c20fcaf95f26f4914380c4fcf+ 1'b1 ;
assign I0a31314c3580f5f9e61e79c133e5d794 =  ~Iafb219f1c8c6883e01fbfb4c887c8d6a+ 1'b1 ;
assign I0e274fd7bfc0388fef95a8ceb939ee91 =  ~I94fc9b0bdd2b0a89a9f6351f1fdd4ff5+ 1'b1 ;
assign Id6f39ddcb73d3f4ec081a365d11d1ef4 =  ~Ia9ceb45f33402293c162cef4037ba007+ 1'b1 ;
assign I807770bfa86d160459d6ec3c0f4d6a0b =  ~I0fa4e12e62e8a30b3b8045143b344b4f+ 1'b1 ;
assign I31c89b8a11a3090bfd74b112cbc474bb =  ~Icec1c637d24ca277bb2e488257e92a40+ 1'b1 ;
assign I79b82cb1bfc72bd5a9d313b9e9c9203c =  ~Ie9aca08b988fad20904545fe070defd5+ 1'b1 ;
assign Ib1046ae03c9a77fd2c0b3e9838e9af87 =  ~Ie82304b2c8583f967649475e309e68fa+ 1'b1 ;
assign Ic63723fd43cbbbde51c233a3cca15d3f =  ~I60da0fb8a2c0669d5f9037ae99b23565+ 1'b1 ;
assign I3abbb59abada1aec6941185f95f738bd =  ~Id8c19a3547c17ed513d2d857adc66885+ 1'b1 ;
assign I8d5bd7039a77ce82ce0f6cbba9c2a076 =  ~Id74984743844e9495ea0f528a391f4b8+ 1'b1 ;
assign I527ad0b9382dd7b6e657dc1a32d8e472 =  ~I9edcdd5b927b3f6b3a4c7cacebeb4a82+ 1'b1 ;
assign I8de02f32e14e719f4930d99743c04a20 =  ~Ic89597a95f50382cd3a2730896735d55+ 1'b1 ;
assign I7614dd5e9628c761dd9b2a512cb1da98 =  ~Ibb7d203dfc75bf6211b09ab94877f93d+ 1'b1 ;
assign Icae7efa4742dd0ad943ee1f67b0c9b14 =  ~Id2f2e6837c83973cb2173454433acb88+ 1'b1 ;
assign Ieb1854b79e9a2bc6cf5aa1c319e8e753 =  ~I1259d5918f8d65b4b22ccfef22fe3afa+ 1'b1 ;
assign Iff50b77f300183ca59a67ccbcc9573c4 =  ~Ib84e8c6e7fd9d7762e6e7e508d5ee40a+ 1'b1 ;
assign I4868604f8178663de759d4c63dc6c4bd =  ~Ia032017912715abde99ffdf5ba732c5f+ 1'b1 ;
assign Ife992a151986c58df4cba79b6bc4ac0a =  ~I55c310bfefb635448ef9c25c5d15987e+ 1'b1 ;
assign I9ab973fb74d9fac5d78eb8fc2c7ecf36 =  ~I92c0f229cf7fdb2cc0fe4d84f4d9b11d+ 1'b1 ;
assign I5ee7916e859b86a98538659401685016 =  ~I5570eb486d238fd96f9a59b174f5a22a+ 1'b1 ;
assign I48c284cefb8cfb5a938a8f23ce4d7f03 =  ~If6f01d24acf4a8b38bdbb1b366cd9a47+ 1'b1 ;
assign I5c1fc666b77a689478654dd29519f458 =  ~Iff29fff36064aa4f9d339d4c62956e61+ 1'b1 ;
assign I38bba98b59184c75ba3b27e1dcf52182 =  ~I818d7cae6f1b80ac452dbfc073ccfe7a+ 1'b1 ;
assign I6905b65403c16b0211643227ece536f6 =  ~I77ecfe991c6ec778495d7d5e5e442eca+ 1'b1 ;
assign I3ed34401bba9d5f229bc98480aedd9a5 =  ~Ie7c6a56e8b6f7756bb5a24bdfd6a855e+ 1'b1 ;
assign Ib4d05804277cddc7f00ac17ac14f5325 =  ~I9f9bc8eb8b2978a3dc529c34516fdf75+ 1'b1 ;
assign I41babdca6d3fa462849592d37b0a7998 =  ~Ie3c0e5a4b00a92357a5d37e527d59b61+ 1'b1 ;
assign I58cfec706dc929ebfdeaca6e01b00c0a =  ~I9b9a9486420e7d4aa105c48dd50aa74d+ 1'b1 ;
assign I7efe3c5b2fc69840a79545e0399ce749 =  ~Id12199a504f7aa298fffaaedd1aacc99+ 1'b1 ;
assign I70e3eeb2b3966676d16a6aa4c85753ab =  ~I813691fd8ea36626d32c8d2562163f32+ 1'b1 ;
assign I2a32d545d1e7beecc7531174c7e8dfbc =  ~I5fd3aaddc3eb8afeb82768b45e2d53d7+ 1'b1 ;
assign Ib8fb40e4ba0ba1f5e9f5a99d1271ed06 =  ~I1ac281eab6c7459e835fe992142b7857+ 1'b1 ;
assign Ica792cb9850a61fa4a8bd8a4b6c6ca05 =  ~I49e5078c9161e8bee00fb76bc00b5288+ 1'b1 ;
assign I779e5997c66649d6d54fd7f0514c47bd =  ~Ia697adf14616bf50d6e8178596b9fa7e+ 1'b1 ;
assign I5aa578b0c2831453683fa44af1878cb8 =  ~Iff3128a26dabe63b015dc6afc98a85a9+ 1'b1 ;
assign I735d6229ef1a4ecda0a1f1dbdfb53fc1 =  ~Ifc04708ee5a7cc2b3f1850db778fa42e+ 1'b1 ;
assign I62affd47512c5e8f0979244115624d97 =  ~Ia405859c9dff67905b2e91bcbc06259e+ 1'b1 ;
assign I14fe27afb3df5531b18dc9604e8dbe65 =  ~I2fec8f62b28575e8f3af756db66fa232+ 1'b1 ;
assign Ib1b1626c84dad8ad13c058f921ffd57d =  ~I98e97c02477032ead66dc50f3f274e5a+ 1'b1 ;
assign Idf4a4bdddb88c21c5afe10a02373a6eb =  ~I9f2dc5add3a4d1e6eb3116c741cd2f82+ 1'b1 ;
assign Iadefc2a3d07ed4b2c3c46b2ab5dec252 =  ~Ie122f7d8a48d7ad29d998b6a14b8e70f+ 1'b1 ;
assign I19315957077b037ffc6415dbb06ef789 =  ~Ib5576c996062391f44066d893dd5cb91+ 1'b1 ;
assign I1f9be09334407fc86c83a7c127e17bbe =  ~If931597aab866a74c3a3ffb1cd429583+ 1'b1 ;
assign I28e17a5af7a7286a2643100d6d058dc0 =  ~I79878bd69ed53785b8a5f025a2a00a4f+ 1'b1 ;
assign Icb2297c397bfe56be251ffb6b249a020 =  ~Iefb0a20652954fc2002154ea874c120a+ 1'b1 ;
assign I64a48984527d660002f1f82c376c7a84 =  ~I646ca66e4e9f24b4fb75b38bf293b4cc+ 1'b1 ;
assign I238b5fc70ce9f05b6322a2691b3a0207 =  ~I051f0d4c44123e3637b84a32c9a00a75+ 1'b1 ;
assign I00c16e7ad3821981032a42d5baa767b3 =  ~I1876f9ec3f6f637ee40cdad7cc347f6f+ 1'b1 ;
assign I42fd5b094da200b33036e6cb8c7d0286 =  ~Ic3d6b8dbec6cf92a9b6a17fb2f75dcd4+ 1'b1 ;
assign I98b7e26a0e9ec9ad750ff87cc0641a73 =  ~I7d89f1db7b1015d34363ad781374de58+ 1'b1 ;
assign I3ec904916870171bf837e162d1030052 =  ~Ife217ec4da1f1477bce034cb3545160f+ 1'b1 ;
assign Iedb11b97900b7dd769d31f8a89521975 =  ~Idc5e5e98508c94b87a760f8eb36fad41+ 1'b1 ;
assign Id0dceec6497c9f13ada07138986d4145 =  ~I9e72b0c823f297535f13a1b3072c2776+ 1'b1 ;
assign Ibfe7d9bac29b8838f20cdcfe8ef7da0c =  ~Ia81da7c58d6636ab70e0cf3e263a12c0+ 1'b1 ;
assign I4d6c95605595942a34573d6ed55eb326 =  ~Ibfc69ef08382c79e30cfafd89bfeff69+ 1'b1 ;
assign Id6d8f32958dfa1a98958a84e7f1aed02 =  ~I2d2afa9165b7121dc8289e9e6cdab5de+ 1'b1 ;
assign I971cdf9ddd1bfff5664eec35f22da335 =  ~I065052693fd8ca87614feb60f7ef37c3+ 1'b1 ;
assign Idd8bc1412a0dc5f489ef253a6164ceea =  ~I13344a81551374f665cbc17c7e94296a+ 1'b1 ;
assign Idbeec36de0128e5924e214877c82bf11 =  ~If5a1d2de0715fa87d191ee5f48171676+ 1'b1 ;
assign I50a9cd240979bc56421bf85011ae99ed =  ~I02b256f74ee86b42ff1eba5e3d242737+ 1'b1 ;
assign I6437095f6bad2d4fb2fbe0361f60bba1 =  ~Ic113fc051eefaef846f440e98f2f8913+ 1'b1 ;
assign Ie9b6eb3bbac26635aa00c38110958d46 =  ~Iabeab9bdd0bd82dd145218b563b5dac1+ 1'b1 ;
assign I9f34e81e3ffb85539a6273babc2a732e =  ~If9ce0a09e3a4e816dda002a24319ac0b+ 1'b1 ;
assign Id0a1ab8472d704001e0eba0317b117d6 =  ~Ib5a7d72c36e41754033a64fbe0718784+ 1'b1 ;
assign I9e632217cd0561d8faa28e4b8850d995 =  ~I41df12c7dee8526abf92b8e98965fa06+ 1'b1 ;
assign Iedeb5b7b2fa8acf1ea083102678710ea =  ~I83dfbd224e7465a6fd769e407182829a+ 1'b1 ;
assign I972431d1f5af0bdf4828e4f85591e358 =  ~Ie57bba5092ec318456365b81b36aaa65+ 1'b1 ;
assign I1f41024b715d8312944ccbf70e95bb40 =  ~Ibcf043d24474ab8c1002d15fde2d7da2+ 1'b1 ;
assign Ia6bb5ca05f5d0af452c994dd50004e1d =  ~I2e3385871c6ed8cf9519f273c8a19fda+ 1'b1 ;
assign I9a1d1d1c862808f9a769cbdb3bc634e1 =  ~I664917b9f44515bf556d69ade4ca408c+ 1'b1 ;
assign I9734eb86f4e73ba217739baf5cb1b13c =  ~I28deacdec0fbd0bce49b654c2620ac38+ 1'b1 ;
assign Ifc0fe00f86569956df72d8a960337e8c =  ~Ibdfc4852c620f573f929584e6b816f35+ 1'b1 ;
assign I223341a807a1d555f759632f67815159 =  ~I5a69b2bbb63ab919ea2270503cd326f1+ 1'b1 ;
assign I6c1f5cdf5f2917118941f4af14d67fef =  ~I2eccd8d60a19481fa595566f51c7aa4e+ 1'b1 ;
assign Ie84e88fd1aa2a0b90aa1715fcd27a329 =  ~I49eb4bba42440657fe04b711eedfa67f+ 1'b1 ;
assign I558f70d7039a8bb58d8ea3f72e43dac0 =  ~I9ed8323951af0de78ae89153cbf9e9eb+ 1'b1 ;
assign I9924269ed3de12f1f2a28893c7f95292 =  ~I1d00816529836546b514f54b1275d39e+ 1'b1 ;
assign If1153befd1396be2798cc14535ddeb8a =  ~Icc58b9a24fb9ef7e8fa5f13a2cc0a0cb+ 1'b1 ;
assign I9bc447b20687fb3e7eff45792bd4dc3a =  ~I9339aef608b029175b488e82f5b3f1bb+ 1'b1 ;
assign If590520f01e452db9867a8d6d5dab29b =  ~Ibd2f24860b701ab46e0c436d774e43f9+ 1'b1 ;
assign Id93ee7d283016ab9b0aaa21237237c54 =  ~I37fe66ec8927f27f646b304500400ccf+ 1'b1 ;
assign Ic1cf03baabaed466fe532e4db3a9ea78 =  ~I4bd6a48f494cf633a857b8ccbd67af68+ 1'b1 ;
assign If3031f9aa8f6eba90eac12db7839fefd =  ~Icd7a7566438dc67e77f138ac814844f0+ 1'b1 ;
assign I0dc2708970ca2b6c092273b6626bacd6 =  ~Ic3d4239413333883dd926c7a42c0a87f+ 1'b1 ;
assign Ia58944aebf0b4f0a7d76a1444fced9de =  ~Ib8298d1ead61bc00eb31599b3087d769+ 1'b1 ;
assign Iedd8e69679d10e05f2889f1d71cf0e7b =  ~I23dbe33ce46f94d3dff1e6d391305609+ 1'b1 ;
assign I90f0d471914a2333b9dc14d6d01cf927 =  ~I138286817f424c76e8a4f30540b0530b+ 1'b1 ;
assign Idceeb22013af64b6bb9f0d773e9ffe9a =  ~I30c645a78b900306864a1ab23e923bde+ 1'b1 ;
assign If43574342e60a625fb6bee5a495e88f3 =  ~Id88681d0fe3ea62530166938503db05a+ 1'b1 ;
assign Id285f055275014d9f23d35f91879afa1 =  ~I808008402174fa4edf42783135c0c3a9+ 1'b1 ;
assign I8c803ab08db372802117de4fa4e2a187 =  ~I3ad4d02ea2e52a49b6fa4f1da9b58149+ 1'b1 ;
assign I13ba48a6b360f3cff5f37ce60cb735c6 =  ~I39486eecb7bbfecf26573a7a5876feb9+ 1'b1 ;
assign I4547cd1dad45dfd01e335e8cf20eadd6 =  ~I21e8ea20029fb2cb62103405b81b21b0+ 1'b1 ;
assign I0a305655b815b0cc159ac1c5f4ce30f8 =  ~Id0b67fa451e276889e02779ddb667904+ 1'b1 ;
assign I3633737da6b74284b0ea9a06c3f5875f =  ~Ic328d25a58ec4559b753da3bcff938de+ 1'b1 ;
assign Ia949c1b338d1cba07cf6bb6572c3e322 =  ~I49c44c2f2522e086c2db8a00647ba35c+ 1'b1 ;
assign I9a0185f8400159415bc0ad6c38284041 =  ~Id4152a04385391294f4b8a18df2cb9ee+ 1'b1 ;
assign I3eeffe43e7deed7ee77a7f5a3bce3cd2 =  ~I5b0213a3df61e94fd0b744a8141f7502+ 1'b1 ;
assign I85af0c31ca7002ae569d9f5ce39943f7 =  ~If0ad11ed403cbbed68614b01e2a3793e+ 1'b1 ;
assign I3dfb8d2fad83fbd807fbfc6330c5b857 =  ~Icfa1170bc73534bee13778bc3b88a2f7+ 1'b1 ;
assign Ic12be21bcba5fa49437cc44dd8a7f064 =  ~Ife1bd938a0dd06d8d3cf30ff41a303b2+ 1'b1 ;
assign I713a384d022d3012e3d0019f5c4ac077 =  ~I4a09cb1b99b476fa6fae0bc44c41a041+ 1'b1 ;
assign I80550019479d0323d0dd7e7d0f767d83 =  ~Ie08cf323944813e4b9e2d59a680ffe8d+ 1'b1 ;
assign Ib8a866f080dd997e0b6c93b6c844d1bc =  ~I85fc307fb52d58550eeecd33bc4207a4+ 1'b1 ;
assign Id542de206d736ee3769ea0bd037cb627 =  ~Id00dd13741fe621d0a240bdc92318f55+ 1'b1 ;
assign I77e6cdb09c92492c3303d0213de9c291 =  ~Idc8e891fd432df75a4eb133ce35ecec4+ 1'b1 ;
assign I788c33a9f94b26f4ce0f515891d06f90 =  ~I2a51cada20cbd14f7d5a289599e68b53+ 1'b1 ;
assign Iaf7074c2b570a296fe2ea8a5a7097ca0 =  ~I65a701d1e083e501544bb0fce24f0c4e+ 1'b1 ;
assign I8964c6d3f8e02866a6ad86553ab05d99 =  ~If3020a9109ac83274b5bafac18d176de+ 1'b1 ;
assign I2aa25edaca90c9dae8ed63b48d333c17 =  ~Iaa6bd55038c2ae911e4df08f707c55f5+ 1'b1 ;
assign I51a440917c7ae23339bec6f8a745c103 =  ~Id49065cedf20e13abac8971534bb8b0e+ 1'b1 ;
assign I56ce875e4619d4d8d6ca2fa0ddee91b1 =  ~I0bb64952d77b59803a561e14b950b9b1+ 1'b1 ;
assign I80607da8f92f5a5d2e4798a62a7b1c5c =  ~I01e295a6ab88c6f34b44efcc32a23233+ 1'b1 ;
assign Ic4dcaa520e26bac40b3876f02074f856 =  ~I2acf864d587b7681ca0fb6e2e2bea617+ 1'b1 ;
assign I3b2714d34081a3b6cccc47fa1638e72e =  ~Idfd0410b37713e8808f8bea81e2af881+ 1'b1 ;
assign I2db1d1ee8f546c00e512875ce2e13cee =  ~I02861f333b5adfd4962356cdf5a11f23+ 1'b1 ;
assign If80a6bb104ff3b2020e909103c104063 =  ~I4ddbc3daa65b111cb0d45e13d62cc292+ 1'b1 ;
assign Iadb72cc5444816fbd132256493930bb4 =  ~Id363d158feb8fec19b5f3d73d84f0068+ 1'b1 ;
assign I3a8ec1ad07bfada3d2c6ffca88b8b678 =  ~I8ec9b7a6e65e727abbed336ce240a4cf+ 1'b1 ;
assign I0aa042b86d9f68d22a49b4eb480a9088 =  ~I128fa1e99b7eb9b6905c2cfd26b95ab4+ 1'b1 ;
assign I89a387374771b68d87d7ff2dcc810829 =  ~I93d459b6da42a205c91c48622f0c5032+ 1'b1 ;
assign I2935b3d5c3bba4dddfc7ae03fa77b229 =  ~I1243cc8d5dddf7dd65b40c0b3b958b9e+ 1'b1 ;
assign I4e0c0248f4aa97d263d64dfec36e3aa2 =  ~I238df7e09d42bc93a972da349a00f511+ 1'b1 ;
assign Ia2871d7493b2727d2cb2fbab596b7e6a =  ~Ic658b2afdc7331653fc84d6372d47418+ 1'b1 ;
assign Ie57adae8873946d6c706074b52a49786 =  ~If39be111eb101c9c983fe0baa9a1cb18+ 1'b1 ;
assign If5ac85646e4b339a19af658f01d0a17f =  ~I9d19d5b7d8b256c1707de97a4549c458+ 1'b1 ;
assign I1c092426f34be030b3e020f40517b0e1 =  ~I6c2fffe204091f7f64aea16b0ac98769+ 1'b1 ;
assign Ic719b72ad271bc7c077067518e6bbb98 =  ~Ic4ba4d2e5c12d9f1dd233d64929f1072+ 1'b1 ;
assign Ib87362230682c88d68a0ba70e25f3c20 =  ~Ia9dec5831998d472d11429e5a7e60ed8+ 1'b1 ;
assign Ifcf097a102f8dc1f912022fed893d222 =  ~Ieaaf52c1e663f260292bc1529718d681+ 1'b1 ;
assign I56483ca3fa550dc59bfa347780cfef7b =  ~I37061896a09588a73445deed73d3746c+ 1'b1 ;
assign I4aa9f61be376458185c3235442c8fda0 =  ~I02f25b80945b6f58193fb37add3da2d8+ 1'b1 ;
assign Id91fde1007d47258273299de80721390 =  ~I19045602bb77f12666ebd44f813db2c5+ 1'b1 ;
assign Id58498c34aff2e1216c189b9df88822c =  ~I4abdc8d5318d2922696a8aaee46ffa59+ 1'b1 ;
assign Ib52e0c68caadcf4dd9636a84f5460e53 =  ~Ie139f2048f346d82623c8fc6d40c9acc+ 1'b1 ;
assign Ie19679053b289bb5a0aad570cc81bd14 =  ~I8d99c96e203fafc81d13ce5aee925d75+ 1'b1 ;
assign I8862c5ef45b723c9abf5d0ab6854a900 =  ~I37b0bdeb3cc54d6a97720c4912c67832+ 1'b1 ;
assign I30db951a07af96a8ddf59360141b9a6a =  ~I08257e9e6c74c60448e22fb9855f0825+ 1'b1 ;
assign I4855a0a0c6426d33014ce6a4c96965ce =  ~I32188cca2fc715698fc05b0fc6506434+ 1'b1 ;
assign I362e8db1791718290bd33a79b4fc0855 =  ~I88f1cbab9b8fa3802345f745d024931c+ 1'b1 ;
assign I773f0508440fb71d73fd82a372cc0a00 =  ~Idf548c0e78bd221bf9f612f27002fae0+ 1'b1 ;
assign I792891cecae468d7a87e12f2da62a718 =  ~Iedfd2e04f5740d283388639dde3ecdb5+ 1'b1 ;
assign I33303820ad094d7a0ab53bca722fc609 =  ~I7088c83eacff6f1dfb134f79d469c8f1+ 1'b1 ;
assign Iff98739de575e25104c0dc30f08912a5 =  ~I6f8431671331f4ca7ea19656e0677cd4+ 1'b1 ;
assign I1952614b64ea451e9d0646dcce5dd1cd =  ~I1e31259e267e04920cbbd16bd7aa18bc+ 1'b1 ;
assign I49c1a7d1c20a25496821ad80c7eff790 =  ~If54d9f8088e67e44cfa3026f5a520fd7+ 1'b1 ;
assign Ie2be17a55e79ca76350e033f227800de =  ~I6fd2c0746407b23aec5dff1e083f5fca+ 1'b1 ;
assign I737a5b06f848cacf0c8da4985c73c66b =  ~Ib2147a19b44d361da628a628fbfaa988+ 1'b1 ;
assign Iab160609bb21501aa55b662d2010357b =  ~Ie804d1f4b241a2de3e9d9c7c876d914a+ 1'b1 ;
assign Ief74f1a9d4a43ee5c9def7b83369bb21 =  ~I6cd1e6db57e06d8f5e60a31f48ae4809+ 1'b1 ;
assign Id144423f50751e661db3860a8487d004 =  ~I3e0e8832d5338423284ac4b2a0c5f3f5+ 1'b1 ;
assign I623352a4f6705b21d461d6b32e85c12b =  ~I6ac006d79e95e222cdc66754b67a08ed+ 1'b1 ;
assign I28d1dc8dc594977b5058b5bb9f6bfc66 =  ~I29087dda1a527842aeb3d35d66c853cb+ 1'b1 ;
assign I5371a83bf9d6f334cf8d1c5b082527e9 =  ~Ia67e5920bbac700dfee52cd96b15963e+ 1'b1 ;
assign If1605d6646fd267e701668a7245b3b44 =  ~I1f6ecd894d90547f661e7a3888d048bb+ 1'b1 ;
assign Idf5eb1ac2c5bd92fa08ed935ae298255 =  ~I3112e793c6e79e1f5da2776e69a34e3c+ 1'b1 ;
assign I44ce30330c4d2d6033a0a970dd2bdd68 =  ~I79152f32b45ed5b4a5302f6460707b01+ 1'b1 ;
assign Ic101b8f56ea1e25c6b752583a1b01242 =  ~I3d16e7d6b190639b88a217f19ac63233+ 1'b1 ;
assign Ib7cf44e681881e55d2d353280a6319d6 =  ~Ia1be780c686163cea54b62d6ede72dc6+ 1'b1 ;
assign I35690f724e964248dbb1e80fb1ea49f8 =  ~Ic398c31a2a6ca89d0236534589a5919b+ 1'b1 ;
assign I5affa2759148a6baf5b9f0cd3122348c =  ~Ie91c3202bc957b350d1915000564392f+ 1'b1 ;
assign Iaeea1f06ff0c6e9cfa43ba14420c3adc =  ~I687957f5300b0d4f50d6893cc556bf25+ 1'b1 ;
assign Iac5a23266c3b038b4b54a916dccdf3a8 =  ~I7816b368e8e8b8dd69383b2c9327120d+ 1'b1 ;
assign Icdfb7f52cc27b1cfcde90a100d29af13 =  ~I5f021f4a664205afbe0761af4c8914f1+ 1'b1 ;
assign I71484d7e00efa02a08b54a1405f2902c =  ~I69728004b59b5206a03a8e2087834f7d+ 1'b1 ;
assign I68a9b0607e69e8b3dae64689eb288a33 =  ~Ibbe1d623f8f5f3aa7fc70197acc6df5e+ 1'b1 ;
assign I2598c48aad48072a7f216b2ab56ee532 =  ~I4cb9f74288811592fd97fdff52bd6fe7+ 1'b1 ;
assign I796e3a193b1b66fa9a04ca60aee11ea1 =  ~Ibb471dbccd39d41e951e98348812e343+ 1'b1 ;
assign Ic96be7e69faf0f43b92618131cf0c98a =  ~I7f37d68f8ddcf8b4d5e99fb51eada873+ 1'b1 ;
assign I648afe4114ce435bf1d13e0ad54425cf =  ~I72ded7153883418a712ef967439d2159+ 1'b1 ;
assign If05d7e30b4717e0a1bfd20b90d0539bd =  ~Ie071e08299bff6bbdbe1f84703aaec08+ 1'b1 ;
assign I5fc356af8a62a1d739cb375fb851e90f =  ~I1b79aa38a39ccfc839260af89aa78e7a+ 1'b1 ;
assign I22f4c5403fbe33d18f97cf21786cdd80 =  ~I7384296e4190d83fb9d9a92cf965125b+ 1'b1 ;
assign I9a1b2b9f924099f1e57fa501ba2e33ba =  ~Ie03034ce6233ca24effe53a2c0c8f6f3+ 1'b1 ;
assign If6253af4ebc430e4937269a5f4989b29 =  ~Ic298f77f42fc1d41cce684790036ecfe+ 1'b1 ;
assign I0427d17423548dbb33cf792883b4be8c =  ~I805269f95afbeb6b93182f68868d08eb+ 1'b1 ;
assign Ie539faf01ae85253e399308fef98afd6 =  ~I881328804c45b06767af51e11182b27b+ 1'b1 ;
assign Iae6e7c42f250cd9223f18f8830fb177d =  ~I958993626e6e44e12f7c1e8026914680+ 1'b1 ;
assign Iff47ec1743b59d7f90e9042af7ce44cb =  ~If31528d1fc3a083ebc364e75cdd9c71f+ 1'b1 ;
assign I1cf4a55ebab332defa32d2922b885285 =  ~I4703b8d5a9033027889bfa8685e09e4f+ 1'b1 ;
assign I284913858691ad5724073b73a820047a =  ~I22d8e84d2db4b07111b7fdc6eef34cc8+ 1'b1 ;
assign I35626ca53adbbf0a3a71cc6fcf43bcb1 =  ~I8b7c6df3b5ea575caab7820c95974608+ 1'b1 ;
assign I0d74ef22d31abcec73c7c582310b1e6d =  ~Ia8aa76bccf7eb310a9356e8b7ea1609d+ 1'b1 ;
assign I15f4cf1aa0ad5ce2bda52df338e677e3 =  ~If9de547bf469b8424f1625e990f72b04+ 1'b1 ;
assign I6c5ca5e68c8844bb1617a2288b5bbc37 =  ~I27d51b2015ea9af9bc345adabdb07b6f+ 1'b1 ;
assign I44343a9491069c3c8ea4fbd6255a5a6c =  ~I93dddce2a0dc01ecb3039fac5cf04011+ 1'b1 ;
assign I1d8318b94d86e1fd28323a5e5684a37b =  ~I746da2c1d5a620eb7e749f72f0f04a06+ 1'b1 ;
assign I825e83bd88575868f4fcc9a8b8729663 =  ~I1e15f8d6fdb4ac732768d0cf73af829e+ 1'b1 ;
assign I3184a16c71cff80c8c90b40e45f114b8 =  ~Ib719e667d7ba857f4f7432a245f4a30f+ 1'b1 ;
assign Iae133550f8bad8357a73e7de1372faa3 =  ~I4c6eec4a0c46e4f5d7c9734df48a16bb+ 1'b1 ;
assign Ibccb4a43c410f698e0fff68553326a77 =  ~I95623ec1fd5516040a9492aae0fc2b70+ 1'b1 ;
assign I72dc7aa294a3af89101ea62a4223170e =  ~I69017b49c11de463fe6d881e5c96a1aa+ 1'b1 ;
assign I91eb3e70921e0b141a344bc57dfbc934 =  ~I4fb9ed32471aa614ce6923f6a2279b36+ 1'b1 ;
assign I1986f22f2269cc135c6ed28d35fb0bd1 =  ~I2f0bc217c8a39d71adc1fc45c10b81c3+ 1'b1 ;
assign Ibef24017bc71de9c002aafa7ce9a784c =  ~I0f1c6bb577ea2b8b2ab636e64378544b+ 1'b1 ;
assign Ieae3ed78fa2c45507066f4e20d96e956 =  ~I7a248af9d606c566e03977e985c280e0+ 1'b1 ;
assign I730fd25ffc7778fd4bb02d33cb3870d6 =  ~I0bf9d47bff47277de1e72518e8d88362+ 1'b1 ;
assign I9a32313f2911b797fb0848f7d97e62b9 =  ~I24b6f4f68f291dc50caf03dc902282cf+ 1'b1 ;
assign I6373e2d64fdb5dd77733b3e4bb405121 =  ~I79335b28eea15735f760b7a8b803e93a+ 1'b1 ;
assign Ib437aa67ab7c13b45d7a4d56ce9e79b8 =  ~I0b14b34b06cfa90539c2abca5639abec+ 1'b1 ;
assign I0cb5c7a759f4c75d4a675f9777f15c5f =  ~I26878777354945712f834740b17dabcb+ 1'b1 ;
assign I0ca91c1426ba14a7b47a081cb3becd19 =  ~I6cc5daed4de5950c02c0a57b993e22fc+ 1'b1 ;
assign I0737e0cc7453e328efab2277bb712ea8 =  ~I52c382d5b0c4829127c011fae402ce04+ 1'b1 ;
assign I456af863661122cc303fccb235f3c7a1 =  ~I46ea9871e867034daa2d0501038f15e0+ 1'b1 ;
assign Idc5916c4800e9f647d51c52444ab6fff =  ~Ibb8a202599550e87831647a93a14181a+ 1'b1 ;
assign I57aca70e2b8d126c120736b2606ed333 =  ~Ibb79f2ce0b6028ebb638fc6661444cf1+ 1'b1 ;
assign Ic6650a6d092b749b4498c08d69cf815e =  ~I0d0c07d65eda2eee01df9c330c0d6f4a+ 1'b1 ;
assign Ic2e3b8f91eb218650c7b9c515c7efe97 =  ~Ie6940736944bac9be609b8d58b2cb13c+ 1'b1 ;
assign I93a084aa1e6881ab8dc905dcdcdfd7ee =  ~I472a71363435cb3ec054e00f9123ae64+ 1'b1 ;
assign I8cba172573be52c5a90bd40e6f40a508 =  ~I553223e9166dcbddd1a51d0f92d68f28+ 1'b1 ;
assign I1cccfd1516af59265731121dde878116 =  ~I495309d795905a53b0a3d3daa4f1f9d0+ 1'b1 ;
assign Ia171bbefe2d20b4c058126c33ef28eb8 =  ~I21d358fd7673c4392f4e4b3d3a858b2c+ 1'b1 ;
assign I84bc44a5d53a8f66b985b70c7ec1ae7c =  ~Ia1a60175112362f015c5531f7c48b90b+ 1'b1 ;
assign I321b104ca3c818018d4b03adfe1110b9 =  ~I5644ece811bddcec04c9e3559c86109d+ 1'b1 ;
assign Ia79b8994da536c86634bf6f54a21145d =  ~I37d2f9d3f05cb90e2d45bd578299885c+ 1'b1 ;
assign I4df55ce80eec5fee295b5a0ae92bd6c8 =  ~Ie7d10f3c0f8b0add66d2cdd4435ccc88+ 1'b1 ;
assign I46593a7956590d870fe680228081a6d2 =  ~I3c37396a1cef2f9e42b8ccc126db6eda+ 1'b1 ;
assign I906e9da31de73ae45579607a014e8b54 =  ~I2f82390734079b8d289d48a6682cc624+ 1'b1 ;
assign If5dd1a1b9e3fc0e67a85da3183480aed =  ~I9061728c3163ae684e8c5aec3e807868+ 1'b1 ;
assign Iadfb1571c78c3f0c05e4ef498267df24 =  ~I672d7ecc28a788c2602aff76187aa568+ 1'b1 ;
assign Icebb43b184c2745cc9da9d01b06bc62f =  ~I660b2fe99cd0bcaac34e9540118b54bc+ 1'b1 ;
assign I6e4b0489ec7333abf2245a1b72a8923d =  ~I6aa263fc2a061d2c4059b08309f860f4+ 1'b1 ;
assign I24ac5dd30526c1d3bc7b941103a66804 =  ~If3aef2d755013d195fd44f734365d7dc+ 1'b1 ;
assign I33681b2292c086fe536dae2aec70903a =  ~I3ad2e0bbff17683824f575deff82c6bc+ 1'b1 ;
assign Ia373ca76c3b15a4148532b3822f82ba5 =  ~I5087dc4b32d29bfd7bad49026fa58a5d+ 1'b1 ;
assign I7d08adbaf66cea04be4891db610bca3f =  ~I8a7d893f3ef6d6a93ba552320d901599+ 1'b1 ;
assign Ic09ed51b20f411683a801eaad61657a3 =  ~Ic057537712e09fa794918e5cde87e084+ 1'b1 ;
assign I6a9af8c9009b5de47ebe9ee8b79d3831 =  ~I0cbab5173052c450504e3a7d15ffda52+ 1'b1 ;
assign Ife18e8a16d4437161b75a93e3dff1b5b =  ~I81ee40feb7abd0fec3faee653f778f5f+ 1'b1 ;
assign I0cde86532c8db1a32d9fbe38a40b91b8 =  ~Ia344347a85d4e6afafa2ee3487e65def+ 1'b1 ;
assign I49c8ec4cd33e6caed8ed7dab779e7ebb =  ~I038fce1597157a3d95bd9579cc2dcbc6+ 1'b1 ;
assign Idb86f95570587a0711d796aac7004c25 =  ~I546585b819c289d855cd098818792e90+ 1'b1 ;
assign I2d1373d0b18992fa46a9607a86d21520 =  ~Ibc3a6609765818327e79519f3e348494+ 1'b1 ;
assign I30f26e090ab14551cbac41883ad8a152 =  ~Id1c71a2a34f9e6239559d28fe2780907+ 1'b1 ;
assign Ib1b4e41ab25733d1d6dd54e1fe81a419 =  ~I1cd6cf5f8119d5e6b4ca40694399b1c2+ 1'b1 ;
assign I146c0d5154a6de44c0536de873904ccf =  ~I15e2a1b4356785d73e2ab5d51f1f5ec0+ 1'b1 ;
assign I8eb9d4839a478a4e28b45a549b5682a4 =  ~I803aeb29e66384bfc62744a841bcc83e+ 1'b1 ;
assign I2501ef991a59512c43693ba9d7db8571 =  ~Ib6e220dd4f54410239dd0c791d84a700+ 1'b1 ;
assign I38213f78fd4dc52f9d2c9b7b22136c1c =  ~I8a009007fec23f4d492b0da1b6b404fa+ 1'b1 ;
assign I49ce91ac152279af421bbc6c4d9b8087 =  ~I5f89adcb1ba235a74639eca119fb2655+ 1'b1 ;
assign I6a2b7bb2cb3ca2ab932c211a68dded55 =  ~I8fd2b001ff154e4760ead2df355c80da+ 1'b1 ;
assign Idaae6ba9da8754615a2c34ef859492db =  ~I581569cc2e63bc68a8466b07ca471b25+ 1'b1 ;
assign Icaca9fc70a3ec6c48c0e41f8168e2bb9 =  ~Ia9cfdea21a65b0270de42cef7ebbf822+ 1'b1 ;
assign I4f69b8ff834c7ab3194bc9390ce0f5f6 =  ~Id66a233d2e312aff939549dfa96a8cf0+ 1'b1 ;
assign I037cb596cd48c5533ed22bc32518d992 =  ~Ie479c12c25a1964c3804936d45725bdc+ 1'b1 ;
assign I94a89577951de90edc4f73b281ad7364 =  ~Ie30d8770ab7e6643fcb67463f6999125+ 1'b1 ;
assign Ib7493a1a384aebaa7999ff1fb867fc6b =  ~I4a17ff532c9341e80f7ed0626f728054+ 1'b1 ;
assign I2ceb9e423696539135c5bae5cc2d8d98 =  ~I597bc1ec224007a78c25f7eea24c2c3e+ 1'b1 ;
assign Ia6bbf236436b2ed22bbaae3b8849de6d =  ~If198ec15fcf66e97e69f88f718979c2b+ 1'b1 ;
assign I33cdaee4676d546dd5507df4704ea1f8 =  ~I6aa13ef29cf7e86ec83affca4fa11e42+ 1'b1 ;
assign Ia44daa9ddc3e4d377267333813d4675f =  ~Ide136b08f4b6211bca8cccf494a0baa5+ 1'b1 ;
assign Ie1f8fff3f43426d6bc39e45322a532ca =  ~Ieeab247764c23256749776b0a164314d+ 1'b1 ;
assign I4ee181895efc22862b6e85802a944095 =  ~I210e9ff7f4588185bd712915954543ce+ 1'b1 ;
assign I5c24ea83cabbb6be089ac084732cb9d6 =  ~I59186d5219833d6dd2e813a2910a61f5+ 1'b1 ;
assign Ifee2342449a3b3d0036ce2ecbc9ae189 =  ~I0c8b2bb61a9c3a67ac7e03e40be2b98e+ 1'b1 ;
assign I70a9a9b8f25066612a50e411ad68e6c4 =  ~Ide24c1f9033e7057262da1bc4762b840+ 1'b1 ;
assign I1870059af857c79d444bef948bb536ef =  ~I4677558b9faf190e7960cfa9b8ee00fd+ 1'b1 ;
assign Iafe61ab12e232a1090123a0f16eefaca =  ~Ie38ab94215851e531d2100b6602d5fa5+ 1'b1 ;
assign I10ca809fe9a04eaf5d7784ba69314178 =  ~I3f5119e8fac99376aa38e4765b8b0f99+ 1'b1 ;
assign I7a1bd0a115b3a1f85cb9c54840f5bf9b =  ~Ie8040301d224f78c1fd18bfe9e29e5ba+ 1'b1 ;
assign I986a564393d944d7d202414431c6d165 =  ~Ied989966cebf0d730633606c5182a249+ 1'b1 ;
assign I464042aaa60a41c7e1faf3d16eeb121d =  ~Ib8818bc4ca106ae38cacd5c20083aa08+ 1'b1 ;
assign I34b9a0bf2b6b562fb36291022ddf5179 =  ~Ibf08556fc39044222321912e84a4436b+ 1'b1 ;
assign I17dd8612b5c7f9dcc90f17e584aab2d3 =  ~I985e2740ac0f656da8f9dd973bca99e6+ 1'b1 ;
assign Id77cf7c05844d83e808a694971145261 =  ~I73012d2d9f6f237bc50bbffc199e012b+ 1'b1 ;
assign I276c1155d766437253f12b25066b84e4 =  ~Iefd0d59e58623b14437b17297fdbf4ff+ 1'b1 ;
assign Id75b386d8076893cb73baca69c3eff59 =  ~I68d2443e98f2fd3fa3baf96f98e1f4bc+ 1'b1 ;
assign If62ddbe87274965cfd83189c6666401e =  ~Ia2d1b6833cd8ed02f05281e508e4d716+ 1'b1 ;
assign I4f73a07452638a610b31e3ee52cb5639 =  ~I512e2251bef73108eb0f3e01e79ca3fb+ 1'b1 ;
assign I2a4faf3344d9bf4ee71da0be8994788a =  ~I9bf64811d14ca8b4c633342ad22669a3+ 1'b1 ;
assign I7d7ad0cbb962a47e229fe9d8406e6fe1 =  ~I45a910acd40d5b9417bdfdc50cddf241+ 1'b1 ;
assign I82988dc2dc83ac61380d2a5cb6551768 =  ~Ibbcf5c5f4528b03508b506c43e4511c4+ 1'b1 ;
assign I058c3a9848fd30010e4742d8682081ac =  ~I2b8b54048e164ef2f1c072517fdfe400+ 1'b1 ;
assign I368121c2534820a7147858c06e58b3fc =  ~Ia48d8883fe4f685477da6b4b05ecd387+ 1'b1 ;
assign I03d4541eeb1440aa72ee490c49977e32 =  ~I276395da1f3f1ae246b082408be2cb80+ 1'b1 ;
assign I75fdf5a355949a87b768b1e67db674e4 =  ~I4d0e2e01d9abf9ce839fe650abfaaddd+ 1'b1 ;
assign I088f4a0af0239602d422324549cb9799 =  ~I7e4e7909094f762c54137cbee99255e5+ 1'b1 ;
assign I787fe66b38237caf805ec14970d154c7 =  ~I761255e100d161b25645ca3a5187e82a+ 1'b1 ;
assign Icef176cff3ae503dbbe2af9ecfc4c859 =  ~Icc2ce1fa3cde69256378ec3f4a07b0fc+ 1'b1 ;
assign Ie0a66e4871bfe94f6716279ecc9ef21c =  ~Idd99afa80ca23644675d3edd60e74fe4+ 1'b1 ;
assign I474adf7a975b405c288058139a08be38 =  ~I486bcb4fb0af80c98c2ea21ac64f7a90+ 1'b1 ;
assign Iebeadb39658f41dcf8719ed413e46144 =  ~I759cca2c0003fc2c2af7709c5ebc59f7+ 1'b1 ;
assign Ie018b0d9f05a86207ae09ca2efac54e2 =  ~I1d5ce9f132cd1f46e96b511c77234e21+ 1'b1 ;
assign I51ee69807609fca0f332c8bc31afd632 =  ~I032e26ea05e88c6d325a810b67e82306+ 1'b1 ;
assign Iee1cb471704b2a8718a68ef93fd2e356 =  ~I0f72df5225a1fec2f276fd3c9138e8c3+ 1'b1 ;
assign I1731c0e3be86eec142c3732ee836e4d5 =  ~I0d18cf087b2335f1b9e1a621acd5379f+ 1'b1 ;
assign Id3b8c0ca32331f94fd98c8dae72bb15d =  ~I7684fc23c57105e856050a45640f2bfd+ 1'b1 ;
assign I6a86b0a82441c6c14436a3e0af6b0fb7 =  ~If778767ab80e59e940deeaa8a0dac99a+ 1'b1 ;
assign I8c92ff598084da7a50f7c68da96620b3 =  ~Idaf86833beb8c334f99291db9302ed29+ 1'b1 ;
assign I8bd1862e7bc2e83e9863389d532e6623 =  ~I6610e8d41cea10498d95850440ce388b+ 1'b1 ;
assign I8053269f8bd78a931878c8350693e1d6 =  ~Ibc653e701eb995e828c8180efaa122c9+ 1'b1 ;
assign I2ff66cdd7314276232715ef2361ad184 =  ~I21d36c49c9c766139b4b01df7c00a8f3+ 1'b1 ;
assign Icf541c76bfaf37fe6111de037d205f15 =  ~I0e4ffded936d7ccfc32b410aec617df8+ 1'b1 ;
assign I68319c8b9febef9f564832429c91b85a =  ~I1a5745021323efb5327d0b893962e852+ 1'b1 ;
assign I127772614218dd7c50d3136b4f174d7a =  ~I65547afdcd7fedb7b44bd51358eec4d2+ 1'b1 ;
assign Ib8d1aea4ad24c6ceb44f2cc672e1ff90 =  ~Iada3eb71e94ff6a6f4e5c702e83036ed+ 1'b1 ;
assign I9ca26c8104bf15f48b19dc3256914544 =  ~I077404a911da16d707a326f18717dc7a+ 1'b1 ;
assign Icc76d9ffc3f3d7b410205eeb8232a33b =  ~I6da1e92759c96aab8b9207a9acb244ab+ 1'b1 ;
assign I7fc4551d8a0445f79b87b4ba5f2ffeaa =  ~If7110182720ffa279b1cec1305cf9889+ 1'b1 ;
assign I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8 =  ~If0e20ea1696ff84329b9928d7f9e3381+ 1'b1 ;
assign Ie34c07af9f6adb9e4b636dce3d0682c0 =  ~I4e69ae6e73a856d4e26203fb9acf3565+ 1'b1 ;
assign Ib869a349250a765d2f8660e0dbdcf312 =  ~I64c939aa568669b4567c21be09ad0e94+ 1'b1 ;
assign I1a4fb631fdc7b5454c266589962ff5f0 =  ~Ia88eb16f68265e322509d541eb457993+ 1'b1 ;
assign I9de4e0e86e9edcf948d9eddf0401b94a =  ~I916f75e5a3858a420ab5cd4c43b13921+ 1'b1 ;
assign Iee7b4838986c962969c00a0bbe53ce0b =  ~Id076f99460a8f73a9fd43467216e8f8e+ 1'b1 ;
assign Id81b11a8ca1dd8989e36cef637ae6aab =  ~Ib4d7aeb8544fbdc36575a55b9f67f2dc+ 1'b1 ;
assign Ibe96deab015b799fe7f69bae8432952c =  ~If65d2514892fb7ee64fa4dc37fc0fed3+ 1'b1 ;
assign I986b52155cc1470299321a4933241ed7 =  ~Ibef07e48768252e9b41baf067bb1ff5d+ 1'b1 ;
assign I04be63a04f3942ce749cc9bd7540e055 =  ~Ib8fb61fa9cb8e92bc57c53a567891895+ 1'b1 ;
assign Ia7adea5b0ec86e9fcd427a5468d72b64 =  ~Id8f5f32cd0757b4d6861d17fcbd6e8d0+ 1'b1 ;
assign Ie8990d8abd23f8f9f79d7fe38c57fa8c =  ~I8be241f29e7eb258e9b3501430820b0d+ 1'b1 ;
assign I9d2f90ddddbdbb525d5f070f32546b64 =  ~Ica8a188ea43e2f28e70b8ea4e2431dc3+ 1'b1 ;
assign I905256d73bdb63bf860e15687350795f =  ~I83ceb726e57d52698b57dc39ce585897+ 1'b1 ;
assign I9adcfc18e4471209edbe9a379e996067 =  ~Ic88e7e05d83ff800b4a941ae4b424557+ 1'b1 ;
assign I3d7d048348bf833f744a9f73889b7802 =  ~I7de81aaac1e5776dfb60eed2d12d4f6d+ 1'b1 ;
assign Id619e8d4040014d0e415ff71c5e0591f =  ~I37058036bd9f4331387ee4a9348541e2+ 1'b1 ;
assign Iaf3de2ef283e03dd72002026e1299224 =  ~I570f85838c418d8501c8ccdc38a53f00+ 1'b1 ;
assign I64551529c0028ec145407be7f5dfef71 =  ~I4aa6f0c0f5163b944f11328888af73e0+ 1'b1 ;
assign I5ebe580a943b65fb16ea722ba101fd05 =  ~Ic7fc1f38ad4e9b2cb472ae75bc3c100c+ 1'b1 ;
assign I0921901599c43b27e701758026dd3ee1 =  ~Ibace8d2fba25834c83b1e57195c81086+ 1'b1 ;
assign I6033532f27c26b2d42bb3ea128f80dfa =  ~Iefc1488e3eb60b99ae08d904a15c5242+ 1'b1 ;




reg  [HAM_LEN-1:0]               HamDist_iir;
reg  [HAM_LEN-1:0]               Ib325dab091dfc3a1a269adb3ea9c75cd;
reg  [HAM_LEN-1:0]               Ifc045af19c3f10d92d2b0dfb4fbbde38;
reg  [HAM_LEN-1:0]               HamDist_iir_prod;

localparam I0c5eab3e4dfde17a8c7261f7827e941c = 50;



assign conv_Sgntin_row_00000_00000 = I5b177dd5c14ad082516b47f550875682;
assign I91679dfab57a372eddc7f9b94a231edb             = conv_qin_00000_00000;
assign conv_Sgntin_row_00000_00001 = I477326720157df2503149125a43ee987;
assign Ic2171967791a0329f3e39fc19d0a6bc8             = conv_qin_00000_00001;
assign conv_Sgntin_row_00000_00002 = I319012bc6fe93d78de57bcace0caaef5;
assign Ic7e35cf8d5cd230b94c40714f16e2418             = conv_qin_00000_00002;
assign conv_Sgntin_row_00000_00003 = I174b6c36f2af82f8047cc76543a3b4ee;
assign I679baea452c3c6d04c53baa88edd8eb3             = conv_qin_00000_00003;
assign conv_Sgntin_row_00000_00004 = I8fd5787ebf758919e7cb75d7419441e8;
assign I75a4cf2948bebc58e12bb039ed273ff2             = conv_qin_00000_00004;
assign conv_Sgntin_row_00000_00005 = I413b1c1985a6c9c6f202e85ff901e3a8;
assign I9d15f76bb68b214057566cba4b511214             = conv_qin_00000_00005;
assign conv_Sgntin_row_00000_00006 = Iea3e35ece9fdb3aff3b9ff5369e9a7e0;
assign I8be20605d26d218911e80a883a90d085             = conv_qin_00000_00006;
assign conv_Sgntin_row_00000_00007 = I30c0fcd89e0cc7c5fa348df7b4fa2ccf;
assign I08a8cd6965c23af6650568b654831b20             = conv_qin_00000_00007;
assign conv_Sgntin_row_00001_00000 = I77b05a8aa92c66a235195a66dc13c0cc;
assign I065a81ba25962785215583e7ece27661             = conv_qin_00001_00000;
assign conv_Sgntin_row_00001_00001 = I876fdba97e755b74532f7ab191fbac14;
assign I71228fe4188ab1d9796081184a422094             = conv_qin_00001_00001;
assign conv_Sgntin_row_00001_00002 = I5590d801fd7fb496019d4c31b7c6d898;
assign Ide9ef5a16d8fe32353c2c2a30e8ee3b0             = conv_qin_00001_00002;
assign conv_Sgntin_row_00001_00003 = I25f1ee9cee4d04bd8fec1fe601d016d7;
assign I0865623d3350645e63fa6e6c9b78ac57             = conv_qin_00001_00003;
assign conv_Sgntin_row_00001_00004 = Ifebcf64858d5e2d07ad7894d6182eb11;
assign Ic10356f9069e3651b9c045c906e63512             = conv_qin_00001_00004;
assign conv_Sgntin_row_00001_00005 = I163cf58b9a308e0439a8dc7c1526e6b5;
assign I43f41bf07836cee48069e9890c1de2a0             = conv_qin_00001_00005;
assign conv_Sgntin_row_00001_00006 = I3347717ba9556e69de30ce7533d4f5a4;
assign Ib8dfd9b8badef282ca00a4f793c3c868             = conv_qin_00001_00006;
assign conv_Sgntin_row_00001_00007 = I5f96a68d20e3ebc71dad4b43305baa20;
assign I2fd872df07f50688486c0d602cfc5549             = conv_qin_00001_00007;
assign conv_Sgntin_row_00002_00000 = Ie117f6ec475f5d6444998af151ce4e69;
assign Iceb7a1d4c23806b8f5824016779ad129             = conv_qin_00002_00000;
assign conv_Sgntin_row_00002_00001 = Ia538dadbd6ae3711740595a18c89b65d;
assign I7b561638da1b4a45ff59be81243e4471             = conv_qin_00002_00001;
assign conv_Sgntin_row_00002_00002 = I141cda06bae0c5666e3bc61c6fe5ad66;
assign Id50edc56fce48130247fdbc42eeff9ea             = conv_qin_00002_00002;
assign conv_Sgntin_row_00002_00003 = Ifb70a30f8bade95f402e71f95fe6644b;
assign Id13c99b7f7500c8195b54627efbc4232             = conv_qin_00002_00003;
assign conv_Sgntin_row_00002_00004 = Ie50aca688b3433fad7565998cb900155;
assign Ia92d2276a8a23521ad1b88df7c27bc2e             = conv_qin_00002_00004;
assign conv_Sgntin_row_00002_00005 = Ied33f18cbb778d5ba744d249f91c950b;
assign Ia96955d9c0a8a587e0afab37c8415d8c             = conv_qin_00002_00005;
assign conv_Sgntin_row_00002_00006 = Ibe97860165dc5d9a076ebd935385ae51;
assign Ia9b5d9ede006c56a6d83905529c77b7b             = conv_qin_00002_00006;
assign conv_Sgntin_row_00002_00007 = Ie46b71f55aef4d00168202431d47dce0;
assign Ie9ab3c88ac62369e3d92d110165a94a8             = conv_qin_00002_00007;
assign conv_Sgntin_row_00003_00000 = I92cb615e2c439914e72ce001256518e4;
assign Iea07d1adf9016a29cffd61d183e268d0             = conv_qin_00003_00000;
assign conv_Sgntin_row_00003_00001 = I7d6a6026eb3c4d06e682523424f9628f;
assign I37e6bc7aff363ed0ed1f84b23c5f3e34             = conv_qin_00003_00001;
assign conv_Sgntin_row_00003_00002 = I06ad520cb02e46d34c45f207d42a9243;
assign I47f17afcd5871fc3ac378316fd3d7ae9             = conv_qin_00003_00002;
assign conv_Sgntin_row_00003_00003 = Ifa3df8b249467cc1e827c69925ef415f;
assign I57015930f5b09a6c6b030ed01dad2177             = conv_qin_00003_00003;
assign conv_Sgntin_row_00003_00004 = I4ba41864bb1d2130c6971e0b2903027a;
assign I26a7fe395eb583258c1ac58aaaa3234a             = conv_qin_00003_00004;
assign conv_Sgntin_row_00003_00005 = Ia67f9b902a21de0414eb8dda52171991;
assign I15a1671def323cd294591564ae6ef8b1             = conv_qin_00003_00005;
assign conv_Sgntin_row_00003_00006 = Idbbf2ce4a30787c5f07c3b908a73da75;
assign Ifeaa99e03bda8ded058f98387de3d49d             = conv_qin_00003_00006;
assign conv_Sgntin_row_00003_00007 = I71d3a999d88e591e102398409b3adebf;
assign If520c1cd27f9d4bc52d0d029f693b660             = conv_qin_00003_00007;
assign conv_Sgntin_row_00004_00000 = If7f3174da35dd39af7f4792aaa649bf1;
assign I40ef50004a60ae58aedc49eb5e6797c9             = conv_qin_00004_00000;
assign conv_Sgntin_row_00004_00001 = I953b975a89adcc88039284970e9b3404;
assign If4132b39ddb92aa02d8d0346fb0e6691             = conv_qin_00004_00001;
assign conv_Sgntin_row_00004_00002 = I5a247475beb737d470f03507e55f5b24;
assign If2af8106efc1f7dd02c074af68278b3d             = conv_qin_00004_00002;
assign conv_Sgntin_row_00004_00003 = I93084ccf5b5e4efaee968b497bb2a775;
assign If8a527cc7f06a9963a80a880d225d34c             = conv_qin_00004_00003;
assign conv_Sgntin_row_00004_00004 = Ibab55499323660588ec82ebd07ab0572;
assign Ic3a431f39c678b7175ed30fde1fa6424             = conv_qin_00004_00004;
assign conv_Sgntin_row_00004_00005 = If9285bf7611bcc5ea6432215c349e021;
assign I4af080cb4e5cc525db95e5f401019e8c             = conv_qin_00004_00005;
assign conv_Sgntin_row_00004_00006 = I3566033cf5c9a06977c9182925750707;
assign Ic6386d7d8813731d612e24b715740275             = conv_qin_00004_00006;
assign conv_Sgntin_row_00004_00007 = I87b10521099179c18652c86d5887c908;
assign Ic512effb493a06ece58a2af155135004             = conv_qin_00004_00007;
assign conv_Sgntin_row_00004_00008 = I13a98f98c54b2e412cd88c96f016c41b;
assign I9b6a674dbcbfcf65f1ae0deb8fc3566d             = conv_qin_00004_00008;
assign conv_Sgntin_row_00004_00009 = I6f7a45fe64ffeda9ed120be3a4519aea;
assign Ib4bdc9069d0c08655f5e87f705943eda             = conv_qin_00004_00009;
assign conv_Sgntin_row_00005_00000 = Iad799775eb657f8973e6dfcf70a9875c;
assign If92db65b39a83e1c699e4cc6d7f9e57b             = conv_qin_00005_00000;
assign conv_Sgntin_row_00005_00001 = I5ec1e530b9007a75a778af4d82ab427b;
assign I0262b30a4efa9f1cfb11d1c3940de9e7             = conv_qin_00005_00001;
assign conv_Sgntin_row_00005_00002 = Idd59a5357d4c835379ed180ac0924bf1;
assign Ie8df350430970b5f1229cda772440f85             = conv_qin_00005_00002;
assign conv_Sgntin_row_00005_00003 = I7a626ec321bf963a5401892a7e3891c7;
assign I8070a3b7d8b1a7ae90c1a2d27aed09aa             = conv_qin_00005_00003;
assign conv_Sgntin_row_00005_00004 = I3342fe0c5d3ee5021892d53eb45bde21;
assign I39bbec42c442d1e8c818f46ad9c096a8             = conv_qin_00005_00004;
assign conv_Sgntin_row_00005_00005 = Ia858ff5551286beffd4cf82f876d30ac;
assign I9bb81dda8102b829441be46460eb8900             = conv_qin_00005_00005;
assign conv_Sgntin_row_00005_00006 = I5402fd208dc7ca81dfd2920a9cfa2715;
assign Ib23edc35fa5bbfe0415fcf0861a22d9b             = conv_qin_00005_00006;
assign conv_Sgntin_row_00005_00007 = Ic32c6734132776c290155a80025fe366;
assign I9cc16a00912e7dfc05fb505a9db23cd8             = conv_qin_00005_00007;
assign conv_Sgntin_row_00005_00008 = I5d92fdff96b9cd64f3af2b28b13e9956;
assign Iccefa45795486757515d95e5908b306a             = conv_qin_00005_00008;
assign conv_Sgntin_row_00005_00009 = I221524a69e18854f029cad30e8f94e8a;
assign Ic3a608b850709286ea0ad2f67425d9ac             = conv_qin_00005_00009;
assign conv_Sgntin_row_00006_00000 = I55e4ad2d71a29ad63b4999d64ac0dc4f;
assign I2213c1a2b831f421707a261f5a58b1b1             = conv_qin_00006_00000;
assign conv_Sgntin_row_00006_00001 = I592a495aecc800236c3470ff8e6adbb5;
assign I4636821315d702a677dc93113872e647             = conv_qin_00006_00001;
assign conv_Sgntin_row_00006_00002 = Ifdb5589982db805a0416e1c01276249a;
assign Iaf8a19fde3de660c3fa925593bebbe0c             = conv_qin_00006_00002;
assign conv_Sgntin_row_00006_00003 = I0c47ccef4b55410286248884a7249703;
assign I0052d562fb3182890c8828e52d437b11             = conv_qin_00006_00003;
assign conv_Sgntin_row_00006_00004 = Ib68deeb7bec4ca3585d1a4dcbf8793f1;
assign I21668ff77cf75570cae97f575cbcf644             = conv_qin_00006_00004;
assign conv_Sgntin_row_00006_00005 = Ia17906696bd0e095d7a5297da2e049ea;
assign Ic279867ebf3055980f3d813d5dc8dec6             = conv_qin_00006_00005;
assign conv_Sgntin_row_00006_00006 = Ic11a6b77b84c44180eb99220a0c4c9f6;
assign Ifc8c6df8904b97674f2970ebc95b523c             = conv_qin_00006_00006;
assign conv_Sgntin_row_00006_00007 = Ie08ad9bd71329858c1742c8f571a1c36;
assign Id88480a0a350bb5fcf01ed5fff0bbd4c             = conv_qin_00006_00007;
assign conv_Sgntin_row_00006_00008 = I8c0c1a0a35f4f7a688f516c567242d39;
assign If38feb4f76f761dce6145731ad235d7f             = conv_qin_00006_00008;
assign conv_Sgntin_row_00006_00009 = Ib105151d91678f81978495ff94b1e651;
assign Ieb528d666fdb708279184bb59eac25d9             = conv_qin_00006_00009;
assign conv_Sgntin_row_00007_00000 = Ie92110d19f4886cdfcfacd0920c06a4e;
assign I631a3300cb6685f47da7781940ec5d27             = conv_qin_00007_00000;
assign conv_Sgntin_row_00007_00001 = Icf3ad912aaeaa0c5cd1ab0edb898d6e8;
assign Ib54d55a70605119e37e9898b940ff636             = conv_qin_00007_00001;
assign conv_Sgntin_row_00007_00002 = I857d3155df0b6dd704514b039c66fa97;
assign I49fb0909ddf66fc0073e6400f1a07844             = conv_qin_00007_00002;
assign conv_Sgntin_row_00007_00003 = I3bc094d67805664859fdcb66f1360e64;
assign Id0eef1adba01447c14a6f005782dd9a2             = conv_qin_00007_00003;
assign conv_Sgntin_row_00007_00004 = Id14074d5230885c38b89b09b130ecf68;
assign I5a9fdec7d7ff99fe33ad6cd8afd9e059             = conv_qin_00007_00004;
assign conv_Sgntin_row_00007_00005 = Ibf312ae4f51fbc44b43848f9df62a45f;
assign I68528be9951f5b8805411711cd11ea59             = conv_qin_00007_00005;
assign conv_Sgntin_row_00007_00006 = If6ce2fa9f0b8bc74442ed8262b5089cf;
assign Ia3450e134e4086c35acbdee1e6042396             = conv_qin_00007_00006;
assign conv_Sgntin_row_00007_00007 = Ibabf61085ca7af8dfc7927b3656a76f7;
assign Ifec374bce7f5507438f550df22d61a01             = conv_qin_00007_00007;
assign conv_Sgntin_row_00007_00008 = Iebecd2d19f9174d87deedc1a273e7baa;
assign Ie87075ac979410cc11099a356966b8a2             = conv_qin_00007_00008;
assign conv_Sgntin_row_00007_00009 = I94a9de743d5bedbea3876de954f479bd;
assign If4d3b31b87c0f723241d35ce7e854eba             = conv_qin_00007_00009;
assign conv_Sgntin_row_00008_00000 = I59c5da6338f431a626c86a065a355c35;
assign Ic53b875b2ddcba11406eb2ca39354757             = conv_qin_00008_00000;
assign conv_Sgntin_row_00008_00001 = I8edf1a08ef943f06ee28771c6e140e28;
assign Ie19b39200436b0bfca13502ad36c21b9             = conv_qin_00008_00001;
assign conv_Sgntin_row_00008_00002 = I1c8024aa9d81704d2dcf63e34853f8cf;
assign I9c981b0614a29386ca5e8ebc06a17f15             = conv_qin_00008_00002;
assign conv_Sgntin_row_00008_00003 = Idc1b8aa2f81a7fbd87e4f5821d14bf01;
assign I9938397dc94002481984f5b560fadc58             = conv_qin_00008_00003;
assign conv_Sgntin_row_00008_00004 = I02812a8a833bb69eb168a1004b6fafdf;
assign I4c366a57920ff090a98a2cb8b9caa00b             = conv_qin_00008_00004;
assign conv_Sgntin_row_00008_00005 = Ic44eab478be232721e7a43d14beca32f;
assign Ieafa9d74d4a61d28ac4a913db460bf33             = conv_qin_00008_00005;
assign conv_Sgntin_row_00008_00006 = Id1dafb7e45b860d506e0c2c91b28142e;
assign Idbf9094c94c931f16fba468b9dd59a25             = conv_qin_00008_00006;
assign conv_Sgntin_row_00008_00007 = I9db50007841762c9a10f6b7e9d40f858;
assign I8d8d95ff26f33f69a182b32ccde23905             = conv_qin_00008_00007;
assign conv_Sgntin_row_00009_00000 = I36ba87b69b5b9dd919319230f697dfad;
assign I8bbe1a2ace8f51aa22cca5d9fc66f136             = conv_qin_00009_00000;
assign conv_Sgntin_row_00009_00001 = Ie7d9730b191781c78391141d95d4f8bd;
assign If0a3b88a66a816b25f17ced5d0e8f775             = conv_qin_00009_00001;
assign conv_Sgntin_row_00009_00002 = Ib774f380e3d7cfd1f5f064e93d8134b4;
assign If7e146da4f3bd255b8457fd6902005f6             = conv_qin_00009_00002;
assign conv_Sgntin_row_00009_00003 = I13b0c9578f7b6b3b7e6704d7b44079c4;
assign I89a3f8d5f760d1a650f85814cbfdc017             = conv_qin_00009_00003;
assign conv_Sgntin_row_00009_00004 = Ia01c82761aeb124cd92fb15ee367ee8b;
assign I3e0e682047f7cc36142e668828cbff1e             = conv_qin_00009_00004;
assign conv_Sgntin_row_00009_00005 = I2db290170ddae8dc52ce07edaf48b365;
assign I596ad7e132f272cb196b74faa8c75aa4             = conv_qin_00009_00005;
assign conv_Sgntin_row_00009_00006 = Ied764ee7730ad129b6f62837ef50774a;
assign I5267fa34449e6eebe891017fc32d0749             = conv_qin_00009_00006;
assign conv_Sgntin_row_00009_00007 = Idc5dd6caa4ed17a63746d30d381a944e;
assign I2dc64c3b06588542b027f997437bee63             = conv_qin_00009_00007;
assign conv_Sgntin_row_00010_00000 = I719a892ad54e63b217c7271741b29cc5;
assign I753f92da60980736440aba814a156f1e             = conv_qin_00010_00000;
assign conv_Sgntin_row_00010_00001 = Ia0c192e590d8c914555b434ce5a634a8;
assign I733605337bf6972630c089d32fd7f98f             = conv_qin_00010_00001;
assign conv_Sgntin_row_00010_00002 = If2b40d249c531e10cc22d1335f350441;
assign Iba70e737d52e6812a67c159520e5192f             = conv_qin_00010_00002;
assign conv_Sgntin_row_00010_00003 = Ibe7e5c2cb9c50eca34a3859d13e83a92;
assign I7d77ac9b64b2e8cae21c6e36947e3ca2             = conv_qin_00010_00003;
assign conv_Sgntin_row_00010_00004 = If0970d9f7b053fce3ced3521b4885588;
assign Icd0622a90782b9c451950e7ab0399567             = conv_qin_00010_00004;
assign conv_Sgntin_row_00010_00005 = I777ee54ff20d0544af18ad8a870d6915;
assign I1487170cb1f3370ad45efc801cefc8ab             = conv_qin_00010_00005;
assign conv_Sgntin_row_00010_00006 = I4edd64d1f1da865b1eb886e22726a033;
assign Ic3ff7ce12c836bf0693252b9a7a7cfe8             = conv_qin_00010_00006;
assign conv_Sgntin_row_00010_00007 = I4dbabfd592b74aef93b819163130ef5e;
assign Ib23d889edb5a6d9f27de977d3b1a2616             = conv_qin_00010_00007;
assign conv_Sgntin_row_00011_00000 = Ifb064c69c7110c014593149ae69c75fb;
assign I8f2986bc015fcc64ac5e5395ac6dd851             = conv_qin_00011_00000;
assign conv_Sgntin_row_00011_00001 = I2c741a5fed7d88e9bdd6b7459feac649;
assign I7d5041a6796c00188f74936d283defe6             = conv_qin_00011_00001;
assign conv_Sgntin_row_00011_00002 = I8a9e516aa824260998d10db758642bb0;
assign I7a2e79d42779ad235bca6ce3757cf588             = conv_qin_00011_00002;
assign conv_Sgntin_row_00011_00003 = I8bb5522183b65583fda83067990b3e94;
assign Icd1da43a4d95230e79dbd35a7ae41066             = conv_qin_00011_00003;
assign conv_Sgntin_row_00011_00004 = Ib0001d7298ad1f3b1c7603173a70d8b5;
assign I5a0f27df5158309f32f0df31e8ae3ae3             = conv_qin_00011_00004;
assign conv_Sgntin_row_00011_00005 = Ibc9a860879ccc58c815b9f6caa23320a;
assign I4255ac1af4367c321567c4e46b06ab25             = conv_qin_00011_00005;
assign conv_Sgntin_row_00011_00006 = I17c9d8f658dd6b2916b645d103f4702a;
assign I72369dedfe36cb22269033cc305b730c             = conv_qin_00011_00006;
assign conv_Sgntin_row_00011_00007 = Iba283e99a57d0a3b78ad2e309c316b65;
assign Ie65a0634454381e24bb3223a333e3ad0             = conv_qin_00011_00007;
assign conv_Sgntin_row_00012_00000 = Ic98c8641d2022080297c54ff2539e75d;
assign Idcb1d8bbdeaed6768c2a418c3048e6ee             = conv_qin_00012_00000;
assign conv_Sgntin_row_00012_00001 = Ia9c273b32d0701c7f185ab2de9e57829;
assign If3e5161254eb9056914c46263b865c10             = conv_qin_00012_00001;
assign conv_Sgntin_row_00012_00002 = Ibf5c141c5cc0a6a20c05b52bf8282476;
assign Ic1faed76fca5a9ceb7db26c2f43623d9             = conv_qin_00012_00002;
assign conv_Sgntin_row_00012_00003 = I2518ccf385b3b677d95983bc550282e8;
assign I1d1a7c5928982c278d068ebd262254da             = conv_qin_00012_00003;
assign conv_Sgntin_row_00012_00004 = I86fefad34d3c864dd0e725133f303b4f;
assign I47b1695a74e4d27389b97543415dcc67             = conv_qin_00012_00004;
assign conv_Sgntin_row_00012_00005 = I180d4f3b23b518271d7cb8189fbeadc5;
assign I5c05da8a222ad5effb9815cbf3ec25f3             = conv_qin_00012_00005;
assign conv_Sgntin_row_00012_00006 = Ic7ebdc317c978eb275eca41d5b9106a5;
assign I6493b3c087d4685a6b3f98c73dc2ff49             = conv_qin_00012_00006;
assign conv_Sgntin_row_00012_00007 = I84057a3b319ab3d6a2ed8f2310f970fc;
assign I2c72248cbe49ec0a0febac2437b8a6dc             = conv_qin_00012_00007;
assign conv_Sgntin_row_00012_00008 = Ifab075b1437495268b6a3be4cb022e71;
assign I6fd1b4395af175eff85b3bfeef4c329b             = conv_qin_00012_00008;
assign conv_Sgntin_row_00012_00009 = I89c5af1a6176cefa1f77ee69996473cb;
assign I2508854bcbab37bd09c9465c377c06aa             = conv_qin_00012_00009;
assign conv_Sgntin_row_00013_00000 = I17a6511072c7fb4846be5844decf17d6;
assign Iba7608ee0a01af103e022bcaf564bf6b             = conv_qin_00013_00000;
assign conv_Sgntin_row_00013_00001 = I9d18ff3465afd8cae63abba68487542e;
assign Ia9642d79bb50567348083b4435c7d66d             = conv_qin_00013_00001;
assign conv_Sgntin_row_00013_00002 = I1e77fe6aeaba852aba34ed37dd53add6;
assign Ice9079fb6e08d629f8c0c9ce332c8f11             = conv_qin_00013_00002;
assign conv_Sgntin_row_00013_00003 = Id38852415486e6989b89a0d85ad6771b;
assign I39ff4663007dbc89b403f3b08a69bb6c             = conv_qin_00013_00003;
assign conv_Sgntin_row_00013_00004 = I89af7644c48a80d7d22f50b008d35841;
assign Ib01cfd833a63500e03333f263805db3d             = conv_qin_00013_00004;
assign conv_Sgntin_row_00013_00005 = Icfc03646b36b971b9fa57d04a26dbfc4;
assign I0f034a8f077b0ab231727b6298e366d8             = conv_qin_00013_00005;
assign conv_Sgntin_row_00013_00006 = I05e739fc87e962848f265e2c73338cac;
assign I17d9e19854cef197fd3267618617efc3             = conv_qin_00013_00006;
assign conv_Sgntin_row_00013_00007 = I624958486d181501c7a8ec2642cb503c;
assign Iacf9640cbf486411d6ceb8fe1a2fd5c9             = conv_qin_00013_00007;
assign conv_Sgntin_row_00013_00008 = Idd775d9fe6fa8dbdbfb07d4071b9caa5;
assign Idc629414f6d0236ce0714cfaae23f065             = conv_qin_00013_00008;
assign conv_Sgntin_row_00013_00009 = I17086dc5193aa55e5c6f56ecd365cc00;
assign Id92a37c091100e9df08e24498ecb4022             = conv_qin_00013_00009;
assign conv_Sgntin_row_00014_00000 = I7e12ad8a8ef857e02f4563b2f3a7f0ca;
assign If6657f90c84ca5e2ba08ec705f34be03             = conv_qin_00014_00000;
assign conv_Sgntin_row_00014_00001 = Ibb35bace971548c9fc98d773d1aff712;
assign Ic51bb9184dfd103703cd0c6ad6edff4b             = conv_qin_00014_00001;
assign conv_Sgntin_row_00014_00002 = I68b585571699a57bc6ba5e8955467119;
assign I4378d139db4b710e3587aa72df22b70d             = conv_qin_00014_00002;
assign conv_Sgntin_row_00014_00003 = If76f04fe0baf171d7df2c0cd849aea2b;
assign Ie88285ce2b9c71de02ebd62e8f44ca72             = conv_qin_00014_00003;
assign conv_Sgntin_row_00014_00004 = I5134b762ac428bed07ce102d8927a418;
assign I88f1b5c12759a5efb2d2ded8483c9ed2             = conv_qin_00014_00004;
assign conv_Sgntin_row_00014_00005 = Id277f5f05551eeb5dec1701056330da1;
assign I6fc8044eb226a14ff1a786ddc96d2414             = conv_qin_00014_00005;
assign conv_Sgntin_row_00014_00006 = Ie886c5effc85f1fe0b6411db4a2cde77;
assign I14cf5d43fc9864820a8a25efcc5c6d86             = conv_qin_00014_00006;
assign conv_Sgntin_row_00014_00007 = I3c10d579f80bd0106506ad047d75f188;
assign I1d9b9ff357667a362f0442f19986f451             = conv_qin_00014_00007;
assign conv_Sgntin_row_00014_00008 = Id18c5a1d4eaa73a94e699e5f9e3c3d35;
assign Id88568dd34fbee42c9cb8cc15ac5c31d             = conv_qin_00014_00008;
assign conv_Sgntin_row_00014_00009 = I9ece87047aec25abc02a5eea72f0e647;
assign Ifaff9dd032cf96487be819c59b03000a             = conv_qin_00014_00009;
assign conv_Sgntin_row_00015_00000 = I12f2f886517647044cc251861721bbb9;
assign I0374ada4fe50717f2158468b7ad205d4             = conv_qin_00015_00000;
assign conv_Sgntin_row_00015_00001 = I27e1d2e0e980216b27b90ea48c061025;
assign Iee6f2484a381bd42e441ff072ec582e4             = conv_qin_00015_00001;
assign conv_Sgntin_row_00015_00002 = I41eff06fe1dea8be4613945de596d3ca;
assign Ifae345c79662c3df3dff0fe68ad68746             = conv_qin_00015_00002;
assign conv_Sgntin_row_00015_00003 = I94e4041b482064334fd0ed92b91bde89;
assign I1eedecb1d8ff505c75be7787199afada             = conv_qin_00015_00003;
assign conv_Sgntin_row_00015_00004 = Ida3d808d100e0bba290f96ed9e744e65;
assign Ie48be9e6b6fd63baa104d0a6a4561a1a             = conv_qin_00015_00004;
assign conv_Sgntin_row_00015_00005 = I4c66570630a650fa7b9bec543f685487;
assign I8eef6ca0a61a21882ea28b3d63735228             = conv_qin_00015_00005;
assign conv_Sgntin_row_00015_00006 = Ib1a40247057324b0bd810c844bf11f51;
assign I99fb9030e8361e57818c07511479a9b8             = conv_qin_00015_00006;
assign conv_Sgntin_row_00015_00007 = Iddc5b5b4501f9f13bcaf22081e5a70f4;
assign Ief67e897e57b96e2ec200e82bbc7caeb             = conv_qin_00015_00007;
assign conv_Sgntin_row_00015_00008 = Ia71cf07b645c58cffe33be1a9a960eb2;
assign Ia445bdc7def7d8c1eec31ab892c25c41             = conv_qin_00015_00008;
assign conv_Sgntin_row_00015_00009 = Ifba3e46933049cb093d2c1809f3a8a3e;
assign Iad166146f7df5e8068fc6efe4d3e4141             = conv_qin_00015_00009;
assign conv_Sgntin_row_00016_00000 = I4acf6d84471cd237f65c9b2391b7a20c;
assign I4ac79b67a8904b95f7912d24af420585             = conv_qin_00016_00000;
assign conv_Sgntin_row_00016_00001 = I17b3a9df6752da6cc987e902e6bbad48;
assign I60ec7459bbe99fce295406bee1f2af46             = conv_qin_00016_00001;
assign conv_Sgntin_row_00016_00002 = I168afc1863f909dbcb6a9230db9f3e00;
assign I6fab46b1766878b26b53f352fee98223             = conv_qin_00016_00002;
assign conv_Sgntin_row_00016_00003 = I989dda9add29306d7b3c0f376822763a;
assign I36ca732e811d67cd742d24fd4cae887b             = conv_qin_00016_00003;
assign conv_Sgntin_row_00017_00000 = I7f7b30f2acbb8e31f50b58096b738254;
assign I355725a804e0df68b4acf96ca98f2448             = conv_qin_00017_00000;
assign conv_Sgntin_row_00017_00001 = I615053b36a1851a06125e2ed5ec7f880;
assign I357137b41bb91e0659b1ac6ead9b5c12             = conv_qin_00017_00001;
assign conv_Sgntin_row_00017_00002 = I9890f7fc708c7b8cf460849b4a30025b;
assign Ie3a336de822ac7baf8486b1618ef1126             = conv_qin_00017_00002;
assign conv_Sgntin_row_00017_00003 = Ibc929201e2eeb3e61cc8f0acbade497a;
assign I354fdd241d5d07f0d8380fe8924e0a8c             = conv_qin_00017_00003;
assign conv_Sgntin_row_00018_00000 = Ia098bbeda8b755ece6b88eac83d03e55;
assign I634484f00590216c0f74f975c9c83400             = conv_qin_00018_00000;
assign conv_Sgntin_row_00018_00001 = I87f34821cd0b58f8855b25c75f2dd32d;
assign Ia89da2f1890524ad3519ab403dd0686c             = conv_qin_00018_00001;
assign conv_Sgntin_row_00018_00002 = Iab2f643f81921ed8464e1bbd9fa8c68e;
assign Ib1357cb20f471f1670ac2448f964f8eb             = conv_qin_00018_00002;
assign conv_Sgntin_row_00018_00003 = Ib0dfbbbca2d3d264065f73b4241caed5;
assign Id38b705f5d2863a020a475ffffc8afd6             = conv_qin_00018_00003;
assign conv_Sgntin_row_00019_00000 = Id20e72ac258d1d1b6cdca1e6c9e3596d;
assign I38c3e3e136acb79c8a0ff850bcc55f16             = conv_qin_00019_00000;
assign conv_Sgntin_row_00019_00001 = I5ebc3047985651f4b9a957d502a97e95;
assign Iedbe9d0e48bd36064f59faea51afddb9             = conv_qin_00019_00001;
assign conv_Sgntin_row_00019_00002 = I53222c82827cab7c770e057ae91bc10e;
assign I6359856a1843d8c8b65dc478bccb3acd             = conv_qin_00019_00002;
assign conv_Sgntin_row_00019_00003 = I339786aa60d4c71d12c65db27ac420fe;
assign Id6e5d67e7bb7c4b999459374ea80459a             = conv_qin_00019_00003;
assign conv_Sgntin_row_00020_00000 = I7a387a1f887c32e9d0f8e89912a8618c;
assign Iad44c932cfa5c249c5e59f8c706173a8             = conv_qin_00020_00000;
assign conv_Sgntin_row_00020_00001 = Ifa09fc1b009d073d5a9973b430c63469;
assign Ic3871325d57b310c95ca02fcaca529eb             = conv_qin_00020_00001;
assign conv_Sgntin_row_00020_00002 = Ia9c8cc5e3becf3d48feedec8fa2c93a4;
assign Ica1997c6c569c1d1f45224fbaa4e6b59             = conv_qin_00020_00002;
assign conv_Sgntin_row_00020_00003 = I4f134c0669b5a6a8c7e03be7eee30c6c;
assign If9c12f8662333fb54a45cfa1bc5da487             = conv_qin_00020_00003;
assign conv_Sgntin_row_00020_00004 = I1c4b29e48d0effac4839037ae5688334;
assign Ieaf14683f40374c4531326d228cb43c3             = conv_qin_00020_00004;
assign conv_Sgntin_row_00020_00005 = I3ade020bbdf8f954821f737439513043;
assign I05341013abd4206eb66fcddfd63bfe26             = conv_qin_00020_00005;
assign conv_Sgntin_row_00021_00000 = Iefe4099ff7e457f6b9fefc83e176c1a0;
assign I78212ae965ab2dcb2eed0b060d6b253f             = conv_qin_00021_00000;
assign conv_Sgntin_row_00021_00001 = I487496233a32f657171b3789590d0522;
assign I29ab844f80c105d247c5c15faa35863c             = conv_qin_00021_00001;
assign conv_Sgntin_row_00021_00002 = I39d3bce4060032a81e6b6a1c1805cfe8;
assign I7ef544597a185b1de63b4ffc4a1d44c2             = conv_qin_00021_00002;
assign conv_Sgntin_row_00021_00003 = I9963d0b24763ed8038b1f3922b8f9548;
assign I27fd0073dbcdee599fbe85cf48806efc             = conv_qin_00021_00003;
assign conv_Sgntin_row_00021_00004 = I5e69e930a318dcb0594a823b3129d650;
assign I5fc3c26d6c5aa893dfd5caa0f677233a             = conv_qin_00021_00004;
assign conv_Sgntin_row_00021_00005 = Ia50526cd3a3174bebc5a7a0889fda661;
assign I15da71a21f5842cb65b543d9bc3e267b             = conv_qin_00021_00005;
assign conv_Sgntin_row_00022_00000 = Ie7470dd75b54d14038de19e4d3043ba9;
assign Ib3b1db2d8b669988c887ed780e439b26             = conv_qin_00022_00000;
assign conv_Sgntin_row_00022_00001 = Ifbc6aa14cd448bbe416897a3671ba857;
assign I5d70bc64cf7b3d3ef4180e082e533237             = conv_qin_00022_00001;
assign conv_Sgntin_row_00022_00002 = I7547c56b32513ad45d775b4502596d9d;
assign I6354a0e638340378124e4df7f3d145b8             = conv_qin_00022_00002;
assign conv_Sgntin_row_00022_00003 = If10f33385e236eaba56cbab8c2883399;
assign I438522d92cce6f7010246424746ca255             = conv_qin_00022_00003;
assign conv_Sgntin_row_00022_00004 = I17d7f36fdade16dbcf621fe302bd7e57;
assign Iab953a8974a1eb619dc0f074c003b5f9             = conv_qin_00022_00004;
assign conv_Sgntin_row_00022_00005 = Ie9f37dba0791359bc426a73639ce33ad;
assign Iccf255fb3422c558465e45226068a16d             = conv_qin_00022_00005;
assign conv_Sgntin_row_00023_00000 = Ifc34f5d6b7a7d0533439794958959856;
assign I35b2c7e9cdc53a98913e1c16a3a47b37             = conv_qin_00023_00000;
assign conv_Sgntin_row_00023_00001 = I87211ac14d832ad3205d47fb83cf256a;
assign Ie33a780b0221084898c9fc5b237b244a             = conv_qin_00023_00001;
assign conv_Sgntin_row_00023_00002 = I17cf58ef5326978c62c03c56090a299f;
assign I9590eb28a81c730b83b92ef7653e71a1             = conv_qin_00023_00002;
assign conv_Sgntin_row_00023_00003 = Id79636d195efff260c430978f0bcee9c;
assign Ib8bf21f32c0e8b9cfa42a53807bfe3a3             = conv_qin_00023_00003;
assign conv_Sgntin_row_00023_00004 = I8015717cd36aabbf2cf4aa3a5c234690;
assign If6f3d91c3c7a43622b9a522492cd83d3             = conv_qin_00023_00004;
assign conv_Sgntin_row_00023_00005 = I9518532a8617fc8290eb6a5e981dea94;
assign I1c2674b2e6b269ed539827412c5199a5             = conv_qin_00023_00005;
assign conv_Sgntin_row_00024_00000 = Ib862ac63c230ccde7fae0e62f9d047fe;
assign I10f14b6433498e3b9e9bf021b60115e8             = conv_qin_00024_00000;
assign conv_Sgntin_row_00024_00001 = I013d84bfd582acc7accf07ec522961fa;
assign I0236c912c6d684bf4862b725be9d5951             = conv_qin_00024_00001;
assign conv_Sgntin_row_00024_00002 = I7cb58e4c486e683faa4acad4756815d5;
assign I92496f68b44a94565af28a2c28d6fbae             = conv_qin_00024_00002;
assign conv_Sgntin_row_00024_00003 = I67d57e38df8cb35ca686ac2eb44e233e;
assign I964e17c41a134c080e9c43412a514f3f             = conv_qin_00024_00003;
assign conv_Sgntin_row_00024_00004 = Ic0c13c9a929c8c46e8702cef74de8955;
assign Id023a6298e65da1f4da3831f5136afc2             = conv_qin_00024_00004;
assign conv_Sgntin_row_00024_00005 = If66524125bfde5aa48ac70c4e448b38f;
assign I6a3f405bb4a0c4448d9b9d3dd95d036c             = conv_qin_00024_00005;
assign conv_Sgntin_row_00025_00000 = Icddb43f9b760a4597a0bb637fb405616;
assign I0b56aa7a1b7549c91dddd3a06ecbaacf             = conv_qin_00025_00000;
assign conv_Sgntin_row_00025_00001 = Ie41ca18c7d11a47e274f9c33f75393ec;
assign I2ba1acca919bddcc22a41a28d43a4e3e             = conv_qin_00025_00001;
assign conv_Sgntin_row_00025_00002 = Idbf4ad11ab2a27044193448c8739fec6;
assign I7208256bb198bfce1be71390b01bc028             = conv_qin_00025_00002;
assign conv_Sgntin_row_00025_00003 = I04864c28351edb33b61a103add6fb875;
assign I9015033ab0caf3fa41dae4de43f24a82             = conv_qin_00025_00003;
assign conv_Sgntin_row_00025_00004 = I431fc2e9533012c8571d8158d4777dea;
assign I5149125aaaad943d891df6a3c2be93a0             = conv_qin_00025_00004;
assign conv_Sgntin_row_00025_00005 = Ic3ec6375998b05a3e48f6c5fe7b3910b;
assign Ib528bb7a64cce4f694081d151fa6fa86             = conv_qin_00025_00005;
assign conv_Sgntin_row_00026_00000 = Ie95662d4faf6b5a4cd5ecfa41697b983;
assign I735db8b0ee0ec98e4cce0030b11508da             = conv_qin_00026_00000;
assign conv_Sgntin_row_00026_00001 = If3b77c41fabcdb283f2c6fdacaa5e9a4;
assign Iaf08bcaaeb15bb0c971432f7f8b16d0a             = conv_qin_00026_00001;
assign conv_Sgntin_row_00026_00002 = I6c765e677f42fe600b848698c8a78349;
assign Ie1681d905517daafcc7584725cd6014c             = conv_qin_00026_00002;
assign conv_Sgntin_row_00026_00003 = Ieca2767ac27170058499d83016447aa7;
assign Ice73589836da9028def6efb24a04dbbd             = conv_qin_00026_00003;
assign conv_Sgntin_row_00026_00004 = I403303228c0df825f67436f4a7e64061;
assign Ie22b94121b58f17af14c75bfb27f96dd             = conv_qin_00026_00004;
assign conv_Sgntin_row_00026_00005 = I0ac421af6e311b6005c3e02e93ff94ce;
assign Iaa40bd3abf668a21e0f87c7bda7b3f69             = conv_qin_00026_00005;
assign conv_Sgntin_row_00027_00000 = I849ee5d34760be03d4285185136aa52e;
assign Ib1a2b31d49ae476e2f1fb9acba2d5af0             = conv_qin_00027_00000;
assign conv_Sgntin_row_00027_00001 = Ifb422c30663eb4824caa72326b238df6;
assign Iadeedf3870f0b1eae98d0f7dbbeff04a             = conv_qin_00027_00001;
assign conv_Sgntin_row_00027_00002 = Ia98de3691917dfb63bebdc3f8655c8be;
assign Iaee6d725a8b2653eeac6d5acb91f8f36             = conv_qin_00027_00002;
assign conv_Sgntin_row_00027_00003 = I67f87fbb746dd937fffc534c596f36c4;
assign Ide604e9bbe35cb55892a4602e18b2527             = conv_qin_00027_00003;
assign conv_Sgntin_row_00027_00004 = I23afd747ecece714e32fbb896b5c022a;
assign I6e37582849c2c98fd15ad92d22c222da             = conv_qin_00027_00004;
assign conv_Sgntin_row_00027_00005 = Ib9db80f43718305a8a8774d8d80c86c9;
assign I919d36a7f6ad42c4bbc23222beb73106             = conv_qin_00027_00005;
assign conv_Sgntin_row_00028_00000 = Ie6212a29c7c6b035cfff4c869f945b68;
assign I42f9b1f8ef24ad56c10086852678b456             = conv_qin_00028_00000;
assign conv_Sgntin_row_00028_00001 = I41ab6fb6ec6ef7ffff70e50f25f217b6;
assign I70ae07db9b44d530be220f06401d3d3d             = conv_qin_00028_00001;
assign conv_Sgntin_row_00028_00002 = I0bce960fcc58938e6a1e01b912eabbf2;
assign I4afdeba4fc2a12a6cbe3567a519367fc             = conv_qin_00028_00002;
assign conv_Sgntin_row_00028_00003 = Ief72606c77113ae37845e4aa4a2ae5e7;
assign I770dff588ee1f52f58bea1921cb23383             = conv_qin_00028_00003;
assign conv_Sgntin_row_00028_00004 = I5ede62333e0f7ddc5446b653ba9a2382;
assign I140078292f7209eccacd53a8bab18016             = conv_qin_00028_00004;
assign conv_Sgntin_row_00028_00005 = I3b775b06b5d78fcd7373c966a62f44ad;
assign I648d2a279dd1f587b1e45eeb35f2fa90             = conv_qin_00028_00005;
assign conv_Sgntin_row_00029_00000 = Ie34534dfd435b3d1cf35e82ca71e83ba;
assign I856fa68463aa5ef1ae53442699d38b33             = conv_qin_00029_00000;
assign conv_Sgntin_row_00029_00001 = I0ec27b590ee6dcdd9c1086105e3b6c23;
assign I6f3be51d69b2b64a04e55b8946d5dd56             = conv_qin_00029_00001;
assign conv_Sgntin_row_00029_00002 = I452e51cca9acec44e36e4efd21b43034;
assign I66528f43f614f0edb715564eba3c77c1             = conv_qin_00029_00002;
assign conv_Sgntin_row_00029_00003 = I946246be5b4745508b7d4b578f83aaa2;
assign I0d9f8c99194d9d6e187b4ad02fcce8b4             = conv_qin_00029_00003;
assign conv_Sgntin_row_00029_00004 = Ib2fe0f68044c11f879e512a200f8099e;
assign I74a4b9365391fd20c34588002ad40547             = conv_qin_00029_00004;
assign conv_Sgntin_row_00029_00005 = If2372a5956f21f97eeb9c76281b6675e;
assign I194a64bef92ecf6714141eaa5d41c9d4             = conv_qin_00029_00005;
assign conv_Sgntin_row_00030_00000 = Ie596289582a73e37f78f4ca4cab21e3c;
assign I7d9ad929660cd212387d893266b681da             = conv_qin_00030_00000;
assign conv_Sgntin_row_00030_00001 = I7b80b4902fe98c10dd72c9eb082346e5;
assign I62d8efd4227cb3dc88aa08b6585fafc8             = conv_qin_00030_00001;
assign conv_Sgntin_row_00030_00002 = I3051f561a5e1131ebf167cb6ccb5adf4;
assign I49f2a06ceb3a59773c65b19f54ff362b             = conv_qin_00030_00002;
assign conv_Sgntin_row_00030_00003 = I388528eaf83566cc56b23485a9c05962;
assign If004de0cac6e5f7701a1fce48c6936d5             = conv_qin_00030_00003;
assign conv_Sgntin_row_00030_00004 = I3ed6426fbdba8aaf1c948cca7442b3a6;
assign I028ce03be0618b816e0ecdf43d4cd6e6             = conv_qin_00030_00004;
assign conv_Sgntin_row_00030_00005 = I7b32c2b108e24750e2a24785668af3ea;
assign Id332e7f482524adeac7f7cdafcf5ca46             = conv_qin_00030_00005;
assign conv_Sgntin_row_00031_00000 = Ib81431cfb3b281555fa7e5b4582a2524;
assign Iabbd1668e0014df518ede5216232834c             = conv_qin_00031_00000;
assign conv_Sgntin_row_00031_00001 = Ie5373b01a92f2ff85be8077cfef2175a;
assign Idcb37cfc357cc088c775409fb9225b51             = conv_qin_00031_00001;
assign conv_Sgntin_row_00031_00002 = I284b23051c85300c2a1e3afe8f25e99e;
assign I2ff3edcdb6158f1e3c9a555aeefc0850             = conv_qin_00031_00002;
assign conv_Sgntin_row_00031_00003 = I71d7f72d83b7410de31e09ea96adb95c;
assign I6b24690f394792edb0d82b3b9e110851             = conv_qin_00031_00003;
assign conv_Sgntin_row_00031_00004 = I4af3e2bf2ebc913ac902b48da672c5b6;
assign I63e45abd4d27219bddcef06108b72021             = conv_qin_00031_00004;
assign conv_Sgntin_row_00031_00005 = I8ec99197a7d823f5745d382c10161430;
assign I226383d68f89db716cfd8d08b837865a             = conv_qin_00031_00005;
assign conv_Sgntin_row_00032_00000 = Ia3559d98eb372b7307f30ad1f7c4c7cd;
assign Ic72f41f9bbf470aee3c9b9b8787b31c3             = conv_qin_00032_00000;
assign conv_Sgntin_row_00032_00001 = I0e8679271ba733bb87c44b6b9f0b6ed2;
assign Ic3d00a27f15f8983a120395082854d6b             = conv_qin_00032_00001;
assign conv_Sgntin_row_00032_00002 = Ia7c9c24f8e993526e76c6915e56908c4;
assign I19bba6a58ad3ef959b33701f82761984             = conv_qin_00032_00002;
assign conv_Sgntin_row_00032_00003 = Ib895fec0b3756932b85962c1d129a03e;
assign I2bdf5d319ba9089a4da34b108f5c5ae5             = conv_qin_00032_00003;
assign conv_Sgntin_row_00033_00000 = I8f1a8a22637d37c3692e808d5eb3d543;
assign I96008f47b9f134c9c4274cfcfb28e550             = conv_qin_00033_00000;
assign conv_Sgntin_row_00033_00001 = Ifad8c7bacf72583f91be27fbe5b7a1e1;
assign I34be4b353cf75603301372840c2f91c2             = conv_qin_00033_00001;
assign conv_Sgntin_row_00033_00002 = I384e50fa8daa639124f083dda56fac00;
assign Iec71fe7fcebccf1ae0d10a5d187fcc44             = conv_qin_00033_00002;
assign conv_Sgntin_row_00033_00003 = I76aab345d13c6678fe37a4a7133cfd7d;
assign Ia91800792941ec7cc60415c3f844e4ed             = conv_qin_00033_00003;
assign conv_Sgntin_row_00034_00000 = Ic76e72b434b47c10ebac3fac4ea50bde;
assign I71412803cc5229025487255aec62ec4f             = conv_qin_00034_00000;
assign conv_Sgntin_row_00034_00001 = I835b902949c2c4c09b757d4d35574a76;
assign Ibd89458312687610aa166a9538968851             = conv_qin_00034_00001;
assign conv_Sgntin_row_00034_00002 = I5f1609647f1e71cef4ba2d605c6c8445;
assign I1c3c4ce44610e04c5eef2fcbc2ea5114             = conv_qin_00034_00002;
assign conv_Sgntin_row_00034_00003 = Ib4f368fa3d3ec11d9ffb2ae9a2ae6310;
assign Id7c507d96098ee7a955af8a48ee5d72a             = conv_qin_00034_00003;
assign conv_Sgntin_row_00035_00000 = Ia1b617e3d141263b51e58c5ef0bd7a89;
assign If1607e907e626902ee26d15020a64c21             = conv_qin_00035_00000;
assign conv_Sgntin_row_00035_00001 = If343015b4815b01dae88bbb6f2017b3d;
assign I3ed5d0fca86f35b3d4b4a89c6147d0cd             = conv_qin_00035_00001;
assign conv_Sgntin_row_00035_00002 = Ic98f33c6a4613534bcc9b6bc4b4f2d17;
assign I599d01cfe6e54d8e45d64446c446818d             = conv_qin_00035_00002;
assign conv_Sgntin_row_00035_00003 = Idd0f3cfc5599481c954a2bfe69f044e5;
assign Ie15e4c1bcdb0e18085d4b320ac6a925c             = conv_qin_00035_00003;
assign conv_Sgntin_row_00036_00000 = Ie74c72742807ae4243748fd27d80d626;
assign I14834fc8e6489775359bcecf5a37ff4d             = conv_qin_00036_00000;
assign conv_Sgntin_row_00036_00001 = Ied8bd4b6fd0e4fbcced6d20eb7435f55;
assign Ic87c3d7762a18772972552162e1d1a8c             = conv_qin_00036_00001;
assign conv_Sgntin_row_00036_00002 = I6cbc06919b9c695d99621db6f8d768cb;
assign I157fdf8775206858c08682db3039b084             = conv_qin_00036_00002;
assign conv_Sgntin_row_00036_00003 = I641539560711ff1824bd90baa0f21f96;
assign I8f0a90e761111a613d2488285534a500             = conv_qin_00036_00003;
assign conv_Sgntin_row_00036_00004 = Ie624c4dad5036a25ca314b94cf3c4b95;
assign I5485d9edcafc6202f6e5f0969979802f             = conv_qin_00036_00004;
assign conv_Sgntin_row_00037_00000 = I8510240df7dc41f85ad58a39868a1fd7;
assign Icbaf92a8e9875bcb19a1d074779a9ea5             = conv_qin_00037_00000;
assign conv_Sgntin_row_00037_00001 = Ibe3d3e6bc58efc2e9d9eb1f96cdfe424;
assign I20c2057240417146df144b518b43d052             = conv_qin_00037_00001;
assign conv_Sgntin_row_00037_00002 = I72939e49bf2d9c6a84e404419fc644a1;
assign Ia30539545e66c4cfc16828140149180a             = conv_qin_00037_00002;
assign conv_Sgntin_row_00037_00003 = I95f0acd4f955058041c035789c3a4d99;
assign I71e101962e766a4d1484b3235359a4b5             = conv_qin_00037_00003;
assign conv_Sgntin_row_00037_00004 = Ibf4b3caa5655cfb6663f9b7e2383bbbf;
assign I7fe364f9f537cbef782e7007848a1c10             = conv_qin_00037_00004;
assign conv_Sgntin_row_00038_00000 = Ia0116a3cebf94318ed5b287960957ad6;
assign Ib0126fb335e32793c400a97c5a4a337c             = conv_qin_00038_00000;
assign conv_Sgntin_row_00038_00001 = Iaaaf373f7e6f55214915b93da9bd71d3;
assign I2993acb61f1abe529f8a60c94a438550             = conv_qin_00038_00001;
assign conv_Sgntin_row_00038_00002 = I0ceb14ac0187d804f9692e0c55b8e941;
assign Ic3b4752136ac08e343933ccc3a4ec47c             = conv_qin_00038_00002;
assign conv_Sgntin_row_00038_00003 = Iea424dd9d8916c4951b8746408b8a521;
assign Ic1efa395cc1fd2c5a1d1559fb169a5a0             = conv_qin_00038_00003;
assign conv_Sgntin_row_00038_00004 = I049d1c09c15def12ba7bae95fc1c3d55;
assign I52dcf5bace9cadcf8a895aaa6a8c1da8             = conv_qin_00038_00004;
assign conv_Sgntin_row_00039_00000 = Ic14760b65c6fe150c3c48e64389a41d8;
assign I6b1d01c3cb8fb51e43cdb788b89816be             = conv_qin_00039_00000;
assign conv_Sgntin_row_00039_00001 = Ibab1d13cd6a4f7b0c79c9f845339e53f;
assign I33b99994abbb5ecf8eed4de39033e4f8             = conv_qin_00039_00001;
assign conv_Sgntin_row_00039_00002 = I2919272e9ae3996a3e1d602ff72ba86d;
assign I39e6d3fb468aa40ea73535e81556ea65             = conv_qin_00039_00002;
assign conv_Sgntin_row_00039_00003 = I1db4ea6916125702e7fb09d0f742e60a;
assign I5b55c285f7e3e78447fee68532ab9f7f             = conv_qin_00039_00003;
assign conv_Sgntin_row_00039_00004 = Ide06ba186ddb179b489ba6e3e209e3e8;
assign I13a9eec6175e695ab8bc4516cf57d6ec             = conv_qin_00039_00004;
assign conv_Sgntin_row_00040_00000 = I6f420c64640dfb0c001f57df7e3b4504;
assign Id0344146d1a53d418add6d2b185377dd             = conv_qin_00040_00000;
assign conv_Sgntin_row_00040_00001 = Id75c23e80cdf25d883806ed20d4ae783;
assign I20590d8fb97ec0b2164ffe17826136a7             = conv_qin_00040_00001;
assign conv_Sgntin_row_00040_00002 = I4d4901ff372f6820ca9c8c29cefa664a;
assign I05370777439b01811fe7f750d2f724f4             = conv_qin_00040_00002;
assign conv_Sgntin_row_00040_00003 = Ice0234f25de4ab1f03a3cb01a2d61dbf;
assign I8cab9fba615b94fd4bb6934325be8ab8             = conv_qin_00040_00003;
assign conv_Sgntin_row_00040_00004 = I1b78785ebe2e7f77a3125a6334c4dc54;
assign Iee73a7c685a4cee03f33d3ef379b1c8a             = conv_qin_00040_00004;
assign conv_Sgntin_row_00041_00000 = I9eb87e62d23bc87d7cd82c0f329f247f;
assign I32fcb28a27356bc6f403528836ea4c1f             = conv_qin_00041_00000;
assign conv_Sgntin_row_00041_00001 = Ied6c684cdd280b41ffab93a026d27282;
assign Ib74a56900c1f8b159ad381f61acee801             = conv_qin_00041_00001;
assign conv_Sgntin_row_00041_00002 = I1ca188bcdebbf41d84f7a5220bd1d195;
assign Ieb38fa62119a5a77c060d6634e051298             = conv_qin_00041_00002;
assign conv_Sgntin_row_00041_00003 = I9322a2a61900943075bbc23c72a3f65d;
assign I86e495dc894d2aace15c1aff89798bf7             = conv_qin_00041_00003;
assign conv_Sgntin_row_00041_00004 = Ie79c93f1703121713fb9401617f349a8;
assign I740dc91716e3906ad078e2c7cc3c925a             = conv_qin_00041_00004;
assign conv_Sgntin_row_00042_00000 = If9a5d830e3ade0fd96b98f5949f165f0;
assign I081b38dbb37d4c14a6a9fd3fefa13daa             = conv_qin_00042_00000;
assign conv_Sgntin_row_00042_00001 = Ie7a68c2b368a295f95571bc4a109b9f1;
assign I633a74e4dfa841c9fd13dbb6564c8493             = conv_qin_00042_00001;
assign conv_Sgntin_row_00042_00002 = I0152dc6e6a7acd72a2144623e63998ef;
assign I0b7b4c0a8503c751229edfe0237cc903             = conv_qin_00042_00002;
assign conv_Sgntin_row_00042_00003 = I9b560d9baf8a7422b0dd84720e924ced;
assign I43b380be6df7df0d354223d0a0d6d6b6             = conv_qin_00042_00003;
assign conv_Sgntin_row_00042_00004 = Icf25f076eec2bf81c899c66f6cfbebc0;
assign I514d2dc697e9b39ba027c418a6df6cb9             = conv_qin_00042_00004;
assign conv_Sgntin_row_00043_00000 = I7332e088bbff69db19c62685e033d26a;
assign I3ea4c33a9419820ed54460eb64134dff             = conv_qin_00043_00000;
assign conv_Sgntin_row_00043_00001 = I1b6abc8fbab3849b285e9f88a4fe867b;
assign I80f3c8559da8e97bc5397bb8b621a0bd             = conv_qin_00043_00001;
assign conv_Sgntin_row_00043_00002 = Ic14f948884da19a272a4760ffaab9ea9;
assign Iaf4ae293c576af16f5f43a8b86c1aa3d             = conv_qin_00043_00002;
assign conv_Sgntin_row_00043_00003 = Ice5f7168aeb940d48093cc9df7cba36b;
assign Ib42816335dd8475dcc78662c4c0786c1             = conv_qin_00043_00003;
assign conv_Sgntin_row_00043_00004 = Ic5c837a0556d1cb66edbf0294d08283a;
assign I782726e317a2aada9e755bcbc4b0d3fa             = conv_qin_00043_00004;
assign conv_Sgntin_row_00044_00000 = I3600031716c2b4e21c9f577d34e033dc;
assign I1eede74f12d37331b399eb7136bc621f             = conv_qin_00044_00000;
assign conv_Sgntin_row_00044_00001 = I859d795a7d141eb777c1f3c038203794;
assign I343c9efe71164c01e9c7d599e032864a             = conv_qin_00044_00001;
assign conv_Sgntin_row_00044_00002 = Ib9c194ec16f435a9357cb344cf25bdcc;
assign Idb72c046c5996fbbd80b706666ffbd92             = conv_qin_00044_00002;
assign conv_Sgntin_row_00044_00003 = I69d82ab774d52c219509e993e7cc4deb;
assign I141fb1cbe09f9abe282cffd4de815d25             = conv_qin_00044_00003;
assign conv_Sgntin_row_00044_00004 = I51ff4bda38746682e3cd4c68118c3216;
assign I11eb26cf0f0b3a334e8f7317bf8d9eb0             = conv_qin_00044_00004;
assign conv_Sgntin_row_00045_00000 = I2eac5b39c6f485c9ae0bd341f894633d;
assign Iad354d876cb9fc72fc0143e6f7da9357             = conv_qin_00045_00000;
assign conv_Sgntin_row_00045_00001 = I12a18a1f8d4416e9bc8abee6ac3dacfc;
assign I92d9fec22d36b1baac8bd78abfc1bbd5             = conv_qin_00045_00001;
assign conv_Sgntin_row_00045_00002 = I45bdd0cfe107da0d57cad1333bf95e3b;
assign I262f2390e77ec486ccd3a6ed05816e2d             = conv_qin_00045_00002;
assign conv_Sgntin_row_00045_00003 = I768720af835b02a8dab376ef23d17a15;
assign I461195b7ae78743e09ee50486ad6ebe5             = conv_qin_00045_00003;
assign conv_Sgntin_row_00045_00004 = I1c074a53e6c0f2467bcdd7c952f51670;
assign I26cb63ba20245b2c332b09e25c4409aa             = conv_qin_00045_00004;
assign conv_Sgntin_row_00046_00000 = Id3de87169c440f95d406693ef77cacd6;
assign Ibac5e7b6d4bf5cd6926358318f0c418f             = conv_qin_00046_00000;
assign conv_Sgntin_row_00046_00001 = Iedc463e359dd3003d9f7e50f3e858e93;
assign I0d53bb5344cabe5fa5ce3ecf7122a260             = conv_qin_00046_00001;
assign conv_Sgntin_row_00046_00002 = I23955b54e486f0f0d21a2809a9472b86;
assign I94f1724740defe5bb7e40041d0e266a0             = conv_qin_00046_00002;
assign conv_Sgntin_row_00046_00003 = I24075f37c6bbd90c83370de1a2e58af2;
assign I6ae2523095237282533e0b5f1c26b488             = conv_qin_00046_00003;
assign conv_Sgntin_row_00046_00004 = I37c49c5a2af240496f5a5706b0d42ea6;
assign Idd7691d31f8d0c09ee988116d574ec59             = conv_qin_00046_00004;
assign conv_Sgntin_row_00047_00000 = I44daa5992b00e7af19adbee70bf01f2b;
assign Ia0d940e16c8cbd4f7544f5a5cd7d83b2             = conv_qin_00047_00000;
assign conv_Sgntin_row_00047_00001 = I457ae11ad90c8478751eb4b42764e158;
assign I23eb1dc4d1c992f804dd04a2d823c778             = conv_qin_00047_00001;
assign conv_Sgntin_row_00047_00002 = Ida3dd5e990ce3c237e9628a9a090901e;
assign Ia630e59cbce82a570ae3890a6c0221e5             = conv_qin_00047_00002;
assign conv_Sgntin_row_00047_00003 = Ifbadefd3a7ab50719a703400ddd742c6;
assign Id1bacd13718f7c29c26b63c239d04dd8             = conv_qin_00047_00003;
assign conv_Sgntin_row_00047_00004 = Ia94c439131e1df5c95fc8ad3cfdba473;
assign Iecc02842a2d2b9b9e8187f2d39e62e05             = conv_qin_00047_00004;
assign conv_Sgntin_row_00048_00000 = Id88a7edf897eea1b4a137141789a04f5;
assign I157bd468200e63385583b9045758d81e             = conv_qin_00048_00000;
assign conv_Sgntin_row_00048_00001 = I70dd1350d65155ee7b562f4c79024a3d;
assign I09e9a3cd4c12d204f760758e873a177b             = conv_qin_00048_00001;
assign conv_Sgntin_row_00048_00002 = Idc445d3f5b3b62562b0ac83e5f17e92a;
assign I32701d9e4b96853c53f0ab651a6a4ba2             = conv_qin_00048_00002;
assign conv_Sgntin_row_00048_00003 = I723a6fee3b2496f23c48b3584f8bf9ce;
assign I5551342f1751fc64f32744a46b9649be             = conv_qin_00048_00003;
assign conv_Sgntin_row_00049_00000 = Ied638fee34f8baed4154b0b72e43a21e;
assign I7a0eada108891aba06cecab5071232c9             = conv_qin_00049_00000;
assign conv_Sgntin_row_00049_00001 = Ief03713f5cf37200373a20d42c7fc9eb;
assign I4df3d4dac24877b14e6d361bafc1a800             = conv_qin_00049_00001;
assign conv_Sgntin_row_00049_00002 = I3ac0799861144b599995318bdade2114;
assign I765a8825e42180a6c63f7b33703bb483             = conv_qin_00049_00002;
assign conv_Sgntin_row_00049_00003 = I648b62fa0bc2185c1756ee531e8e34de;
assign Iff7c29299f005c1cd5a16b64601e727e             = conv_qin_00049_00003;
assign conv_Sgntin_row_00050_00000 = I1b43f29e0ddb72467befd6f3a9c1c829;
assign I3c128efc9f80c9b8334bf7b61de71b43             = conv_qin_00050_00000;
assign conv_Sgntin_row_00050_00001 = Ic07c650e6e49892a41cfaf3a37471426;
assign Ied00d87af99ae55144fdde41ebfc1357             = conv_qin_00050_00001;
assign conv_Sgntin_row_00050_00002 = I4082b3564c1949a19ed35bd5a88e1ef4;
assign If2539da6722562bbf31786fd0036666a             = conv_qin_00050_00002;
assign conv_Sgntin_row_00050_00003 = Ife631f9a3c4c64a3d92aa9586ae75f3c;
assign I17a5446e942bcc1dc2c96930e0a87a70             = conv_qin_00050_00003;
assign conv_Sgntin_row_00051_00000 = Id0f4dbb72da33748d8baf723c5a32567;
assign Ia5eba52d169755c507b9e0094e467fab             = conv_qin_00051_00000;
assign conv_Sgntin_row_00051_00001 = I44ccc3ae897109dd51f9afeef93daca4;
assign Ib9ceb8315f0cd848f861bab677c2c694             = conv_qin_00051_00001;
assign conv_Sgntin_row_00051_00002 = I73bbf90b625d56f663ad10f9d21d8e76;
assign I8e96c69e7d872be23229353808c34953             = conv_qin_00051_00002;
assign conv_Sgntin_row_00051_00003 = Iaac1d82f0846fce1bd88ebf8e60300ac;
assign I719b67f84e07e90dfd29a8cd5d94cf39             = conv_qin_00051_00003;
assign conv_Sgntin_row_00052_00000 = I002820a37fa7c6c504c487df4368e2cf;
assign I3e4754acc31d99bc71525789bdee0c1a             = conv_qin_00052_00000;
assign conv_Sgntin_row_00052_00001 = Ib0bb71b1f8829347b3a9a7543f9dd964;
assign I0899e8fec1a7209cd94757c0b2f87c9a             = conv_qin_00052_00001;
assign conv_Sgntin_row_00052_00002 = I1dd4671765f8826c2fe20c592c5e32c8;
assign Ied029d0bdea3bf134744c99426fa72dc             = conv_qin_00052_00002;
assign conv_Sgntin_row_00052_00003 = I3175159add7b814df637c2db8feb43f6;
assign I5aba6218461e8d571be03a3ef041ebaa             = conv_qin_00052_00003;
assign conv_Sgntin_row_00052_00004 = I48cd09f035f668536cd288a23010b07b;
assign I2c835dfb3596b8bf057a7cc21122c81f             = conv_qin_00052_00004;
assign conv_Sgntin_row_00053_00000 = I76992221b1edff5684c482df7ac4693d;
assign If6e745bb85abba7282dae1f6f701225e             = conv_qin_00053_00000;
assign conv_Sgntin_row_00053_00001 = Ib13436ad16a37d656d6b1ee95b9aee20;
assign I918c46173eebc5b2a95e041cfd91d958             = conv_qin_00053_00001;
assign conv_Sgntin_row_00053_00002 = I47b0847946b0e00961233ac0101fa2a7;
assign Ic8be2c94235fb40f78da33179ce4873a             = conv_qin_00053_00002;
assign conv_Sgntin_row_00053_00003 = If2042aede3390bd208a281f0380c95a4;
assign Ia3104c69fb4f7abfb5efa3874169a7ad             = conv_qin_00053_00003;
assign conv_Sgntin_row_00053_00004 = I119b2e5c2fea5338244c4019884af26f;
assign Ib71b3d357c98dcdfae5c777ca3082275             = conv_qin_00053_00004;
assign conv_Sgntin_row_00054_00000 = I3751f191f5009322acb7c9be4f8d7129;
assign Iadfc60386481092ae85cc148a2c40abb             = conv_qin_00054_00000;
assign conv_Sgntin_row_00054_00001 = I14fa7aebb608d4a3d67176ba27d34d9a;
assign Ie21a2c9b22e7bf8425fb5c0f33e5f4f7             = conv_qin_00054_00001;
assign conv_Sgntin_row_00054_00002 = I7b813d83b13bb7bc13940cf5714c06ba;
assign I7c3291f0250d13ca94802b0b071a95c6             = conv_qin_00054_00002;
assign conv_Sgntin_row_00054_00003 = I0eaa22f5eca8f33dd254fe241017a098;
assign If79d1d378f7c6fd29fc3335ec5f5c51d             = conv_qin_00054_00003;
assign conv_Sgntin_row_00054_00004 = I2bd34b2fd12f12bc301fd0d5d69c0fb6;
assign I086bf19f620c8a8f6888e775cb1ed7f4             = conv_qin_00054_00004;
assign conv_Sgntin_row_00055_00000 = Ie517386cb5832e406fefc5e85eb2e7d1;
assign I4a8abfa0896ce414d9b98093ef84455f             = conv_qin_00055_00000;
assign conv_Sgntin_row_00055_00001 = I3fd0fa3b774d30a267d61e9427d09f3f;
assign Ic7147944f8835e26b9838fdbdc18ca41             = conv_qin_00055_00001;
assign conv_Sgntin_row_00055_00002 = I4ee312036de8c08300c358edcff1e1e9;
assign I7e393e6c1d1bc44daaab120d55f5dd59             = conv_qin_00055_00002;
assign conv_Sgntin_row_00055_00003 = I1d98943b01a6a2d8c4db18b98dd62f5c;
assign I356d747600182675699a2d2634d4c5ce             = conv_qin_00055_00003;
assign conv_Sgntin_row_00055_00004 = Ib715b1e0061b84ce614a30d961a83e7e;
assign I802c554d5b04af6b949677819a4966ed             = conv_qin_00055_00004;
assign conv_Sgntin_row_00056_00000 = Idc07dc30c0a957e474546ac7a60df38f;
assign I4f8792c18bd07b23e82bbc44b4ca947f             = conv_qin_00056_00000;
assign conv_Sgntin_row_00056_00001 = Ifc640243288c9b37b7eb9e00351b23f0;
assign I3459d98131faef5a5040a03847890b55             = conv_qin_00056_00001;
assign conv_Sgntin_row_00056_00002 = Ie83fa8157a7cce44c2e25f46ce897dbb;
assign I512cc8f6519aa08aee18225b56d47c9f             = conv_qin_00056_00002;
assign conv_Sgntin_row_00056_00003 = I570c036d0237c53bb069c52d621e539e;
assign I4a41999cea9357a85c73a0af509eeac9             = conv_qin_00056_00003;
assign conv_Sgntin_row_00056_00004 = Ief8c2838abac83370fd7ec25c06d509b;
assign Iceefb06cb3715e1b41e6f7d89420e5ba             = conv_qin_00056_00004;
assign conv_Sgntin_row_00057_00000 = Iad90879acba3fc2101829549264960f3;
assign Iaa5b2807e5cc2403c5787eeb3d10ca6b             = conv_qin_00057_00000;
assign conv_Sgntin_row_00057_00001 = I951dedd7af44c3865a8f36888432d0c9;
assign Iace01234164c8a9f7c98eeb83268745b             = conv_qin_00057_00001;
assign conv_Sgntin_row_00057_00002 = Ia7606050c683ecefc510ba92ac539a9c;
assign I22c8ccd4a9018ad1c129aa058bf579d8             = conv_qin_00057_00002;
assign conv_Sgntin_row_00057_00003 = Id3b089fb6edd5bcfdbca142fddd5ff89;
assign I87d6a5d30c3e4202cf51f33c7a770c51             = conv_qin_00057_00003;
assign conv_Sgntin_row_00057_00004 = I561d79eb079915c0b1732cbddb119c2d;
assign I56948bc48c0220893d68004615a6ebaa             = conv_qin_00057_00004;
assign conv_Sgntin_row_00058_00000 = I2eb08ebaa07a1004638cdd61a7209b7d;
assign I698b1dbc9d8664d1c86c7a763d97b3b7             = conv_qin_00058_00000;
assign conv_Sgntin_row_00058_00001 = I46e1047bca2b38e62b4de80d1d2249de;
assign I68b575fcbc5321d4d26a22bcdbb506f6             = conv_qin_00058_00001;
assign conv_Sgntin_row_00058_00002 = I41796b587316c600bf583edc62649bd8;
assign Ib6aded6c73a8cc3cb964b0ae895b859e             = conv_qin_00058_00002;
assign conv_Sgntin_row_00058_00003 = I0a569f6536789efb7ad2377c11842830;
assign I6ca8a1fa2c72b1c61d11dc7d1ba5f37b             = conv_qin_00058_00003;
assign conv_Sgntin_row_00058_00004 = I8bb75bf828d5ef337fa6a965808e4638;
assign Iec1368f034655d61354ab5b5e94d7d89             = conv_qin_00058_00004;
assign conv_Sgntin_row_00059_00000 = I47cbb92d2284aef7b9e56e88f0ba6f7e;
assign I08ece7cd684e593e02321612b7a88cee             = conv_qin_00059_00000;
assign conv_Sgntin_row_00059_00001 = Ib99e1b93fb7fbda260d93eea3d24c3e9;
assign Icdcd83341f6b5c404f91ec7e97d0550c             = conv_qin_00059_00001;
assign conv_Sgntin_row_00059_00002 = Iee6e52d75c093a24eb4e5e0b45feb256;
assign I82f266e5792cdb6e7ebd264e246161f5             = conv_qin_00059_00002;
assign conv_Sgntin_row_00059_00003 = I19b73c5c93a71e90f620572f23f0e6d2;
assign Ie1b7257c99831ec5864f65958ecf14fb             = conv_qin_00059_00003;
assign conv_Sgntin_row_00059_00004 = I11ba339c8250d07b497c88a39a6df1ac;
assign I1e43c0aeeb8a2461d208eba24967af30             = conv_qin_00059_00004;
assign conv_Sgntin_row_00060_00000 = I8a4c1f23212ff846400651b100add502;
assign I11c1fc94a3bd6dffa17e1571cc6ae97c             = conv_qin_00060_00000;
assign conv_Sgntin_row_00060_00001 = Ief18a19d451f05f6051e3cc8de16d73c;
assign Ica6707efd6d44ba6bbb87c0593a3d828             = conv_qin_00060_00001;
assign conv_Sgntin_row_00060_00002 = I7009c18515dd43d8dd2e5d1ee6779641;
assign I939368b76d98b43826c68c7f468a5632             = conv_qin_00060_00002;
assign conv_Sgntin_row_00060_00003 = I173aa69cf52114e223ac1410d90b4bfe;
assign Ia6eb85b127cf9c1a437611556296b967             = conv_qin_00060_00003;
assign conv_Sgntin_row_00061_00000 = Iada5bc4a51dc1bf57bb9cca11326bdff;
assign I93bb43c1b89d4c70a57bdc019d64fd22             = conv_qin_00061_00000;
assign conv_Sgntin_row_00061_00001 = Ib6fbe376477afa58bfcc17a8564f78b2;
assign Iae449b74e50e0907feae9e60f2329426             = conv_qin_00061_00001;
assign conv_Sgntin_row_00061_00002 = Id48fe0672aa98f987162931527e9f9bc;
assign Ibfacfe5b83819afe7fbd4bffa2d6d4e2             = conv_qin_00061_00002;
assign conv_Sgntin_row_00061_00003 = Ia4e89e99acb95f4183474b94798ca35d;
assign Ieba89aa901e61218074af53a2484a74b             = conv_qin_00061_00003;
assign conv_Sgntin_row_00062_00000 = Ic1927bb3335f6a28c0816eba12d3975e;
assign Ie0ee5445c56a5f9b41640b57422206de             = conv_qin_00062_00000;
assign conv_Sgntin_row_00062_00001 = I5b8a1e1a6b904b0f6822c224ee0486e3;
assign Iacbb4daf5ce5c7eb1a2afe30d0cb5382             = conv_qin_00062_00001;
assign conv_Sgntin_row_00062_00002 = I8be4711146486fea913843e497065b50;
assign If08370fd0e8af818c6db20f43e74034d             = conv_qin_00062_00002;
assign conv_Sgntin_row_00062_00003 = If4c36727ab1c29bf78f72e8acfc00d7c;
assign I8b3b875c6c07bd97ba598a5139156fa4             = conv_qin_00062_00003;
assign conv_Sgntin_row_00063_00000 = I9b096ce09467c10f448496fda13987d2;
assign I680be647bf2a62e0ee9b5d379dc87b4f             = conv_qin_00063_00000;
assign conv_Sgntin_row_00063_00001 = I57b7b48f13436b19a8d6a47e014eb41f;
assign Icbfbb37bad6344005dd233b3605a784f             = conv_qin_00063_00001;
assign conv_Sgntin_row_00063_00002 = I5446c1c323774715371c73bd1be66697;
assign I83330fef69470d2f5def8e6d7d9c50d2             = conv_qin_00063_00002;
assign conv_Sgntin_row_00063_00003 = I6426943b4ab66f17c2b7b399ccc7a6a9;
assign I7b33ddad346077928620344542b9481e             = conv_qin_00063_00003;
assign conv_Sgntin_row_00064_00000 = I595665d8128bb87ab62741d7ac520a4b;
assign I8d0a1ae4c47edf1f2b99d1175aaa7197             = conv_qin_00064_00000;
assign conv_Sgntin_row_00064_00001 = Ic920452d5997a8477724fa78c86c0fba;
assign Ie5757e7b1647ab7d43cdbcf98cbb77fc             = conv_qin_00064_00001;
assign conv_Sgntin_row_00064_00002 = I3a8e9e7d2cd6751e8500a5567cef5acc;
assign I0539d598bbe3d50940329a282c801328             = conv_qin_00064_00002;
assign conv_Sgntin_row_00064_00003 = Ib0dadebad37d9ea9d01350054872863c;
assign I8acc93b34974c1e708b0e1591f7b2d3d             = conv_qin_00064_00003;
assign conv_Sgntin_row_00064_00004 = Iddcffa815489773b3688fd68dba18bd8;
assign I11d967a5c5d14c88b5587d4cfed1d05f             = conv_qin_00064_00004;
assign conv_Sgntin_row_00065_00000 = Ife0952b85f14a960007b67646b0cd969;
assign I6da2b3a481ee71b85f3087b36b399288             = conv_qin_00065_00000;
assign conv_Sgntin_row_00065_00001 = I4d54dd2ee2f32909098d3cc2b6689220;
assign I280e20c20c0b4f26278b3de9b2ff84e4             = conv_qin_00065_00001;
assign conv_Sgntin_row_00065_00002 = I797c9cb725f88c07be28f017871d17f8;
assign I544f6263f16cd5e0b7cf28c511a8f6e3             = conv_qin_00065_00002;
assign conv_Sgntin_row_00065_00003 = Ie165d0729542c81ca89f45d15e0afd3d;
assign Ie11da10808c4ca84f399535df6261307             = conv_qin_00065_00003;
assign conv_Sgntin_row_00065_00004 = Id00642563679fa9a6696f8e7bbdf6576;
assign I27458d76b3ac6520fb379405c6b2956f             = conv_qin_00065_00004;
assign conv_Sgntin_row_00066_00000 = I258c45897919cec5c6acaddee7f3a41b;
assign I508bbade361787127e1a2e8687ec884c             = conv_qin_00066_00000;
assign conv_Sgntin_row_00066_00001 = I1e11f0088959aa40b4ad1a047b59caf4;
assign Ic19486b6ab0373b9c0ad8f7597782d8f             = conv_qin_00066_00001;
assign conv_Sgntin_row_00066_00002 = Idce46f6d03376bea1ba361e8c59f8bd1;
assign Ib8e68a77ad8b9e7cf415bee17645c3f9             = conv_qin_00066_00002;
assign conv_Sgntin_row_00066_00003 = If17c0096ce34b88007247bf4c429d5c4;
assign Ie84be0ae8311d906eff08f7f5b214943             = conv_qin_00066_00003;
assign conv_Sgntin_row_00066_00004 = Ifda1c55899cd3506853cc82b450b3936;
assign I2525111a2fb5f10d64bbd16e148653b8             = conv_qin_00066_00004;
assign conv_Sgntin_row_00067_00000 = Ic69094123b75ae36e3e54f179a9f2cb5;
assign I691c84d81c60a462e28e2b2bae3ea845             = conv_qin_00067_00000;
assign conv_Sgntin_row_00067_00001 = Id182a776b03f48fb139c28194ae7ab6b;
assign I4904ab14b19fa1b6befc218bc7be3842             = conv_qin_00067_00001;
assign conv_Sgntin_row_00067_00002 = I65171c9ee8449407484e5c82d13c6751;
assign I0ff382edfc8051459657ffa3899f5f73             = conv_qin_00067_00002;
assign conv_Sgntin_row_00067_00003 = I92eb6f60c14ee9eecb01718b01ea980f;
assign I8f94dbafaac589ac9f14b56d4556ff96             = conv_qin_00067_00003;
assign conv_Sgntin_row_00067_00004 = Ib5d1a7cdbcba0b654c12063d4f1768e1;
assign I7b7cbcd1c6d2a2eeaaff474536a69eed             = conv_qin_00067_00004;
assign conv_Sgntin_row_00068_00000 = I07abbbd75d91018ac53f53e64cffafb9;
assign I58dc9cce6384160c0a85c6efb3319cdb             = conv_qin_00068_00000;
assign conv_Sgntin_row_00068_00001 = I4cdc955fa9afc75c2c977de4ec540e1e;
assign Icde3e6dbcf985682041f30903ad95572             = conv_qin_00068_00001;
assign conv_Sgntin_row_00068_00002 = Ie79ce8adeef2c3c24a3386f054d0cf5b;
assign I644ee0055a55f54ab3544bb532e39c61             = conv_qin_00068_00002;
assign conv_Sgntin_row_00068_00003 = Ifc2963762403a00c4f3662b2863c991e;
assign Ic90b98708faa8c8b75d4bd9a52c292f7             = conv_qin_00068_00003;
assign conv_Sgntin_row_00068_00004 = I5e8ed024e2f2548bb375a2ecf1918a5f;
assign Id2a7f0781d18dccc7c4e0b383b7cddfa             = conv_qin_00068_00004;
assign conv_Sgntin_row_00069_00000 = I256050251d23250854ff337bef28e460;
assign I734e601f5f9d568a44a48834559e04db             = conv_qin_00069_00000;
assign conv_Sgntin_row_00069_00001 = I20ffba20af04b99954bf719589e90d1a;
assign I749e987266a20840bb8a4b1a2a2fc5b0             = conv_qin_00069_00001;
assign conv_Sgntin_row_00069_00002 = I7353ebf3a1cde89d2bb3fa667f7f5485;
assign I9d2864024148337277523ef7fa2e1600             = conv_qin_00069_00002;
assign conv_Sgntin_row_00069_00003 = I97e82e5f6775d1e31537b891597223bd;
assign I754563caea429d3d0e22df5d193b84eb             = conv_qin_00069_00003;
assign conv_Sgntin_row_00069_00004 = Id25deba967318f049de8163e67262f4b;
assign If8bc141d98ebe1be7fa81cde5c65868e             = conv_qin_00069_00004;
assign conv_Sgntin_row_00070_00000 = If876ca6a14ffb4323503ed46666bc25f;
assign I11094e852295755925c3c61f1df81643             = conv_qin_00070_00000;
assign conv_Sgntin_row_00070_00001 = I5109afc4dc91780e05704ea5e1399e3e;
assign Ic419255414995e7168afb97b051fa64f             = conv_qin_00070_00001;
assign conv_Sgntin_row_00070_00002 = I621b20d29d3a9a9f41065bc3c3bbd2d8;
assign I202f88fdc946494d55fc8831c2e8a34c             = conv_qin_00070_00002;
assign conv_Sgntin_row_00070_00003 = I76fd9005abd511c3c5bf6c77de8bf2f3;
assign Ib60d4ac0fcadcdfce5a14fb92f58423f             = conv_qin_00070_00003;
assign conv_Sgntin_row_00070_00004 = I925f6b549a25cdc8f85152eb21ea3b58;
assign I8645e1326c66f5efef4b9c923599d1a3             = conv_qin_00070_00004;
assign conv_Sgntin_row_00071_00000 = Ib42d37576e3aff3d205f1f8822cc58b5;
assign I2afeb2a7b199c0c6738938f156ae4274             = conv_qin_00071_00000;
assign conv_Sgntin_row_00071_00001 = I3ce10718a2211184999663c3c2493cc1;
assign I7992ea31927b4f0e268462a3b0f18c5d             = conv_qin_00071_00001;
assign conv_Sgntin_row_00071_00002 = I06b48093d4c9b0327c3efc6fa4ca7daf;
assign I484545c4d2c869d79eb17f51e11070a3             = conv_qin_00071_00002;
assign conv_Sgntin_row_00071_00003 = Ie8e29053f122a9247b0dec291c6ef4f3;
assign I280fa9d114e227cd649bf0e55e845651             = conv_qin_00071_00003;
assign conv_Sgntin_row_00071_00004 = I9b49e1acb81ef5b088b808d2e4ce9954;
assign I0426ef66185128dd1ef4dbb68dcda585             = conv_qin_00071_00004;
assign conv_Sgntin_row_00072_00000 = I364ed3f83c49626bc3b939e53524d9c7;
assign I7a2e554d07bbea291f2cfc18694fca3a             = conv_qin_00072_00000;
assign conv_Sgntin_row_00072_00001 = I8188dd7cb03854c6f709de06ff785d91;
assign Iace8b3b3a4c16763132b5aaa6b24212d             = conv_qin_00072_00001;
assign conv_Sgntin_row_00072_00002 = Ie7cfdd25541414ff3f8d6e5d7677fbe5;
assign Ib2f5f5fc77ea8b529f2471c54388f2d1             = conv_qin_00072_00002;
assign conv_Sgntin_row_00072_00003 = I6386a4dd26e7c36165dc265b3a2c93cf;
assign Iddd954df5bae9b4240e0512f746669a9             = conv_qin_00072_00003;
assign conv_Sgntin_row_00073_00000 = Ia659126b51468cfef48c97a135a71500;
assign Ie5f8620371236cb11c9e88c16b509ee8             = conv_qin_00073_00000;
assign conv_Sgntin_row_00073_00001 = I866b30a63b3b5fb708934a1cbb0e1d9a;
assign Idf600b93ee1018ecf969ed7944b6bc7b             = conv_qin_00073_00001;
assign conv_Sgntin_row_00073_00002 = I2b7822d5d77aaed61eee87570564df76;
assign I7f90f96c0260560ad5e6dc7448b2670a             = conv_qin_00073_00002;
assign conv_Sgntin_row_00073_00003 = Ia20709f08cfff3a51d4af1e81d640400;
assign I29e940970d87e8e09b26ab1b0b8f2286             = conv_qin_00073_00003;
assign conv_Sgntin_row_00074_00000 = If1c0a3726041f70e508d68cbf6e40e04;
assign If4d75f83299a21802b6fbe136913489f             = conv_qin_00074_00000;
assign conv_Sgntin_row_00074_00001 = I019e399a1cef87745e025a7d74e94db0;
assign Ibba4e82d1510ddc16eb4ef64893cec02             = conv_qin_00074_00001;
assign conv_Sgntin_row_00074_00002 = I0dccb8eaad52ce4d780696a8485420f1;
assign I108c269ceec4adcff9afeda01101b838             = conv_qin_00074_00002;
assign conv_Sgntin_row_00074_00003 = I1ff042bdb52aac5d69791e96e2f9706c;
assign I488f6d9676aa85a55d030bf12e8997a7             = conv_qin_00074_00003;
assign conv_Sgntin_row_00075_00000 = Ice1ce5b4c30841dd92268559ebadafcf;
assign I5395ee57418c31e11cf847f0f514ec19             = conv_qin_00075_00000;
assign conv_Sgntin_row_00075_00001 = I3d149293f106ae8680c7f4702daa0bd6;
assign Ie9b9221b2122087cd5f309570b6d31ca             = conv_qin_00075_00001;
assign conv_Sgntin_row_00075_00002 = Id17ada8dae3f9810d1892d34f2288859;
assign I4eadce87f47df6d8f0e4acd057de5a09             = conv_qin_00075_00002;
assign conv_Sgntin_row_00075_00003 = Iaa2cbf59f6f61198b4fcf5a741cd5bc8;
assign I99d761b75ade1fb2e8afbb1a77752609             = conv_qin_00075_00003;
assign conv_Sgntin_row_00076_00000 = I3eeeb1949945032d6c1759875426b733;
assign Iff125392fa39afebae1637a19c4e23ec             = conv_qin_00076_00000;
assign conv_Sgntin_row_00076_00001 = If2dfcbf493b761fb5d7c622e739b23f3;
assign I9c633aa620cca127b0ff8cf882178e76             = conv_qin_00076_00001;
assign conv_Sgntin_row_00076_00002 = I3f5053e519a928640ae49cf4e5b39d1e;
assign I4e08021c0235fafb60200aab97827a8f             = conv_qin_00076_00002;
assign conv_Sgntin_row_00076_00003 = I01c94743a11042e75638ba6618356203;
assign Iac4e3d20178049f9c59abf374752dccc             = conv_qin_00076_00003;
assign conv_Sgntin_row_00077_00000 = Ic2b000c3b2ca3beff2d427caab04701a;
assign I3e59b2419c7dd1553b792d536208514e             = conv_qin_00077_00000;
assign conv_Sgntin_row_00077_00001 = I1c2ee281cd47a8414851c5e1c758ea65;
assign I86255756ddd1f88b74e070b19f8c3bfa             = conv_qin_00077_00001;
assign conv_Sgntin_row_00077_00002 = Ia3ef2f70c5abaa852586a33c505aee0d;
assign I91a6408a11fab36a8ba3dbd3f895a803             = conv_qin_00077_00002;
assign conv_Sgntin_row_00077_00003 = I0a0340a0e52145f3597accfe4a4e8624;
assign I618d33f26badabfa578908903a613bce             = conv_qin_00077_00003;
assign conv_Sgntin_row_00078_00000 = I3c3c22bf63e55a81ae91b1dd1ef615a0;
assign I8d7c1fe2e33bbd45379b0325a3c5e989             = conv_qin_00078_00000;
assign conv_Sgntin_row_00078_00001 = Ib02268d5048c7c8e83118070e927453f;
assign I56bf74b5890ec67090f499afdc0a9c88             = conv_qin_00078_00001;
assign conv_Sgntin_row_00078_00002 = I30be0b18e4415ca50f2d8149efaaafe6;
assign I739267bcc50c54b8a685cb3c6afc5cc1             = conv_qin_00078_00002;
assign conv_Sgntin_row_00078_00003 = I3bb4d24caaa0882a75125e466070f0b1;
assign I822d7973afe090b2764335f1b72dfd0e             = conv_qin_00078_00003;
assign conv_Sgntin_row_00079_00000 = Iaf36ce8598a29573979c683a5e2cf9fd;
assign Ibddfda6413e3dd2f483c3174ea836b6a             = conv_qin_00079_00000;
assign conv_Sgntin_row_00079_00001 = I82f0e5a32d1bcd761a74f1f9ce8c88ba;
assign Ie421da1dc5aaea57c50d0c7d9c5a2717             = conv_qin_00079_00001;
assign conv_Sgntin_row_00079_00002 = I659322a9fd0d5eac514437b02e0491b3;
assign Iebf769a6bdaf214c1006c55c608d4eda             = conv_qin_00079_00002;
assign conv_Sgntin_row_00079_00003 = I44ead0ab5ccc53226fccc03024643771;
assign I12c1035353e553b3b6a13bb174ce6020             = conv_qin_00079_00003;
assign conv_Sgntin_row_00080_00000 = Idc2a9c6dd8d2aa912548c918c8a488f4;
assign Ibaf2f1f8bda2f6b932dc30f8369c0e1f             = conv_qin_00080_00000;
assign conv_Sgntin_row_00080_00001 = I08f22261d5713c0636d77c7938f592d6;
assign I88a61cf72347d695489909d0819332ab             = conv_qin_00080_00001;
assign conv_Sgntin_row_00080_00002 = I04c734eb876aa722e84d6b9edd297978;
assign I39289e6385a9bc378a9b8dd440249a7f             = conv_qin_00080_00002;
assign conv_Sgntin_row_00080_00003 = Iaded125f7fd5c833e7206dd7071069be;
assign Ia6d61947d36fc128c689808c82db80f6             = conv_qin_00080_00003;
assign conv_Sgntin_row_00081_00000 = I98febac90cccb5fc1f3d966b6e38c4d3;
assign Ief5cbddfbfb98fce4812a676849b9a98             = conv_qin_00081_00000;
assign conv_Sgntin_row_00081_00001 = I0038305f94aaefe2cd1a243580d95932;
assign I3ca2b9b77ed8d78a10aff42a07a53b07             = conv_qin_00081_00001;
assign conv_Sgntin_row_00081_00002 = I0d41bef808860bde56d48792764612d5;
assign Ic5467e42aa377c6ffd8f70673808774f             = conv_qin_00081_00002;
assign conv_Sgntin_row_00081_00003 = I373be7c3f9511a2906584e33e5048abf;
assign Ie9b042f686381739b9ff219041f1e0ce             = conv_qin_00081_00003;
assign conv_Sgntin_row_00082_00000 = I2c8f4a147b363d9c5ef0e080d9a9ed40;
assign I694d471fd353eb54aae08a2afa7b645a             = conv_qin_00082_00000;
assign conv_Sgntin_row_00082_00001 = I9171019227f35760d02d0c8ce786f4d3;
assign I15fafe2baba4d2f28037023a81ce0a81             = conv_qin_00082_00001;
assign conv_Sgntin_row_00082_00002 = I669d34b955d2991ebbb31c149ad1b6f8;
assign I1c85a2d1df6749a194072eb731506bfe             = conv_qin_00082_00002;
assign conv_Sgntin_row_00082_00003 = Ie0b5f51835ebdb508a596eeebf0e4847;
assign I0c4268c01aed70ce4fc71531bf4bb862             = conv_qin_00082_00003;
assign conv_Sgntin_row_00083_00000 = Ie644d131c4f2c603e8e64c5581fdf822;
assign I7d4924388dc5373ad7936dca76797473             = conv_qin_00083_00000;
assign conv_Sgntin_row_00083_00001 = Ib70e99c3acc76286a6811bcacc9284de;
assign Ifa43d74fa91b7b9884969f575ef9ca8e             = conv_qin_00083_00001;
assign conv_Sgntin_row_00083_00002 = I263aad78110a1136eb7012c6983b2a8d;
assign I3ee10f6a7785a236db317515fdd23a2d             = conv_qin_00083_00002;
assign conv_Sgntin_row_00083_00003 = Iddb75e0197b9a76b36a59ac2a7ccdf3a;
assign Ia34e42f8de91fa4861b0c6cac5dcfc29             = conv_qin_00083_00003;
assign conv_Sgntin_row_00084_00000 = I8e873fb2321eea82bb590a92411e2e2c;
assign I46894c6526983bf1ce4b503159131b41             = conv_qin_00084_00000;
assign conv_Sgntin_row_00084_00001 = I6cde57127c5bd2732e71ecb7738fad6d;
assign Icb82c9ff4cb58159a1c3115c6fdd5f8c             = conv_qin_00084_00001;
assign conv_Sgntin_row_00084_00002 = Iae6ed7748692f2edf1aa9d73380075f0;
assign I3ec5819176ad4b0895a9118d90ab22b5             = conv_qin_00084_00002;
assign conv_Sgntin_row_00084_00003 = I08c03198b9599b2f4590e3022e398f7c;
assign Ib7c5850b4f7cc77be2048d114a2128d9             = conv_qin_00084_00003;
assign conv_Sgntin_row_00085_00000 = Ia62832d325f86160285c4d1a790a32cb;
assign I4fbdc4ee57a3be42b62d9bd43078d6ef             = conv_qin_00085_00000;
assign conv_Sgntin_row_00085_00001 = I2f23d4cdb6f5f827513aa60266936e4f;
assign Ib3367565e4456da15e7c2315dccdb5e4             = conv_qin_00085_00001;
assign conv_Sgntin_row_00085_00002 = I4b99891bed4f5c149cd4a5b4f1dde0f0;
assign I4accbad1b451ed2b622e15ef9ae16d13             = conv_qin_00085_00002;
assign conv_Sgntin_row_00085_00003 = Ia4f3cff223e24815ee1d86bf41756f06;
assign I32bb50faa2b246b2d3b462a79be597c5             = conv_qin_00085_00003;
assign conv_Sgntin_row_00086_00000 = Ice82cfe55a5f226746e59e5c8beb46be;
assign I33bddb0adcc2af7b12a83bf843036385             = conv_qin_00086_00000;
assign conv_Sgntin_row_00086_00001 = I09031235f61238b0e32ff52641aab70e;
assign I2c926fd9d306e9ae13364e07c4b0395b             = conv_qin_00086_00001;
assign conv_Sgntin_row_00086_00002 = I9d7614d286377329eb3999213889b707;
assign I8e517c401d62dbb10dcc96ab536f6afb             = conv_qin_00086_00002;
assign conv_Sgntin_row_00086_00003 = I56592e1452c4b559af19465b30230ec0;
assign Idc6d40a49f05c5422758cee50f787eb1             = conv_qin_00086_00003;
assign conv_Sgntin_row_00087_00000 = I384d5377ee6b8f7eb2db23a2e444ddbc;
assign Ia6308e16fae5428f4ab6560f5b21479a             = conv_qin_00087_00000;
assign conv_Sgntin_row_00087_00001 = I477a920e2326828bf026b0a6b6a18e2b;
assign I448f126fd3932d5065abbe7bb2d92c56             = conv_qin_00087_00001;
assign conv_Sgntin_row_00087_00002 = I5196382b75d16892d550f17893de15ec;
assign I960768a84aec9d5b8bc7c1c523024a25             = conv_qin_00087_00002;
assign conv_Sgntin_row_00087_00003 = I213ce488e5345fa405a9c5df297d6f74;
assign Ide1d7dc22a4b271ef764df14ac22366a             = conv_qin_00087_00003;
assign conv_Sgntin_row_00088_00000 = I5ad7eb9d3ce7c712515254f892d1670d;
assign Id9364a29fd79b52d0442e18dc0227854             = conv_qin_00088_00000;
assign conv_Sgntin_row_00088_00001 = I914dedc1d5e5e21c9b8d07ec0ecc01f9;
assign I2b2bd845428c49346ef8e94e95b618f8             = conv_qin_00088_00001;
assign conv_Sgntin_row_00088_00002 = Iefac1e428116a797c2c0803410ac5601;
assign I7ace6778ac86b3e05939a3fcc716136f             = conv_qin_00088_00002;
assign conv_Sgntin_row_00089_00000 = Ib534288c2cf976b6ec85db743bc2a823;
assign Id113cab2dd1949d32e3c1c15273185c8             = conv_qin_00089_00000;
assign conv_Sgntin_row_00089_00001 = I90023493600924a76d2192080cf6194e;
assign I103f1449c78c47396d6a54dc1c810934             = conv_qin_00089_00001;
assign conv_Sgntin_row_00089_00002 = I8b419d5827e5b1af9649d602401c189a;
assign I044e01e8d2df46e03f00a0af2beb0bf5             = conv_qin_00089_00002;
assign conv_Sgntin_row_00090_00000 = I485f9d1104a965d5d035feef912a2ca8;
assign I816704585ad393f685731104ad3ec64f             = conv_qin_00090_00000;
assign conv_Sgntin_row_00090_00001 = I474f6bd977f4197742d0bddb3bece684;
assign I53121a39de0bcba91a4d0438be2ae958             = conv_qin_00090_00001;
assign conv_Sgntin_row_00090_00002 = Ie989550c9101de382056dd60d5da0e01;
assign I45a7ddcda2662e36b7617dfe64514346             = conv_qin_00090_00002;
assign conv_Sgntin_row_00091_00000 = I9b76f0121a3f7e887e7121db50024ab4;
assign Ie317e5ea2ca4ba2060d0f491290af96f             = conv_qin_00091_00000;
assign conv_Sgntin_row_00091_00001 = Ic3fb524ab434e80b3289c9241b65d224;
assign I58703e8b6d04f8c69ac38f5fcfdc4efc             = conv_qin_00091_00001;
assign conv_Sgntin_row_00091_00002 = I259010e323e1e8dcd9dd719091131f6c;
assign Idada779a1ac7b844867571d77054b657             = conv_qin_00091_00002;
assign conv_Sgntin_row_00092_00000 = I30d615203b697787ead37394953925cc;
assign I5ea02b5349cd4d99ccbcb6b26f0cfdd7             = conv_qin_00092_00000;
assign conv_Sgntin_row_00092_00001 = Ic9146d8b3dd0c612073b70b8a8791e8c;
assign I30b0b1d54912c1a41a02a25ab238bb54             = conv_qin_00092_00001;
assign conv_Sgntin_row_00092_00002 = I3e0b41bee4c76eb5f3340ad23bfa01ad;
assign Iee6da3120d73373627b25ab7c0dedd28             = conv_qin_00092_00002;
assign conv_Sgntin_row_00092_00003 = I389ac86954fd70464c9550e3fed4ed33;
assign Ieeba01b18a244ab8c0ac263c138fabcc             = conv_qin_00092_00003;
assign conv_Sgntin_row_00093_00000 = If4cb744ee52b6ae793431cd038069b57;
assign I6404d0df952b5bf8292c753e4c6f35d8             = conv_qin_00093_00000;
assign conv_Sgntin_row_00093_00001 = Ic3cb34aae74c5f1a870b3635f8a40764;
assign I913d818403024510c55b65b56a38dd89             = conv_qin_00093_00001;
assign conv_Sgntin_row_00093_00002 = I877e8d94236c3d8b0a31858a98fba5d6;
assign Iadf927d18644a232ad1f1eba7db82934             = conv_qin_00093_00002;
assign conv_Sgntin_row_00093_00003 = I77371f0e55b4684d1af196ed52d3d997;
assign Ie4c9797a955778694dd8615219cb51e7             = conv_qin_00093_00003;
assign conv_Sgntin_row_00094_00000 = I83c7d177eec2dad0a924557cdc91ba77;
assign I5510b88bfd65811b3200adf4ef975b48             = conv_qin_00094_00000;
assign conv_Sgntin_row_00094_00001 = Ib1073489d63ea33d7f3892f4ff875358;
assign I7774313f1ae5a2de98855aad572b3676             = conv_qin_00094_00001;
assign conv_Sgntin_row_00094_00002 = Ieefbb5d6f4ac1e586832c5c0f513c5a2;
assign I46ee30b46020d91707689f3468f00e26             = conv_qin_00094_00002;
assign conv_Sgntin_row_00094_00003 = I5a21996f5724a2a49fcf8e928c01b062;
assign I28a5ed4c239e64c76bb6e566b50cfd23             = conv_qin_00094_00003;
assign conv_Sgntin_row_00095_00000 = Iea1297491d1dfe98f395d8c73808a893;
assign I529f92b82248efe2cf64f7da0ec8283c             = conv_qin_00095_00000;
assign conv_Sgntin_row_00095_00001 = Ie9236599cea94cfb603c6b977fdbb44a;
assign I7846bc2cc11e08d05f7c853c4920d555             = conv_qin_00095_00001;
assign conv_Sgntin_row_00095_00002 = If8fe5af7e5c3c97b5a713f6bcf919f1f;
assign I7607af5d98e8070e3d15cee23cdf877e             = conv_qin_00095_00002;
assign conv_Sgntin_row_00095_00003 = Id46108963921efa50aff64d4dd7d1701;
assign I79a705ee1e414fe4a5fb14e9b3ce9597             = conv_qin_00095_00003;
assign conv_Sgntin_row_00096_00000 = Ife25829fb3c5023b7d69bbaadf9cf77e;
assign Ica3a41ace27f7d94377981079952f4f7             = conv_qin_00096_00000;
assign conv_Sgntin_row_00096_00001 = I3375fff5ee0d4b4b12c5a70fbdee59fe;
assign Ib730fdb59198f23d1e590f6d6039e96a             = conv_qin_00096_00001;
assign conv_Sgntin_row_00096_00002 = I68c35d63dc95baff41b4dc27a86d2342;
assign I31243de90dc2a1656ca9d5e03bdd78da             = conv_qin_00096_00002;
assign conv_Sgntin_row_00096_00003 = I8da50e5093acefb6f809aed64564a53e;
assign I04f90a907f10a7fa1ae3591b48094d5c             = conv_qin_00096_00003;
assign conv_Sgntin_row_00097_00000 = If988b82b86db1f4ff6d3695f7b0197e4;
assign Icfe1a689e33b2b9aa9dba692d6d610b9             = conv_qin_00097_00000;
assign conv_Sgntin_row_00097_00001 = Ia9f5ce4603af279bbd9b486b67016482;
assign I56b3a97dc3037f0bb2eed93a9482c813             = conv_qin_00097_00001;
assign conv_Sgntin_row_00097_00002 = I0c5539373b3868d0664a92157b4b4226;
assign I282d2eb4e74e034694e33273b9cb19d5             = conv_qin_00097_00002;
assign conv_Sgntin_row_00097_00003 = I03b0694777d0160a83cbc82ac1397736;
assign I31d25b1b49e65216e90b39aa27acd6be             = conv_qin_00097_00003;
assign conv_Sgntin_row_00098_00000 = I10fca5f2cbf5e2bc3433c0dda579a051;
assign I85d95015a9ce27a18ccbf73bbbcdbd70             = conv_qin_00098_00000;
assign conv_Sgntin_row_00098_00001 = Iaa1e981134f5a5c02983c49562683bc5;
assign Iff7950f24f0a6b0073942c37fff49d37             = conv_qin_00098_00001;
assign conv_Sgntin_row_00098_00002 = I6eea5fde8e2517554ad6ba25018572dc;
assign I6072331f838d82329a07a4ffa340c7b6             = conv_qin_00098_00002;
assign conv_Sgntin_row_00098_00003 = I85c2bffb93569d9fe1b1bcb10b98bcac;
assign I1f6540c5f037d861dee2c0091cba01ec             = conv_qin_00098_00003;
assign conv_Sgntin_row_00099_00000 = I9eaf4e9ebe07717503ff69b51f0e1905;
assign I56ea52c50a188ec47e48740839a031c9             = conv_qin_00099_00000;
assign conv_Sgntin_row_00099_00001 = I23c8b64e433af0bd00cef44e38df99f8;
assign Ie1f41720e296ced1b74cb325b666d88f             = conv_qin_00099_00001;
assign conv_Sgntin_row_00099_00002 = I7bfb4c5d9e22d1bd8811844d9c74dff8;
assign Ib3a0307176d424a4733720416d71069d             = conv_qin_00099_00002;
assign conv_Sgntin_row_00099_00003 = Id00274c88b93867a80606343add1cdab;
assign I9632bb500b7faaaaeb649d74c21cbe8c             = conv_qin_00099_00003;
assign conv_Sgntin_row_00100_00000 = I7741e239c16828889d488cc87647c154;
assign I8522c402e654d007abffcb0e904af5e6             = conv_qin_00100_00000;
assign conv_Sgntin_row_00100_00001 = Ic828cdd5dfde844df4c150921af2a443;
assign I2605f078c1a9006c93855a9a2b0cf6b9             = conv_qin_00100_00001;
assign conv_Sgntin_row_00100_00002 = I61e829cbf7d6c0ef8ddc11677981e2cf;
assign Idd0217a35c3adc8abc7bb581a5df7a2d             = conv_qin_00100_00002;
assign conv_Sgntin_row_00101_00000 = I7050adb9d06f767549b7f35c4679e391;
assign Ib57ef2f577cca54713c16717cbbd1ce9             = conv_qin_00101_00000;
assign conv_Sgntin_row_00101_00001 = Idc5fb0f3a04ab32948e249e088a11b11;
assign I2e11a697d7f17ac30302eadb500de72d             = conv_qin_00101_00001;
assign conv_Sgntin_row_00101_00002 = I9e8ae2aed048068b01b3bd46f30baae8;
assign Ic05b46168884322644db4e331d37d759             = conv_qin_00101_00002;
assign conv_Sgntin_row_00102_00000 = If43dd31198c8a0da6fabd194cf13bb70;
assign I2f34af0036985cd94ade9cc905bec065             = conv_qin_00102_00000;
assign conv_Sgntin_row_00102_00001 = Ic0732810fd355d59a3168be896a0f9ac;
assign I56fc99a22960232b305d6e683c66fcc7             = conv_qin_00102_00001;
assign conv_Sgntin_row_00102_00002 = I7dab71adbe62687846fc027d2789451d;
assign I53c88dc237bb2cd02d50fd7f0a168a48             = conv_qin_00102_00002;
assign conv_Sgntin_row_00103_00000 = Ib16548d471f0a4f4625852ea04335dcc;
assign I21de4f6194dec9e3c401934db92c25e7             = conv_qin_00103_00000;
assign conv_Sgntin_row_00103_00001 = Iff2f1716cbd73b406d8f07c22dc79fc8;
assign I2a9c673cdd7ded79e09ada38c0f47e6f             = conv_qin_00103_00001;
assign conv_Sgntin_row_00103_00002 = If1295608bd218ed60922a0b95bf1d098;
assign I7450d4ab3ef0227e93a02bfd620d047b             = conv_qin_00103_00002;
assign conv_Sgntin_row_00104_00000 = Ib051eb1091a85f85a1e50007f1b27cab;
assign Ide86f019e9573706c25bd8b4552396a8             = conv_qin_00104_00000;
assign conv_Sgntin_row_00104_00001 = Ibdad0ab78e4404c852e60a2b04c3a5f6;
assign I07b417cdcc99eaea3413f563e26ddc73             = conv_qin_00104_00001;
assign conv_Sgntin_row_00104_00002 = I5fdd8e1550feaecd81b82069fe73ed7e;
assign I8eba6f14f42701d22859fbea94bd1871             = conv_qin_00104_00002;
assign conv_Sgntin_row_00104_00003 = Ib4ae1cedd09d72c235765a6cd7e91366;
assign I49b64469d298012dbb131d879bff38d6             = conv_qin_00104_00003;
assign conv_Sgntin_row_00104_00004 = Idf04e08c120ed116af14a62659675b44;
assign I2b16e5b4e279bb29c3c675b72083e5fe             = conv_qin_00104_00004;
assign conv_Sgntin_row_00105_00000 = If6a5dc79c0f6ce348956286737a369d8;
assign I5d5701435c96f1078e741921b56e3c65             = conv_qin_00105_00000;
assign conv_Sgntin_row_00105_00001 = I6d4fc81ced37c159303c243af04d345e;
assign I761983331fb6e3c6c437b3f1660f0b6b             = conv_qin_00105_00001;
assign conv_Sgntin_row_00105_00002 = Iba1c0ebd9cefeb0dd7f690bdbbbfec58;
assign If7f373506cac70f8ba1222db135c27e8             = conv_qin_00105_00002;
assign conv_Sgntin_row_00105_00003 = I3472ee8c06644490252e606b62bf9bd5;
assign I5ce8b2f633011e89356243a1a71edeb6             = conv_qin_00105_00003;
assign conv_Sgntin_row_00105_00004 = Ieb7614ad1b1bfed3e2b0089a72fe214a;
assign I70c92e8ada46476d15ef4b3c620d2601             = conv_qin_00105_00004;
assign conv_Sgntin_row_00106_00000 = Ia8e304ca12c82e41cb8e4de7be199394;
assign I644e83f0a7d432fba38ffb2d99088eca             = conv_qin_00106_00000;
assign conv_Sgntin_row_00106_00001 = Ia2c5fe53cb5b318fa63d09881609655f;
assign I73203143fe37933c16fff873c1abf512             = conv_qin_00106_00001;
assign conv_Sgntin_row_00106_00002 = Ic124975d36a292816146a2fe61ab3ab9;
assign I039f05d5be891a37e04556f1eae674d2             = conv_qin_00106_00002;
assign conv_Sgntin_row_00106_00003 = I3eab1582cc42db0ac7739386cce2a712;
assign I8ad3627f171eadcc960a688ac0afcbc0             = conv_qin_00106_00003;
assign conv_Sgntin_row_00106_00004 = I589062eca318b25dfe5735da455b6fe1;
assign Ib193b07804d6d5f111b06bda487bfa5f             = conv_qin_00106_00004;
assign conv_Sgntin_row_00107_00000 = I05721e06a1acdcc0571907c7d853f18c;
assign I51e98035b35a35fdc52f5bab8f19c152             = conv_qin_00107_00000;
assign conv_Sgntin_row_00107_00001 = I1e93f0470d2818249f1c28ef2a399a0e;
assign Idcada1bfb3c0d1f2a09aab58a2071a57             = conv_qin_00107_00001;
assign conv_Sgntin_row_00107_00002 = I453dd7d7c0a2f003f0b67e909630d641;
assign I94c4e11670b4233fa072517a8f19c901             = conv_qin_00107_00002;
assign conv_Sgntin_row_00107_00003 = I6387919f2426c283e2d70e471cda54a6;
assign I09b5273bb15d48a7fd78559930fa6d1c             = conv_qin_00107_00003;
assign conv_Sgntin_row_00107_00004 = If3db87afb3ea184c9e4020c5e45cb161;
assign I885433b0ab16c6d87abe45af13c9e529             = conv_qin_00107_00004;
assign conv_Sgntin_row_00108_00000 = I7979161aa1e2262ebea862004c387697;
assign I5ed85845c39337c37791f16e718069b4             = conv_qin_00108_00000;
assign conv_Sgntin_row_00108_00001 = Iaddc1f2e822fd2fe9d9046d759a82cb4;
assign I1cd93172cf5996bc870063aa642188a2             = conv_qin_00108_00001;
assign conv_Sgntin_row_00108_00002 = Ia14bc1fcd5bbdcb60b8e68298f7d716a;
assign I198c055930cb89d0390c336eda8fed4f             = conv_qin_00108_00002;
assign conv_Sgntin_row_00109_00000 = I04aacd95d9e44657f616e01c9053f0fb;
assign I15943aa74e9fbbaebdc0d54eb6a3bffa             = conv_qin_00109_00000;
assign conv_Sgntin_row_00109_00001 = Ia8974083bfd064f2c27dcd421490fcfd;
assign Ifb00ae47340bc99669c71da34cccc59e             = conv_qin_00109_00001;
assign conv_Sgntin_row_00109_00002 = I268b60cb371b3d46dc3f8b0009f541b1;
assign I688a2c72e69b217d2673e8da75146a83             = conv_qin_00109_00002;
assign conv_Sgntin_row_00110_00000 = Ibeb8c72b90b50c6897224ca1a792fa56;
assign Ia1a0d8d7dfd6e877f15cce773f85f5b7             = conv_qin_00110_00000;
assign conv_Sgntin_row_00110_00001 = Ie232799bd6c4ec99e24c78f3ad798265;
assign Id4451722e8e2393d627dcd0175dc9903             = conv_qin_00110_00001;
assign conv_Sgntin_row_00110_00002 = If2cd93b57cd1c2b91ee7a73a97dd19f2;
assign I3b6fde4ed14cd68af1468ae1d4cc1a22             = conv_qin_00110_00002;
assign conv_Sgntin_row_00111_00000 = I0987c561670b7b2b6683303c1be39561;
assign I57d0920119f8901bd4dea2d5f8fb5d90             = conv_qin_00111_00000;
assign conv_Sgntin_row_00111_00001 = I3b30b4ab00a49e10a75587aa324d6132;
assign I80a89644e278e96b1cd1c4b7f764dc34             = conv_qin_00111_00001;
assign conv_Sgntin_row_00111_00002 = Id81305359a07db527e49fda05cd2784f;
assign I5d3df1e7563630311f56143ee6d97a8e             = conv_qin_00111_00002;
assign conv_Sgntin_row_00112_00000 = I8b2a79aa4ac88e6b4ca8188a7852022e;
assign Ib57795a63d642a73456324bab41384b6             = conv_qin_00112_00000;
assign conv_Sgntin_row_00112_00001 = I6b5645cdde4b35a16fe3e91d90caaa4e;
assign I2370042234b0e93bb66e44b97fca3e43             = conv_qin_00112_00001;
assign conv_Sgntin_row_00112_00002 = Ibc48fabc172f27ebce18d0a9b5120dc5;
assign Ia86740e870d8063f0266b68ad6d7481d             = conv_qin_00112_00002;
assign conv_Sgntin_row_00112_00003 = Id8292eca087c1a17dc8b5a572a76f21f;
assign I90a7ea789d3bf7f9126c786474a56da0             = conv_qin_00112_00003;
assign conv_Sgntin_row_00113_00000 = I6ef260ef75e47b011a46ba2080ac3684;
assign Ia4b671f3360f3ce55db0dc0e4d78ddbe             = conv_qin_00113_00000;
assign conv_Sgntin_row_00113_00001 = I34e6e9d2153e4a70ee36ab85e72d5318;
assign Id96e744d9b10dcddd1ae0115ea57a76a             = conv_qin_00113_00001;
assign conv_Sgntin_row_00113_00002 = Idf1ecab26889c4adcb835fda6b1cb368;
assign I4d226dd2f0bfcdbea6a2e6a6613c1b64             = conv_qin_00113_00002;
assign conv_Sgntin_row_00113_00003 = Iddb19725b093506e5e521d8d68dcb8e1;
assign I5029424c9d9fe923eeb858b1e62cd758             = conv_qin_00113_00003;
assign conv_Sgntin_row_00114_00000 = If8572800d5d80cc92dd917b60447b63b;
assign I992e7c551b4aa818606c3465d33eb798             = conv_qin_00114_00000;
assign conv_Sgntin_row_00114_00001 = I3566f2779e860008b1a5d305366a07c9;
assign I97f2b15ce0a74e68d5a4438111adcb0a             = conv_qin_00114_00001;
assign conv_Sgntin_row_00114_00002 = Ia9f1e580e8f441394d719d52a7bad688;
assign Ia0886ce792e062e22d0c224158cdfb7d             = conv_qin_00114_00002;
assign conv_Sgntin_row_00114_00003 = I0b573d3a86a3111451da661e46384876;
assign I1e805c70d50c2765b4a03ad2982dc421             = conv_qin_00114_00003;
assign conv_Sgntin_row_00115_00000 = Icb0841ecf142687c3aa23e68f01c927c;
assign Id9b9a8fe43992ec0793845715dd2226c             = conv_qin_00115_00000;
assign conv_Sgntin_row_00115_00001 = Ibfcfd3151af0d82bfce293ada44059b3;
assign Ia6a7f9beaceb08d81012f0e72171252f             = conv_qin_00115_00001;
assign conv_Sgntin_row_00115_00002 = I220e32641265b46527ca61111f7ebf1b;
assign I0a9a09b0ab43d2a0f1d1d01e13f0333c             = conv_qin_00115_00002;
assign conv_Sgntin_row_00115_00003 = I0ff479e61d1a0cede88ebffb073c60be;
assign Iba58175a7fd5c5da650222193caff0b3             = conv_qin_00115_00003;
assign conv_Sgntin_row_00116_00000 = I8e87530a131b5a73cad6df68b9e4967f;
assign I5dd29fd1a73df5662d2b636e7285bad9             = conv_qin_00116_00000;
assign conv_Sgntin_row_00116_00001 = Iee17ece482d04964d3c21a092ec955a4;
assign I7c19a79f441ecbb73685db5a505e7479             = conv_qin_00116_00001;
assign conv_Sgntin_row_00116_00002 = Icd6f8f5df6b4ca4c81855e974db76526;
assign I7401a0501ba69c5559fbf00c77e58dc5             = conv_qin_00116_00002;
assign conv_Sgntin_row_00117_00000 = I2bdf4736022e5da7294a0e851006a124;
assign I89537301987d6da0dbe6cff3caab3ff4             = conv_qin_00117_00000;
assign conv_Sgntin_row_00117_00001 = I1c7e41b9cb1bdb6f649c88c0ed3f4100;
assign I9aaa036a6158d11c235bdc8406d79f4c             = conv_qin_00117_00001;
assign conv_Sgntin_row_00117_00002 = I7ce064a756dad56d37684d5d7d168047;
assign Idd9f7ea657ea9cdcb45a7e4b573b9d50             = conv_qin_00117_00002;
assign conv_Sgntin_row_00118_00000 = Ic62fc602da3d16fe13d03a49a21269d0;
assign I89013d61c1ea8da8b1c6071cc21c316f             = conv_qin_00118_00000;
assign conv_Sgntin_row_00118_00001 = I5364deb983adc2ae505ed2b8c57f876d;
assign I1f00849ea055a7893df386aed162a7b6             = conv_qin_00118_00001;
assign conv_Sgntin_row_00118_00002 = Ied2ea62cfb21602645babc36e27b8218;
assign I53f275395dd6be17961a5edc3e8da7f2             = conv_qin_00118_00002;
assign conv_Sgntin_row_00119_00000 = I2ff317d57f59747c4524ef4278d51092;
assign I6ac24c46319a787daa5c545de8c6eeea             = conv_qin_00119_00000;
assign conv_Sgntin_row_00119_00001 = I6e92a48aaab94074a555efa9bd1e7243;
assign If4d5b48882e9e628cf51ad2ac2f38c22             = conv_qin_00119_00001;
assign conv_Sgntin_row_00119_00002 = I79b85da6e5ce0b02ebd1619115c98e24;
assign Icab010d78cd66b02e089c74f04bf4e75             = conv_qin_00119_00002;
assign conv_Sgntin_row_00120_00000 = Ie68b31360c12a83c6095254b6f14603c;
assign I84c88b631bed5311cb6e99e58941149e             = conv_qin_00120_00000;
assign conv_Sgntin_row_00120_00001 = I00d3f14b20e1ea7d726533386e0eba27;
assign I5c942076b173cf527e1be2ddb8560e84             = conv_qin_00120_00001;
assign conv_Sgntin_row_00120_00002 = I579c7926e7b78f4ffc606adc10522f53;
assign Ibed2a63af723a7abf96dacf1951e5266             = conv_qin_00120_00002;
assign conv_Sgntin_row_00120_00003 = I837183265ee22d080e81fea468ab0887;
assign I242a30bdc8699d8ff550b25dd53d6c59             = conv_qin_00120_00003;
assign conv_Sgntin_row_00120_00004 = I8e1ddd7e4185c28caa71d30bc28138f3;
assign I376a48b7e0195a5aacc76a0ad8bd14b2             = conv_qin_00120_00004;
assign conv_Sgntin_row_00121_00000 = I9539fcc40d26b13015a864718b116d5b;
assign I21b062856ced09cb9131c01b5e166f32             = conv_qin_00121_00000;
assign conv_Sgntin_row_00121_00001 = I02849282dd1bd663fd39baccf41762f9;
assign I6b3cd79aa87235ff174c0299b855dd3d             = conv_qin_00121_00001;
assign conv_Sgntin_row_00121_00002 = I5d6e576b0fa7e3219aaf9ccc345085b8;
assign I814b62120953991f9da055f118967e05             = conv_qin_00121_00002;
assign conv_Sgntin_row_00121_00003 = Ic0191941cb968bbd7644c21767423d2e;
assign I3f33901c407a87e10d86c13c83dd52eb             = conv_qin_00121_00003;
assign conv_Sgntin_row_00121_00004 = Iab0bff1633e2f3ea0bfbc291f3ab5d29;
assign I241622b0367dde514f96ece55c8c3964             = conv_qin_00121_00004;
assign conv_Sgntin_row_00122_00000 = I8850ab26807dcd55fefadf6310729ca7;
assign If9efe7a1c359ec03014a52870ac13aec             = conv_qin_00122_00000;
assign conv_Sgntin_row_00122_00001 = Ice59d2af73d0b0f2ae91a2ef0c2b7f04;
assign Ibc73d07e0c97a6fcae791e04106cb082             = conv_qin_00122_00001;
assign conv_Sgntin_row_00122_00002 = Ic4efba3932e598784f5b9ad6ad04772d;
assign I2f3ab9654e515a54e22e73d6c130ccc3             = conv_qin_00122_00002;
assign conv_Sgntin_row_00122_00003 = I9ad2f6fd2d7f68011fc926ec9abd5c34;
assign Idf6875955525d80dc660ce956f4a84e7             = conv_qin_00122_00003;
assign conv_Sgntin_row_00122_00004 = I5f0751fceaa008feba5c6867ced453dc;
assign If94a1abfb972f63629d07e64dc23863c             = conv_qin_00122_00004;
assign conv_Sgntin_row_00123_00000 = Ifdabf743a8cb46b7053000ff48ea0c60;
assign I0c0060fe260afa3cdc72f35ffb6938ff             = conv_qin_00123_00000;
assign conv_Sgntin_row_00123_00001 = Ie562ebb336e476a81f20a652d4cb20f1;
assign I6627bcdbaa8afb115123777abd45435b             = conv_qin_00123_00001;
assign conv_Sgntin_row_00123_00002 = Iefdb8bd28839af9413a3906cbfe715e6;
assign I70d32affde22f9dcb2d77430fca39069             = conv_qin_00123_00002;
assign conv_Sgntin_row_00123_00003 = Ib9d58222da98f29fa302b4896594fe26;
assign I76060709de3ea188748849f043c59ac0             = conv_qin_00123_00003;
assign conv_Sgntin_row_00123_00004 = I9f6751c15237c20b0cf2175575195ea7;
assign I07b9b1f4fa01b16cc69356057d3b6154             = conv_qin_00123_00004;
assign conv_Sgntin_row_00124_00000 = I081e2595b18f306a74d070203447ecf6;
assign Iabf572c97b48c6a7dcc19e56676e3a82             = conv_qin_00124_00000;
assign conv_Sgntin_row_00124_00001 = I3b84dad6d0dd8730312b3e20c6d5a2a8;
assign I5814a85c45fd0f7be21ed325235fe4b7             = conv_qin_00124_00001;
assign conv_Sgntin_row_00124_00002 = I6ea50be10bc990a1206cdc9e28e0c4c2;
assign I2288a6ad3b748b716249f4adc42d52c4             = conv_qin_00124_00002;
assign conv_Sgntin_row_00125_00000 = Ifc1da524e7670772834d521a6fc4c96f;
assign I60cbd4369e7ba9b6532f279e5c59084c             = conv_qin_00125_00000;
assign conv_Sgntin_row_00125_00001 = Ie2d946edaddd3c87f328e861f3e72c0a;
assign I95361d5f524ccb9feb42811af5c482e2             = conv_qin_00125_00001;
assign conv_Sgntin_row_00125_00002 = I43c2fab87f70ea883321ab82de85f133;
assign I022df337bcc05ac5648b8ae2e42f3a76             = conv_qin_00125_00002;
assign conv_Sgntin_row_00126_00000 = I24645082ef16129eed1c574f5fc601ca;
assign I2ead0e9941e2280309ab53535b1e1ac1             = conv_qin_00126_00000;
assign conv_Sgntin_row_00126_00001 = Idb1efe99b5d7fd567a7f82cfd52f7eb8;
assign I3e5139f24e3d082eb31b0e61ea9fa1aa             = conv_qin_00126_00001;
assign conv_Sgntin_row_00126_00002 = I1af02ed6cf00d4cb0704b5e44c83bfa3;
assign I60d9a7f95fb8623753002ecaf9a4efcc             = conv_qin_00126_00002;
assign conv_Sgntin_row_00127_00000 = Ie8c0fac00a9de74870e59cbf9e87a39b;
assign I93b69bfb228db4b569a6772179d603be             = conv_qin_00127_00000;
assign conv_Sgntin_row_00127_00001 = Ie4827dc0983c1a63053c08de6e36d375;
assign I85c4d3d6c8408c6f38741257ed177ca6             = conv_qin_00127_00001;
assign conv_Sgntin_row_00127_00002 = Ib71611afdd0381cc1884f5ddbbae1acc;
assign I23a74ea5e7174d95e6d16a5e85ac236b             = conv_qin_00127_00002;
assign conv_Sgntin_row_00128_00000 = Idf8d15c7bd7705b9aafbda09c3a5b46c;
assign Ide530e6f4622c8a7b101b6dce9650e42             = conv_qin_00128_00000;
assign conv_Sgntin_row_00128_00001 = I7f720a18542528f0c9bfb14f699ff4da;
assign Ic95191bccb18e26c10e56be395ca6b1a             = conv_qin_00128_00001;
assign conv_Sgntin_row_00128_00002 = I70a4926e9e6a05fa9ee51a26988862fe;
assign Id0f75e19b94541ed5c5c352d13390d2d             = conv_qin_00128_00002;
assign conv_Sgntin_row_00128_00003 = I38fc49afce0298846ae8ed63ae715e81;
assign Ie697d28d757df82b3901564bda43251c             = conv_qin_00128_00003;
assign conv_Sgntin_row_00129_00000 = Ic6fd9592d2ffcb8f4ca83c6f0bd19975;
assign Iaf0bbbe791bb71d0f557dc71caa5fb87             = conv_qin_00129_00000;
assign conv_Sgntin_row_00129_00001 = Ie4cda4648f6ceb76b8fb74f290ab6439;
assign Ie4ae993ddb776bdffec843db0def2f5c             = conv_qin_00129_00001;
assign conv_Sgntin_row_00129_00002 = I5707d30ca29842b6a96cfaeb44ac6668;
assign I4dca2dd40a7127ce44f83b430a34c738             = conv_qin_00129_00002;
assign conv_Sgntin_row_00129_00003 = Iddc3e44d83e8253e5129b6cbf5082df7;
assign I8572aedc94f7243ce5eacb332c81eae2             = conv_qin_00129_00003;
assign conv_Sgntin_row_00130_00000 = I94009bb7239be96243902ab0f0abea7e;
assign I4102100fa5f1dd299af0190862efcc42             = conv_qin_00130_00000;
assign conv_Sgntin_row_00130_00001 = Ic308610ea8bb62ecb6094192e02dbdba;
assign I224bbdf94ac86c5c376d1db4f4d4e060             = conv_qin_00130_00001;
assign conv_Sgntin_row_00130_00002 = I85654bd3a07b4329aba17d8b27777f4e;
assign I6d83efa9f988328f487e9232bf2633a2             = conv_qin_00130_00002;
assign conv_Sgntin_row_00130_00003 = I975a87bdda30c5b6be8d2f0e4b107450;
assign I6734123aaf6320da75638b212812732f             = conv_qin_00130_00003;
assign conv_Sgntin_row_00131_00000 = I8bd2a9d90074500698b302cb8db7f03a;
assign I52403a0454e5fa002e79eaab7ea497bd             = conv_qin_00131_00000;
assign conv_Sgntin_row_00131_00001 = Ib5ee5a6ffc45ed1fece0822dc4619b57;
assign I96fe3eb633eff6958ac575b997460bb9             = conv_qin_00131_00001;
assign conv_Sgntin_row_00131_00002 = I235c3a9fd3e8ea1cee762c10bc8e2c53;
assign I69f563e7b7ad483893ac9c4684349769             = conv_qin_00131_00002;
assign conv_Sgntin_row_00131_00003 = I582bd96afa764ded148202f738b7a1df;
assign I7f6dc6f0f403c58f9aaaa70c2383a666             = conv_qin_00131_00003;
assign conv_Sgntin_row_00132_00000 = I5490039998187a1a2efc3549e3dee7d6;
assign I4f1221ce7880729fe584b42ef3afe6b2             = conv_qin_00132_00000;
assign conv_Sgntin_row_00132_00001 = I0615acb0f7cf79b5f6ae8e91cb525dc9;
assign Ic08e85346f61da036a15345a13ac12f0             = conv_qin_00132_00001;
assign conv_Sgntin_row_00132_00002 = I7ec15b73b2811b44e1e50c74a9f921e9;
assign I9160d11439c5140c0109b5190eb82e6b             = conv_qin_00132_00002;
assign conv_Sgntin_row_00132_00003 = I6fb88d97bc9ed37a06b729020a1df140;
assign I66391978843c39b6acbdb4847a01050a             = conv_qin_00132_00003;
assign conv_Sgntin_row_00133_00000 = Ic5cb81c821716a8aabf8cc2283ff73ba;
assign I6a6eb62960b616043415406ebfc21346             = conv_qin_00133_00000;
assign conv_Sgntin_row_00133_00001 = Iffa06a336949f56f4e5a88a06d8b7e60;
assign Id667c80003b5541de9f84d3b8709c828             = conv_qin_00133_00001;
assign conv_Sgntin_row_00133_00002 = Ic68f500938d80460ffdb33a0adc48298;
assign Ia030c08757123aae947f86ab8bfb6d94             = conv_qin_00133_00002;
assign conv_Sgntin_row_00133_00003 = I1500943c4a550e78fc169437b0a663b7;
assign I4f756e4125c8af5c412944b273e01cb0             = conv_qin_00133_00003;
assign conv_Sgntin_row_00134_00000 = I22f5bb821a2571d1764978fd76c8f1d0;
assign Iaec1f186cb4a65da21d41e637fc628f7             = conv_qin_00134_00000;
assign conv_Sgntin_row_00134_00001 = Id962beade26396738ba0e97f67d5e261;
assign I123a212546a8ac394051425db4924812             = conv_qin_00134_00001;
assign conv_Sgntin_row_00134_00002 = I7c965c047d862c973d09a81abe03a845;
assign I730634ea15ac94d241f3ad2d6393a227             = conv_qin_00134_00002;
assign conv_Sgntin_row_00134_00003 = I0b83f4ef8ba9badb27e81b32765ec5b6;
assign Id2c9f7ac95de07148c54803f69347f56             = conv_qin_00134_00003;
assign conv_Sgntin_row_00135_00000 = I42ae0c42360c977b35429ce290516a6f;
assign I45c5e6710240685bf54b73b0d7a64271             = conv_qin_00135_00000;
assign conv_Sgntin_row_00135_00001 = Ia03836a4e93d2f36513227d1dfaea0fa;
assign Iebdc41368d57498a04fa73e30b10a966             = conv_qin_00135_00001;
assign conv_Sgntin_row_00135_00002 = I6d423a7d17e05a3c597ec6ef6c5a7cba;
assign I47b878f27c30f79a37e97e022307e9e9             = conv_qin_00135_00002;
assign conv_Sgntin_row_00135_00003 = I2c420acf428e44cdd9ca9998e276f258;
assign I5061e13a179d27e1ba5f89ce8ee0fd4a             = conv_qin_00135_00003;
assign conv_Sgntin_row_00136_00000 = I14bf11ad80890227e47fda26ae1b9c24;
assign Ic7ff9cde71054c1ee9eef81eabdd7061             = conv_qin_00136_00000;
assign conv_Sgntin_row_00136_00001 = Idd474d80b50992537d6f527faf279800;
assign Ia0a02781c674fe5d769206448d475245             = conv_qin_00136_00001;
assign conv_Sgntin_row_00136_00002 = I2eed3d32a27d51036e17c4a21382b4c1;
assign Id66c47fd69c175a4393e975a269cf053             = conv_qin_00136_00002;
assign conv_Sgntin_row_00136_00003 = Ic7b6dae3017b55dd3cd27423d5f1b0ec;
assign I0f7c32fc1548fb49b8041f55c157498a             = conv_qin_00136_00003;
assign conv_Sgntin_row_00137_00000 = Iae7b72abf4d3c536330a229e3836b441;
assign I4939f69abb1eac56d5021e06406a93b5             = conv_qin_00137_00000;
assign conv_Sgntin_row_00137_00001 = Idc5e98f6958786ccf95d39b922b42ea9;
assign Ife1190f76c2e251704c2960c23330a48             = conv_qin_00137_00001;
assign conv_Sgntin_row_00137_00002 = I2a4bbedf880a9a7b4e1bf946f9f96c0e;
assign Ib06b60cf9933dd8952206c5f3ccced8e             = conv_qin_00137_00002;
assign conv_Sgntin_row_00137_00003 = I4a91a7c9b2a0f3552b8f2ef4e2398be2;
assign I89ffab735ee30423c82e079ed98216c5             = conv_qin_00137_00003;
assign conv_Sgntin_row_00138_00000 = I3b8cdfb1440732ce98cd1676e05a2af1;
assign I634f0ce28934600a1a31ab0d8e59b4a9             = conv_qin_00138_00000;
assign conv_Sgntin_row_00138_00001 = I3fbd40faa4c3b78b547b8348c466fd1f;
assign I1a24e98165afa62bd14986911a36fb6e             = conv_qin_00138_00001;
assign conv_Sgntin_row_00138_00002 = Id6b508145cd21ba088ab8fda34577c35;
assign I9c4b34b5fb1d59c132bcaeb6258675df             = conv_qin_00138_00002;
assign conv_Sgntin_row_00138_00003 = I99ff29c7ba68b5d0819f1e1bead51287;
assign I9494921d8487ee0b314f75cf0380fd2f             = conv_qin_00138_00003;
assign conv_Sgntin_row_00139_00000 = I2aea17846a53e2eb2968581ee2c48226;
assign Ibaf00a6780325882067a79f0c4d693d2             = conv_qin_00139_00000;
assign conv_Sgntin_row_00139_00001 = Ibf2a253afde05c905d0b2404c5a808a0;
assign Ic23e01562c8a753fd70c343297be288a             = conv_qin_00139_00001;
assign conv_Sgntin_row_00139_00002 = I24f82a3f2c0e8df486fe495dd95cf8bc;
assign I61cc8a0f49e393721a62a776e4793deb             = conv_qin_00139_00002;
assign conv_Sgntin_row_00139_00003 = If06b00be0356a2be5074d958ddcdb2f9;
assign If2b3e7d1541cbd8ffc2b4cfc3ad13a57             = conv_qin_00139_00003;
assign conv_Sgntin_row_00140_00000 = Iae5d6faac1f5685cb1d400ee2b1d85e0;
assign I71afab29cdb962e1f1ca21b61dfb50c6             = conv_qin_00140_00000;
assign conv_Sgntin_row_00140_00001 = Ia98a6f01e4eb5bc74d50d350e79be426;
assign Ia284f974dd8a526f31eb81ed71a06e94             = conv_qin_00140_00001;
assign conv_Sgntin_row_00140_00002 = Iabb01dc9980b4879a7356712b51df0d6;
assign I3e3ce8b4ead150a6eae2e5c701c7b598             = conv_qin_00140_00002;
assign conv_Sgntin_row_00140_00003 = I604283449f13c7b225ea03f99f2e296a;
assign Idf3d79da44f2d686f5bd43c3c1427430             = conv_qin_00140_00003;
assign conv_Sgntin_row_00141_00000 = I68b152a599887c0039dd9d45c528c219;
assign Iefd370d0df1a93639af482f78a1e8706             = conv_qin_00141_00000;
assign conv_Sgntin_row_00141_00001 = I24135210c23b2422a42c90ee25594191;
assign I3ed2da9b53daac0852a06ad1acfad21b             = conv_qin_00141_00001;
assign conv_Sgntin_row_00141_00002 = If4308ed204e33952c9931f8fe257aca4;
assign I453fdf4fbb5af5bd28a20d7643da9eb2             = conv_qin_00141_00002;
assign conv_Sgntin_row_00141_00003 = I2b600e5f5c146ee97c4044c08e1f5ad5;
assign If8125ad3c9e7f0a2b84106064d320996             = conv_qin_00141_00003;
assign conv_Sgntin_row_00142_00000 = I852d5295a32984af00c95f6d9389555e;
assign Ifb6c65a00d9a2c31d8b1119b949828d8             = conv_qin_00142_00000;
assign conv_Sgntin_row_00142_00001 = I33ee415d85e2bcd8f975d34b880f6ea7;
assign I43f2b69c6b427de3095c44d4166b77cd             = conv_qin_00142_00001;
assign conv_Sgntin_row_00142_00002 = Ifb89e7ad8ef661959d82b7c22f187243;
assign Ie9cce5746a83479a567bbaeac6dbf497             = conv_qin_00142_00002;
assign conv_Sgntin_row_00142_00003 = I9fe16403fc21bb1159a5e0305fd1ef69;
assign Ic9018b88fa91fb638bbab0613795ae13             = conv_qin_00142_00003;
assign conv_Sgntin_row_00143_00000 = I207a0f6184a0b3be71766a8b47ea5535;
assign I56873feb8418005b5661c7382f2dbeec             = conv_qin_00143_00000;
assign conv_Sgntin_row_00143_00001 = I86ba73ee348f80e2f9891d2ebc8a02ed;
assign Iefdcb71f2903b11f5cb0b8857f7a1727             = conv_qin_00143_00001;
assign conv_Sgntin_row_00143_00002 = Ib6ae81df8db1dae269437861ee11ec0d;
assign Ic57eb4a034247a4c952d8224ea9f2bac             = conv_qin_00143_00002;
assign conv_Sgntin_row_00143_00003 = Iabdb9374e5caee281c25b003624b2c4e;
assign Iad4ea0196eb32f9a152c9e6fe5059e46             = conv_qin_00143_00003;
assign conv_Sgntin_row_00144_00000 = Ie5d9cc18b2dd300132470f206452ff17;
assign Iadbd245bf842aebb456417579a3e6296             = conv_qin_00144_00000;
assign conv_Sgntin_row_00144_00001 = I1b695aa715615662eff7065c742b0859;
assign I9c15a6a5c0db11ede80ff6d04c9a56d8             = conv_qin_00144_00001;
assign conv_Sgntin_row_00144_00002 = Id0ab747d92288f23cef793567b2363d1;
assign Ie95f1a7e0effcec0aa423dc803056a13             = conv_qin_00144_00002;
assign conv_Sgntin_row_00144_00003 = Ibd12036702fe60b57354b3aac921559d;
assign Ia8ff29ed728e7f2ae4213f00328b495d             = conv_qin_00144_00003;
assign conv_Sgntin_row_00145_00000 = I671de3d408b5b783541663c7f1e3a6fa;
assign I7103aa739616a39c03e675ea0efb0335             = conv_qin_00145_00000;
assign conv_Sgntin_row_00145_00001 = Ibe01835305315fab50269c72ef849b61;
assign I5827bc87b5db1801b7db16e1e61515db             = conv_qin_00145_00001;
assign conv_Sgntin_row_00145_00002 = I138fb0c48f2d27e3315e237d9e61d653;
assign I5b4305bef5b4350c1d7ae143667afddd             = conv_qin_00145_00002;
assign conv_Sgntin_row_00145_00003 = Ib1639811de6eb1c38257800c201fb704;
assign I70717726200ec02929f679ef05496455             = conv_qin_00145_00003;
assign conv_Sgntin_row_00146_00000 = I169d8f2bb5fde5b202b4239b7a7f1ed5;
assign I16e3559c63ebfed83d6698fc9a9cd93a             = conv_qin_00146_00000;
assign conv_Sgntin_row_00146_00001 = I2b97a79c90f6578c8b2f321f8d598cc8;
assign Ie7f3f1d6cee7f02ae1b17740ed54c049             = conv_qin_00146_00001;
assign conv_Sgntin_row_00146_00002 = Ieed4c810a5bb69de112522dcf00b16ed;
assign If5dfdadb3868ed5a495007362f7db648             = conv_qin_00146_00002;
assign conv_Sgntin_row_00146_00003 = If926d98f659e8fe4bbf36ad2c5c852c5;
assign Iaf1e4c7dae6ad89567836877c08f57d2             = conv_qin_00146_00003;
assign conv_Sgntin_row_00147_00000 = I8ca17b6cf35e1b1f8f601604575d3f27;
assign I88c10c47ae424fbdcb852fbf1e94127c             = conv_qin_00147_00000;
assign conv_Sgntin_row_00147_00001 = I9a6923c6368526a53ef70e16471386ef;
assign I06c7728ef64be8311f48d10d766d0c44             = conv_qin_00147_00001;
assign conv_Sgntin_row_00147_00002 = Iaf82668eb49248709540f2f529f1b3e4;
assign I02cbb4255db2b21ea32140f9e9ddb36b             = conv_qin_00147_00002;
assign conv_Sgntin_row_00147_00003 = I211f8d7f97ebb8eb3e50313513abfb1b;
assign Icd09aa81e9b43528af73e23b2f0f80cb             = conv_qin_00147_00003;
assign conv_Sgntin_row_00148_00000 = I0fd2f706e374a4eb57ee26ab50201e15;
assign I6ff7b86cd7f63f9243646f1be10b2577             = conv_qin_00148_00000;
assign conv_Sgntin_row_00148_00001 = I83ecf12f3b38fc14c3b75e47b71ecc09;
assign Ie631e40caade823a196370fc3358f042             = conv_qin_00148_00001;
assign conv_Sgntin_row_00148_00002 = I304ac9f96945546cdf1b6f1fa7136731;
assign I6ebb2b94f0f80425f8401ae823d92a1d             = conv_qin_00148_00002;
assign conv_Sgntin_row_00149_00000 = If5ae6fbf843fdeee17945bc5ce81aec8;
assign I8c35c5b343b552c22000e194c517ca12             = conv_qin_00149_00000;
assign conv_Sgntin_row_00149_00001 = Ie039ab562e9cf90289047b5425186123;
assign I37dca40506d61bdeab1255ed4892ca20             = conv_qin_00149_00001;
assign conv_Sgntin_row_00149_00002 = I7a9800418bd5c195fc47a72370680b56;
assign I4a2c3204a6a9936d4a215b46c0ffd045             = conv_qin_00149_00002;
assign conv_Sgntin_row_00150_00000 = I9b8023f4dced915cd52c91bc9d4ed78f;
assign Iee367c535d9c39f872d2ec043e7e7b33             = conv_qin_00150_00000;
assign conv_Sgntin_row_00150_00001 = I49d35ec6369de10afb15be8e0cf135c3;
assign I67347c413b5efd8ff9e0d5bc7ab2a047             = conv_qin_00150_00001;
assign conv_Sgntin_row_00150_00002 = I5f6a61c9f0c67510e148e596f553a4d6;
assign Ib02c0694762c4815448b2c8d3df767c2             = conv_qin_00150_00002;
assign conv_Sgntin_row_00151_00000 = I48e3309c61918c3991852b45d9c72ea5;
assign Ie76b0739aec66f8860870e66e87a6445             = conv_qin_00151_00000;
assign conv_Sgntin_row_00151_00001 = Ifa6e3541f5e12bf9677ffc51d0392749;
assign I613d4b1e3b9e812b785c9cf14fefdfe6             = conv_qin_00151_00001;
assign conv_Sgntin_row_00151_00002 = I8e313ceb21359bcc44114ab217b1c394;
assign I98cee6efbbe565d3a4de16703189782f             = conv_qin_00151_00002;
assign conv_Sgntin_row_00152_00000 = I3c0a621dbef864fd1f566bc2e47f32c6;
assign I4a777f0dd62b19dd340ad31517c4e789             = conv_qin_00152_00000;
assign conv_Sgntin_row_00152_00001 = Ie61f299252b8fecfd3e8634b64df5a90;
assign I1e50c90010a3df1a8ce1cff811cc7a0c             = conv_qin_00152_00001;
assign conv_Sgntin_row_00152_00002 = I33ddee677715877c11a1df45cbfb01ac;
assign Ia642db613c0ec1ca4e69afde7a14a839             = conv_qin_00152_00002;
assign conv_Sgntin_row_00152_00003 = I4c9518755c33d725221ad79ee6badba9;
assign Ibf981c01a9d44cbea3c6d8ead92bc2ab             = conv_qin_00152_00003;
assign conv_Sgntin_row_00153_00000 = I5cac08dabbb6de3b01c821d4db93a8e3;
assign Ib6ea4a822da2ea32e0abf6cf8a33d295             = conv_qin_00153_00000;
assign conv_Sgntin_row_00153_00001 = I1e96d5af3d0e3fdce39530dfd0131a7d;
assign I2eb90278aaa54b9c8212b3b4af7c3617             = conv_qin_00153_00001;
assign conv_Sgntin_row_00153_00002 = I373841aa2bcbad8232d54ac9035a3ef9;
assign I45bc13ae0e0554a79c62cd9c6aa8f2a5             = conv_qin_00153_00002;
assign conv_Sgntin_row_00153_00003 = I3c3cffec9f47c9979cb9503f222f370c;
assign I864c33e8ea204d20a9baef4584f22d4e             = conv_qin_00153_00003;
assign conv_Sgntin_row_00154_00000 = Ib62b02ddf0f57bee49838d19783ef6c3;
assign I9905e2686b350e8a6e7f790563a91294             = conv_qin_00154_00000;
assign conv_Sgntin_row_00154_00001 = I182b43872d50de6f7afb700f178b160e;
assign Icc93450a007cee4c0a42717ed7600528             = conv_qin_00154_00001;
assign conv_Sgntin_row_00154_00002 = Iddcfab4a7022e0f12fd20cb34e9b9d02;
assign Ic4a6c02880a9aead7353332708e3f388             = conv_qin_00154_00002;
assign conv_Sgntin_row_00154_00003 = I68d6769541fdc3df321e192f645c667f;
assign I6ad3228e0e2e1f19648d73e83ba5a229             = conv_qin_00154_00003;
assign conv_Sgntin_row_00155_00000 = Id051f1d5454802e0eb37e22248efe8ca;
assign I995d2809ffaf0ecda6a004d01cb9c8c4             = conv_qin_00155_00000;
assign conv_Sgntin_row_00155_00001 = Ib08897f9216599042f7b97b137e07fe1;
assign Idefa29d4d4e2a6e9147f84893520096f             = conv_qin_00155_00001;
assign conv_Sgntin_row_00155_00002 = Id1dce2b9eafc35fa71df33ada4aac539;
assign Ic044d7419cc43736d278c2df33b4a3cc             = conv_qin_00155_00002;
assign conv_Sgntin_row_00155_00003 = Ided55428cbb77f454c2607ac783d7548;
assign Ie099210a99a4899c53baf39559592690             = conv_qin_00155_00003;
assign conv_Sgntin_row_00156_00000 = I275cd09649a750edb8ae8313e4e1e279;
assign Icd2e75e47cab1d539ba9ff1b6e1d7155             = conv_qin_00156_00000;
assign conv_Sgntin_row_00156_00001 = If533578cacb685a95afbb8e1c05d3c07;
assign Ia1ee5579358b564de06c08ca418a9bf4             = conv_qin_00156_00001;
assign conv_Sgntin_row_00156_00002 = I8879df010bbdf6e5fc9370e2fb3289b4;
assign Id3e0c98bff2636e216b4d3a0ffd51054             = conv_qin_00156_00002;
assign conv_Sgntin_row_00156_00003 = Ifd3d4f3e2a388b3c70e7704d6351e0ba;
assign Ieeec71d9df4613555fade2ced7b3baf1             = conv_qin_00156_00003;
assign conv_Sgntin_row_00157_00000 = I7c791c854d0bc28e8dd787545f8fbda0;
assign Ifc8ece44a4e68c3117eda9e65f3084d2             = conv_qin_00157_00000;
assign conv_Sgntin_row_00157_00001 = I90b3708abdf742370f06cc513ee307e1;
assign I65354f2069de0c25bbe7cd50fbe892aa             = conv_qin_00157_00001;
assign conv_Sgntin_row_00157_00002 = I9a403c511fe2d44472ab319a9477199c;
assign Ife1164cad7cda4aa9a08d94dfe86add6             = conv_qin_00157_00002;
assign conv_Sgntin_row_00157_00003 = I17d32f292758416fe02527dfd938fa0d;
assign I4931884e3544af182bcda9061091a42d             = conv_qin_00157_00003;
assign conv_Sgntin_row_00158_00000 = I446857735e680cae93a24dccb59b1924;
assign I0296d01fd3f9a269a617efd4beea9b8b             = conv_qin_00158_00000;
assign conv_Sgntin_row_00158_00001 = Ie536879e6fa9be65376d7f00e0fc40d0;
assign I106deaff50b8480eac31ddbae2ec7c61             = conv_qin_00158_00001;
assign conv_Sgntin_row_00158_00002 = I3ade5535a79ce83857481ac771cd8618;
assign I5669856f88f5e2c98f64df696db76414             = conv_qin_00158_00002;
assign conv_Sgntin_row_00158_00003 = I9ce3942aba354c1fd7d6b9a39c994d7b;
assign Ib3fb10da528d450251764a9b9ede0dba             = conv_qin_00158_00003;
assign conv_Sgntin_row_00159_00000 = I40a223380fb4414a3f26a08cb90025ec;
assign I9747a02384abb1c2dd1f52b3a5a999cc             = conv_qin_00159_00000;
assign conv_Sgntin_row_00159_00001 = Id0b1c46fa4caa63a4c63a44ba3c5ef8a;
assign I2795d21d343b83a69146314a2407cfa2             = conv_qin_00159_00001;
assign conv_Sgntin_row_00159_00002 = I88a89b2d938552458dab9bc34728959b;
assign I1b7a401bc11741e6f011fb9895b5c797             = conv_qin_00159_00002;
assign conv_Sgntin_row_00159_00003 = I2c6c6041c9c69c84f4d64af6458955f5;
assign Icdc9e676957b2223d60c413331fa982f             = conv_qin_00159_00003;
assign conv_Sgntin_row_00160_00000 = I0c616f736879c28a5222de3d6f49a587;
assign Ib196f5bcf9152703dc32c5101076600a             = conv_qin_00160_00000;
assign conv_Sgntin_row_00160_00001 = I44f170d02bae7fe044456e125a98451d;
assign I165653ab165cfafe2b74cd441331f9e1             = conv_qin_00160_00001;
assign conv_Sgntin_row_00160_00002 = Iefbdf686d9452a62cb99cf023a4d9fe7;
assign I340c98b886123c541a1b8d9fc8a6d48c             = conv_qin_00160_00002;
assign conv_Sgntin_row_00160_00003 = I830a4fffe1244e071eb82c28ddc4a308;
assign I381f6051282c062ccf53866830344cd4             = conv_qin_00160_00003;
assign conv_Sgntin_row_00161_00000 = I620b8ecdcaccc1ec80ebcf9fa6af0017;
assign I9fe11f6c8147391aa4a5afd1a4e4f731             = conv_qin_00161_00000;
assign conv_Sgntin_row_00161_00001 = I94460b6ce7b776bcc5eca149eab80c26;
assign Ibf80bb564263ea85bd886a8617f09bb2             = conv_qin_00161_00001;
assign conv_Sgntin_row_00161_00002 = Ic3ba4531855366e9a060cec1c7694844;
assign I72b1bb104bf2843f161448baf7aab44b             = conv_qin_00161_00002;
assign conv_Sgntin_row_00161_00003 = Ifad8e46fc3844bbfaf434a14f6b5869d;
assign Icfc21935c007fbbceb2a67ebe1a68a0b             = conv_qin_00161_00003;
assign conv_Sgntin_row_00162_00000 = Iec91b3ca3b54010755d57f8b8ea4a544;
assign I8922487573e02d684a3d71448c3828f5             = conv_qin_00162_00000;
assign conv_Sgntin_row_00162_00001 = Idc6b6357741c9887a9db1037ccc2d922;
assign I68bb1f26f878862f288c1f57049cf58b             = conv_qin_00162_00001;
assign conv_Sgntin_row_00162_00002 = I21e72a7e5870151c3247d15121e5fb4f;
assign I848ed394bd4f0b199d11c0ff458394a7             = conv_qin_00162_00002;
assign conv_Sgntin_row_00162_00003 = I10a6c6a8fdb0003de1f360c148777d0f;
assign I120d597a80158374726e064fb0f099fb             = conv_qin_00162_00003;
assign conv_Sgntin_row_00163_00000 = Id806a2df1c4519bbbe811791cb4072f9;
assign I1c85c8f73ef80a6808c6aec0c8eca8ab             = conv_qin_00163_00000;
assign conv_Sgntin_row_00163_00001 = I472352e7027b9df2fa957d9fd68443ff;
assign I50383e3d7c172eedfa00aa50a9faac4c             = conv_qin_00163_00001;
assign conv_Sgntin_row_00163_00002 = I74cbc0ec3bb682e0f927890eef8d7a58;
assign I4c971e714427664c59c6371e14781bae             = conv_qin_00163_00002;
assign conv_Sgntin_row_00163_00003 = I4cde586fc28f8d03fc9934d56f7ff7b8;
assign I2520aa556aadf851f58f0b1820498730             = conv_qin_00163_00003;
assign conv_Sgntin_row_00164_00000 = Ibd59d0e5a062f149bd0e91ba76985a13;
assign I524e78ae6a4204e17ba4532dba047d4b             = conv_qin_00164_00000;
assign conv_Sgntin_row_00164_00001 = I51e14ece9ab6607f83e6ba27f3f046a9;
assign Id1fbbe0594dae272856566522633bb3d             = conv_qin_00164_00001;
assign conv_Sgntin_row_00164_00002 = I433dd5092cf1851cd196feade3cfa6d8;
assign I432aa7cb844286c442356954f8814260             = conv_qin_00164_00002;
assign conv_Sgntin_row_00164_00003 = Ib83a067fb08e118dcf794902beef9405;
assign I6203f49a08107f7185ebadeecf2c16b0             = conv_qin_00164_00003;
assign conv_Sgntin_row_00165_00000 = Ic4c6f707f461cebbc4c93f2ba664ae7b;
assign I4e8ebc46bc068c3f9889d970db131112             = conv_qin_00165_00000;
assign conv_Sgntin_row_00165_00001 = Icc67656ad2dd3fffae4e5abe02f8fff9;
assign Ie1817cbf3a80dae435a5571dfbd2f5ad             = conv_qin_00165_00001;
assign conv_Sgntin_row_00165_00002 = Ib6124faff821158c6a2c9a9c454ab68c;
assign I92678f5b52c9c55556ff7f17f0f607b7             = conv_qin_00165_00002;
assign conv_Sgntin_row_00165_00003 = I358cf9609272a4562423a85f9b2f56bf;
assign Ia706fb593b63cebbee0321c154cb859b             = conv_qin_00165_00003;
assign conv_Sgntin_row_00166_00000 = Ic04828ba2db8239b093043c27476d345;
assign Ib75747cb32130d44b338ed8c8af8ca11             = conv_qin_00166_00000;
assign conv_Sgntin_row_00166_00001 = I38352b363fa37f6f822fbc1a39100968;
assign I43493f70f0336453d77caf7f27503daa             = conv_qin_00166_00001;
assign conv_Sgntin_row_00166_00002 = I759409e242eaeb144a53e630a8cfd514;
assign I7fb3b66cb48521f8715f66bf5642cdb2             = conv_qin_00166_00002;
assign conv_Sgntin_row_00166_00003 = Ic1e9d9113150ad57954c0e369259dc62;
assign Ia4b5f2b07556629673fc6576bc49a5dc             = conv_qin_00166_00003;
assign conv_Sgntin_row_00167_00000 = Ibe6b8c57d7ff47b6fdad5fadf1f6b841;
assign Id1659ccdeaea3e59eb2d3f65a65ebd05             = conv_qin_00167_00000;
assign conv_Sgntin_row_00167_00001 = Ic9b72b2a91d951cf08cf54ed215ecaa8;
assign I9ec9f389d0489908d497487e44c6edcd             = conv_qin_00167_00001;
assign conv_Sgntin_row_00167_00002 = Ied19cb51636bfb029ba8a2c390f97105;
assign I6714551e8885ef5e4490673fe1b2dad1             = conv_qin_00167_00002;
assign conv_Sgntin_row_00167_00003 = If7fe3f5ccbb5b279e41fd183c8ff3974;
assign Ic532c6b85b156f821e0742f47239a65c             = conv_qin_00167_00003;

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
          start_d2 <= 1'b0;
          start_d3 <= 1'b0;
          //start_d4 <= 1'b0;
          //start_d5 <= 1'b0;
          start_d6 <= 1'b0;
          start_d7 <= 1'b0;
          start_d8 <= 1'b0;
          start_d9 <= 1'b0;
       end else begin
          start_d2 <= start_dec | iter_start_int;//start_d1;
          start_d3 <= start_d2;
          //start_d4 <= start_d3;
          //start_d5 <= start_d4;
          start_d6 <= start_d5;
          start_d7 <= start_d6;
          start_d8 <= start_d7;
          start_d9 <= start_d8 ;
       end
   end


assign flogtanh_00000_00000 = ~I5f68368511b59d2e365cc91b806b334e+ 1;
assign flogtanh_00000_00001 = ~I71e4d98dca37256fcc84248a26d703e2+ 1;
assign flogtanh_00000_00002 = ~Ib8380902ac4082f834744ddef6d0cc6a+ 1;
assign flogtanh_00000_00003 = ~I9570f8498d95bee230bb3c5e720bb857+ 1;
assign flogtanh_00000_00004 = ~I55c425102db0a6838012a165c0597680+ 1;
assign flogtanh_00000_00005 = ~Ic970a88c435a85d21ed71c6060b8a8e4+ 1;
assign flogtanh_00000_00006 = ~Iec8dc328edd6cbaa2d697e05ed222746+ 1;
assign flogtanh_00000_00007 = ~I16d2084ccfb102c3bafc701872f5ef2d+ 1;
assign flogtanh_00000_00008 = ~Id680a9affed622577164b3a8380494f5+ 1;
assign flogtanh_00000_00009 = ~Ifcd68be4bea38622d2d57d3a4e6fc5bb+ 1;
assign flogtanh_00000_00010 = ~I16deb9107193a3536979e4b5e5654b9c+ 1;
assign flogtanh_00000_00011 = ~I28cac65a4db3f708cc90a1b023bfe894+ 1;
assign flogtanh_00000_00012 = ~Ie763738b7faf253837e1c45de255cb5e+ 1;
assign flogtanh_00000_00013 = ~Icfef12499b53cd84f0aae067f30c17d0+ 1;
assign flogtanh_00000_00014 = ~I0982b8d7f99aceb8871c9c10448f54c5+ 1;
assign flogtanh_00000_00015 = ~I6c661048307c23c699d4b3636564de0f+ 1;
assign flogtanh_00000_00016 = ~I786dfcaa131b99c254aaff15bd2c2b6d+ 1;
assign flogtanh_00000_00017 = ~I2b49d74cb130542f2ca99534e2c513b1+ 1;
assign flogtanh_00000_00018 = ~I0f6cb7a5a31d6f2f6178632c0c898bc6+ 1;
assign flogtanh_00000_00019 = ~I03bea609a189246a2375b355df47cf81+ 1;
assign flogtanh_00000_00020 = ~If56555b7cf539750706cf678030ccdb2+ 1;
assign flogtanh_00000_00021 = ~I94e89b3a841f9760e3967c97e86d7160+ 1;
assign flogtanh_00001_00000 = ~I8cab6f6faf0758f26d1a8851fae43896+ 1;
assign flogtanh_00001_00001 = ~I6ecf7249e6151477fe74a79d0b126b21+ 1;
assign flogtanh_00001_00002 = ~I3753b2c4ba8f1bee70def390a96586b0+ 1;
assign flogtanh_00001_00003 = ~I9b919f3d4ee3f33506b87bcdaf2d43a3+ 1;
assign flogtanh_00001_00004 = ~Ib3be128b6704cc04c61e0fc9814dcf20+ 1;
assign flogtanh_00001_00005 = ~If365a3c3ef86dca7c7315b91298c2db8+ 1;
assign flogtanh_00001_00006 = ~I83560e8d0f8cd37815cca6336fb2208d+ 1;
assign flogtanh_00001_00007 = ~I099441ae3d3dffe49b18bc578af54dc7+ 1;
assign flogtanh_00001_00008 = ~I58f89947eead94b5054a0fea3520ae33+ 1;
assign flogtanh_00001_00009 = ~Ibf565bf1803ed43120fa54b80f6f1f29+ 1;
assign flogtanh_00001_00010 = ~I619957528c630e7f64924a25127c93fb+ 1;
assign flogtanh_00001_00011 = ~If3cc31fd16469339470702045fc6d0da+ 1;
assign flogtanh_00001_00012 = ~I338ccc17dc6158aec0129c8b0c02c429+ 1;
assign flogtanh_00001_00013 = ~I83d71a89f35eb73265ee3e54184e1277+ 1;
assign flogtanh_00001_00014 = ~I7362f08ed4e4ae309dfbfda112c56ad6+ 1;
assign flogtanh_00001_00015 = ~I8be4be8471625db0749e6385f87d2dcc+ 1;
assign flogtanh_00001_00016 = ~I3d6a685a1913bd8be01fddbce1edec2e+ 1;
assign flogtanh_00001_00017 = ~Ifd77e040c5f82790b1d5636a42fca602+ 1;
assign flogtanh_00001_00018 = ~Ifbe479e5cab3cba43444bec1e12e72a0+ 1;
assign flogtanh_00001_00019 = ~Ia784f35a5a46837b69eb048dabf84052+ 1;
assign flogtanh_00001_00020 = ~I8d0f440df332ea96e2d56eec490fbd51+ 1;
assign flogtanh_00001_00021 = ~I8d431a0524241fa54cf6dd1e79de4c74+ 1;
assign flogtanh_00002_00000 = ~If49f97cc0c42b23ce393b534015559a0+ 1;
assign flogtanh_00002_00001 = ~Ie932a22a7f1fa37087cbc9e8d73efef4+ 1;
assign flogtanh_00002_00002 = ~I2956687a5fc2fba7149889624ef85647+ 1;
assign flogtanh_00002_00003 = ~Iebf28886bd39c2540c90e808a9c20d3d+ 1;
assign flogtanh_00002_00004 = ~I8d4f3e64c8e3b0710a4a6b30d27c8be8+ 1;
assign flogtanh_00002_00005 = ~I16e3f3a6802fd206654bb622fa1393fe+ 1;
assign flogtanh_00002_00006 = ~I4b5713aee09999592256c407d4b8a95a+ 1;
assign flogtanh_00002_00007 = ~Ieb1dbb98d5e5bda5b9ce803857f2ca26+ 1;
assign flogtanh_00002_00008 = ~Ife1c8d014675240a94f1133a78703ed5+ 1;
assign flogtanh_00002_00009 = ~I94d9412a7b43fa0bd4b9a6d32d313fc7+ 1;
assign flogtanh_00002_00010 = ~If13e359e530823319046ce20027445dd+ 1;
assign flogtanh_00002_00011 = ~I221777352b48c4e228c6637410113854+ 1;
assign flogtanh_00002_00012 = ~I1ee46fec2b82cf8e5142f8e2ac5d9d8a+ 1;
assign flogtanh_00002_00013 = ~Ie45aaf966aa0a94803050b5f43d69e6c+ 1;
assign flogtanh_00002_00014 = ~I88aedd7f52399f5fd435c3415f2218ca+ 1;
assign flogtanh_00002_00015 = ~I7651176b0a74846108fbaabc5cc4900a+ 1;
assign flogtanh_00002_00016 = ~I57ac487adc18165136e9b3c7c50f95ad+ 1;
assign flogtanh_00002_00017 = ~Ic95668328a2121027436f682bac50b9c+ 1;
assign flogtanh_00002_00018 = ~I118726375ca9381e45f001965fcefc5b+ 1;
assign flogtanh_00002_00019 = ~Ic8d47ff5d6c31601a57df868da78c2d4+ 1;
assign flogtanh_00002_00020 = ~I7cdc5ada6fc68ee31fd4062e2ff004d3+ 1;
assign flogtanh_00002_00021 = ~I59547aacdcfde31dc016ec2acbb2f4b4+ 1;
assign flogtanh_00003_00000 = ~Ia7f53f0cd86055da72c13ac474f052a1+ 1;
assign flogtanh_00003_00001 = ~I915054f2fbb8b93516d8748a3e3e29e2+ 1;
assign flogtanh_00003_00002 = ~If257757fa31c2f4cc9ec322e4ecccf83+ 1;
assign flogtanh_00003_00003 = ~If91268e2b84df18785cd6a53e53eb4e9+ 1;
assign flogtanh_00003_00004 = ~Ia072f1d679429d3c3180f8eb67fc7dd7+ 1;
assign flogtanh_00003_00005 = ~I91a8168d3b087ab3891cd6d479427b95+ 1;
assign flogtanh_00003_00006 = ~Id1dce8c1542f1279badb381aca3c9b51+ 1;
assign flogtanh_00003_00007 = ~I8983f003c30a218543f39f5bbcd9a25c+ 1;
assign flogtanh_00003_00008 = ~Id1b5c33bc63f75561b7cce6fc0981c69+ 1;
assign flogtanh_00003_00009 = ~I003f95fb8f2027efa41a1936e8b53986+ 1;
assign flogtanh_00003_00010 = ~Ie16dc913f571ae73ce03d755077345a9+ 1;
assign flogtanh_00003_00011 = ~I86e53eed5b857c439039238bb486067c+ 1;
assign flogtanh_00003_00012 = ~I89433799cfa534afd66e8d6b9f1b62b9+ 1;
assign flogtanh_00003_00013 = ~I80f2e8f6743e28e86e4d85b295e2f768+ 1;
assign flogtanh_00003_00014 = ~I1391018fb93372ccc2fcc08700e38b65+ 1;
assign flogtanh_00003_00015 = ~I8fd26d47ecd4cdd08294cf6133468d17+ 1;
assign flogtanh_00003_00016 = ~I7097c9518bb3351818b96f31ed49c6d3+ 1;
assign flogtanh_00003_00017 = ~Id683d693cd50645c3d6d657aa1c8bdb2+ 1;
assign flogtanh_00003_00018 = ~I88bd8012c93dd9e2ed52ea5e9b8b0004+ 1;
assign flogtanh_00003_00019 = ~Ia8d3667adc34b2b50acf7edb970538d8+ 1;
assign flogtanh_00003_00020 = ~I3f0bba472e912f11dea8e788fbc1cb63+ 1;
assign flogtanh_00003_00021 = ~I6dc671e73b4e9c70cabfdeaac2e5c40b+ 1;
assign flogtanh_00004_00000 = ~Ia6255a136d5f36ea6cba654bd5823850+ 1;
assign flogtanh_00004_00001 = ~I2b9584392ef9a7828ff57bd4c522a302+ 1;
assign flogtanh_00004_00002 = ~I6c1235e88ae444a96ea64fd1bfd04d8f+ 1;
assign flogtanh_00004_00003 = ~Id09b8242c22851fb960d55222fe733d4+ 1;
assign flogtanh_00004_00004 = ~Ie355fa27abbc41291eaf08f2cf9a6ff7+ 1;
assign flogtanh_00004_00005 = ~I566224393f6bb27bfd8b0b0d6b8e53d6+ 1;
assign flogtanh_00004_00006 = ~I8fcad6e7d5ffc9f79eaaf634f6fe8cda+ 1;
assign flogtanh_00004_00007 = ~I6f0f74dcc830fdcb0af9df75a2b722f7+ 1;
assign flogtanh_00004_00008 = ~Idd95fd099dd2b53c46d02f09575b8032+ 1;
assign flogtanh_00004_00009 = ~I0f277bc88d46a4e6e9f1f2c410b503fd+ 1;
assign flogtanh_00004_00010 = ~I66b92f1de2cf408c3af53b161a6ffa60+ 1;
assign flogtanh_00004_00011 = ~Id28d9545e8d20ac080fbac5e345692da+ 1;
assign flogtanh_00004_00012 = ~I4a5cfd6ebd47cda4fa2e06ba9ad6e5b2+ 1;
assign flogtanh_00004_00013 = ~I62bda8dc70e0b5eb38abe094bbe92fc6+ 1;
assign flogtanh_00004_00014 = ~I223b05d94c09b095d1988df121aa5e37+ 1;
assign flogtanh_00004_00015 = ~I5f73e5faf1aca83ee0a415c9ac4a1b9a+ 1;
assign flogtanh_00004_00016 = ~I75f9d3a41019dca3044a1c2cf7069662+ 1;
assign flogtanh_00004_00017 = ~I820fa56328e3919970dd64adb1d4d8e7+ 1;
assign flogtanh_00004_00018 = ~I05eadf11cdc6c2f2b021e33f2438fa49+ 1;
assign flogtanh_00004_00019 = ~I2c487770d606451440eecf358202db32+ 1;
assign flogtanh_00004_00020 = ~I082aa8c413d7ef8f054b1c2857cbe39f+ 1;
assign flogtanh_00004_00021 = ~I420e2c5a8745133f6263a71b458f1e2f+ 1;
assign flogtanh_00004_00022 = ~I4b8d520ee88fd39d83a16432e962f731+ 1;
assign flogtanh_00005_00000 = ~Ia3f7f07ddb09ea33218afe14281ac3c6+ 1;
assign flogtanh_00005_00001 = ~I25aefb53f59a00abe88b9dcf6be6907a+ 1;
assign flogtanh_00005_00002 = ~I22c3140a8db02352d2e2a2a11eeba117+ 1;
assign flogtanh_00005_00003 = ~I954dd66f60316803a8f13a39c460a39a+ 1;
assign flogtanh_00005_00004 = ~I37b3988d699a1ed42923e3fd1584ecc0+ 1;
assign flogtanh_00005_00005 = ~If79bc5a35cb55036a367efb88c7d5510+ 1;
assign flogtanh_00005_00006 = ~Ideab06dc2448a6950cd1a06a0c90c2c6+ 1;
assign flogtanh_00005_00007 = ~I1d7d7a68fc53b8be89c4637ac8f29380+ 1;
assign flogtanh_00005_00008 = ~Ib34ad1d14978608d1440f59998a31672+ 1;
assign flogtanh_00005_00009 = ~Id081512cd113e4d09df0fb13e443d76b+ 1;
assign flogtanh_00005_00010 = ~I57a0f8c3710cf8e216d6dc2420f7621c+ 1;
assign flogtanh_00005_00011 = ~Iaa164a078c8cdaad694a053c9c1e0313+ 1;
assign flogtanh_00005_00012 = ~I7eb76b3d17296fdae702d8f820f1428d+ 1;
assign flogtanh_00005_00013 = ~I00ecb5e329390023b318a2ceba0df231+ 1;
assign flogtanh_00005_00014 = ~Iea32ebc385c6cfc9212ff37973a0a05d+ 1;
assign flogtanh_00005_00015 = ~If845af0d620024f04525244753ba5d18+ 1;
assign flogtanh_00005_00016 = ~I08e907b0619bec3ef2cf4cb3779e0794+ 1;
assign flogtanh_00005_00017 = ~I68e5b12792a86dda0576742831d3b728+ 1;
assign flogtanh_00005_00018 = ~I72db05084d30d7c59ba1cb06d3b09400+ 1;
assign flogtanh_00005_00019 = ~Ib1f1aef6c0a9291553b62fd555feb2e7+ 1;
assign flogtanh_00005_00020 = ~Ib504b808f724ca6032e7c746517cd4fd+ 1;
assign flogtanh_00005_00021 = ~Ia47f7fb27f2d965cfd2989569c257356+ 1;
assign flogtanh_00005_00022 = ~If2b17f9e9186542117f43d0dd342326e+ 1;
assign flogtanh_00006_00000 = ~I6c4ba0863ab4c8d1a56324a4d89ccbeb+ 1;
assign flogtanh_00006_00001 = ~I4dbd1bb8f1641f15e3a4f1e309962811+ 1;
assign flogtanh_00006_00002 = ~I26781ef851ed43c6f88ff1215cddca6b+ 1;
assign flogtanh_00006_00003 = ~Ia349e1f7c10a63ddccb3f300c73b4572+ 1;
assign flogtanh_00006_00004 = ~I50c4e1d3a3f63b93bc36b5141226fb3c+ 1;
assign flogtanh_00006_00005 = ~I12334038c2be8634c47869f397503019+ 1;
assign flogtanh_00006_00006 = ~I64692d5168554dfd7ce1c7a046aecf72+ 1;
assign flogtanh_00006_00007 = ~Ia4b438844530fff602ea04e72b07db8d+ 1;
assign flogtanh_00006_00008 = ~I9574759e112f27778f3645d5d49126b7+ 1;
assign flogtanh_00006_00009 = ~I2ffb7c2ad09bac694ef13ec41e5de327+ 1;
assign flogtanh_00006_00010 = ~Ib190f589f4d663dbc0a3c166a8dcf5fa+ 1;
assign flogtanh_00006_00011 = ~I459c59ac61179d74170db53bf45ba89e+ 1;
assign flogtanh_00006_00012 = ~Ie5e432a991aff25577639f1b4ffd594f+ 1;
assign flogtanh_00006_00013 = ~I72064a6a84ff956d76a5aa590bbc05a9+ 1;
assign flogtanh_00006_00014 = ~Iea74ecbac92e1b8f2ec7ad68d10b8e7d+ 1;
assign flogtanh_00006_00015 = ~I4f72d0db9fcc358c6fbec9964fbe0bbb+ 1;
assign flogtanh_00006_00016 = ~Ifd958901d2ea2284f506e04a058012fa+ 1;
assign flogtanh_00006_00017 = ~Ie317bbd70b9092b840c0f2713204fb9d+ 1;
assign flogtanh_00006_00018 = ~I2f9e56d570e72714a06c59aa9e4334c0+ 1;
assign flogtanh_00006_00019 = ~I5b53fd45210b92703cb10d583f471ab9+ 1;
assign flogtanh_00006_00020 = ~I8edbe77bacf1975e014faeee6b861980+ 1;
assign flogtanh_00006_00021 = ~I174fcbc2ee01fc55edbc8238e5da7f0c+ 1;
assign flogtanh_00006_00022 = ~Id4dc304aef5f35f6ceb91796c278e716+ 1;
assign flogtanh_00007_00000 = ~I0cbdfae6f75a639eb591d9c0022f5838+ 1;
assign flogtanh_00007_00001 = ~I088898ee932a96c14f2f0f568f5455b6+ 1;
assign flogtanh_00007_00002 = ~Ide0abde3644a4fafb436aa59768d016e+ 1;
assign flogtanh_00007_00003 = ~I08581dc8d42be712cfb36d744f2786e0+ 1;
assign flogtanh_00007_00004 = ~I29fb3830a5fc5922f1ec687a38941e97+ 1;
assign flogtanh_00007_00005 = ~I715d59fb27e519a9b76bdd8b5139a619+ 1;
assign flogtanh_00007_00006 = ~Ibe6a876a041198a581c95457a7d1fcf8+ 1;
assign flogtanh_00007_00007 = ~Iec078a95a69b081cfb5e987ba9c5a613+ 1;
assign flogtanh_00007_00008 = ~I0e8f3f56bce3be1ee4d5f780a2f2a9fe+ 1;
assign flogtanh_00007_00009 = ~Ia73cacadbf80c0701a5b5b430c0d5c98+ 1;
assign flogtanh_00007_00010 = ~Ic634d26fc09589a29a160e4efb5613a8+ 1;
assign flogtanh_00007_00011 = ~Ie1374cac341cf353b1863dae9f544e8b+ 1;
assign flogtanh_00007_00012 = ~Ia07447985347e9a7f3739bd98867cdfb+ 1;
assign flogtanh_00007_00013 = ~I2121318f589878b4a9260625f97de518+ 1;
assign flogtanh_00007_00014 = ~Ibd8424c228f87f85df3da6204edff2b5+ 1;
assign flogtanh_00007_00015 = ~I8a7fb51566bf215af214cd2fb5209974+ 1;
assign flogtanh_00007_00016 = ~I7c0f872988488ac69815d288885dfd2f+ 1;
assign flogtanh_00007_00017 = ~I3521b10b97b0e74888ce385cfc772945+ 1;
assign flogtanh_00007_00018 = ~I58f0b81a46549cab8e74ecbc285df23a+ 1;
assign flogtanh_00007_00019 = ~I7095040b38bf9d6b5229c11d2a0d7c57+ 1;
assign flogtanh_00007_00020 = ~I675ab6c4fb93b006f3fcafc985fbc405+ 1;
assign flogtanh_00007_00021 = ~I239a992ebb62899120a74b1c9e6cc4b4+ 1;
assign flogtanh_00007_00022 = ~I927c870d09285dcb47e6d399f319471e+ 1;
assign flogtanh_00008_00000 = ~Ie23ed3ee61f468f59f2baf661cb7f85d+ 1;
assign flogtanh_00008_00001 = ~I68e58664be09261e5a80d6f8ecdd1b60+ 1;
assign flogtanh_00008_00002 = ~Id2808e0f40992c79ead4da7c734e5b79+ 1;
assign flogtanh_00008_00003 = ~Icb2b390266bff241a688961136db0f51+ 1;
assign flogtanh_00008_00004 = ~I54cfd68212d97a2cc8241ef429429453+ 1;
assign flogtanh_00008_00005 = ~I8d4e3962525c424786ae822a6981a5e6+ 1;
assign flogtanh_00008_00006 = ~I1a5f22b4e326d1684c0a8c7a7e754ab4+ 1;
assign flogtanh_00008_00007 = ~I8c2e0c83a8204d6b21e0e3e458d56f05+ 1;
assign flogtanh_00008_00008 = ~Ie0622ff815747e4a9f368c74787026ec+ 1;
assign flogtanh_00008_00009 = ~I5ffed139764d90825b9f2eddacd0eddc+ 1;
assign flogtanh_00009_00000 = ~I5a3297f48e1045273db6522744582b05+ 1;
assign flogtanh_00009_00001 = ~I9858bb2a3cc458aca5bf7eb077ee55dd+ 1;
assign flogtanh_00009_00002 = ~I6e7e27bb176196e4493bf9c45ca19719+ 1;
assign flogtanh_00009_00003 = ~I4cff1804df738cbf4f940c775236df9c+ 1;
assign flogtanh_00009_00004 = ~I0c1e22375d5e023c24519901b92eceb5+ 1;
assign flogtanh_00009_00005 = ~Ida5b16851dc06534844a0b037d74feb3+ 1;
assign flogtanh_00009_00006 = ~Iac3cb5b4481687fcf430c8bf52cfb74d+ 1;
assign flogtanh_00009_00007 = ~Ia1499972c4995268acd828c1289f353d+ 1;
assign flogtanh_00009_00008 = ~Ie559401a3a913400dc5e3e5641297fa6+ 1;
assign flogtanh_00009_00009 = ~Ie0667fbe76244eaec0b155d69dcc9447+ 1;
assign flogtanh_00010_00000 = ~I1d0f031e8ae9c0335d501d1565118220+ 1;
assign flogtanh_00010_00001 = ~Ie2c801b2de066c3218d7312615b7bfda+ 1;
assign flogtanh_00010_00002 = ~I64c4bb0d40d80ec52aab61ce46954f43+ 1;
assign flogtanh_00010_00003 = ~I512f57a40c7c8cb2f040bdde73e44ca3+ 1;
assign flogtanh_00010_00004 = ~Id60cbf534604e5dba988050ef5abe625+ 1;
assign flogtanh_00010_00005 = ~I37998a91d20db2248ebdd8e661d42f70+ 1;
assign flogtanh_00010_00006 = ~Ib65ff82aff398f6ff7ba711a36f41ee4+ 1;
assign flogtanh_00010_00007 = ~I3d1dd8b9c7c6d3913f7ac369ad7e625c+ 1;
assign flogtanh_00010_00008 = ~I097722547450582dc5776bdaff914741+ 1;
assign flogtanh_00010_00009 = ~Id4a213e494f9c9be0fd1a307e87c756a+ 1;
assign flogtanh_00011_00000 = ~I21594c8b0169efd7c2aa6cbc31f4a901+ 1;
assign flogtanh_00011_00001 = ~I15022e1b349eee259d3567837283dbf6+ 1;
assign flogtanh_00011_00002 = ~I1070940dc2ef6e8ee3d1227ec9ff3162+ 1;
assign flogtanh_00011_00003 = ~I8922cc37cde6ba132f632743113e42af+ 1;
assign flogtanh_00011_00004 = ~Ia66c399023e500ed67197dcf236f5d42+ 1;
assign flogtanh_00011_00005 = ~I1171dc208d5db1024dc3f09a90c78ca0+ 1;
assign flogtanh_00011_00006 = ~Ic28b148967a5b3d05409976fa9001ac8+ 1;
assign flogtanh_00011_00007 = ~I79fe46308b93fbb24245fe1c75edf4a5+ 1;
assign flogtanh_00011_00008 = ~I3bfcd63e92f1949234ab1d2701dbb499+ 1;
assign flogtanh_00011_00009 = ~I5e2331edf6e881e9f3a8c47eebda0ac4+ 1;
assign flogtanh_00012_00000 = ~I4b66c202450986ef0df05e979cc8bc7f+ 1;
assign flogtanh_00012_00001 = ~I737daf208eccf95feb3192897586cdce+ 1;
assign flogtanh_00012_00002 = ~I29c8133231cfda17668bbe7b692bdfe2+ 1;
assign flogtanh_00012_00003 = ~Id9d56f09595e80d66c2ac300f7d1d972+ 1;
assign flogtanh_00012_00004 = ~I97e89a2ee18d2688d7c1a640318a1e0d+ 1;
assign flogtanh_00013_00000 = ~Ife123bf57fe693dabe6aeaa236c4e058+ 1;
assign flogtanh_00013_00001 = ~I0c0d844fe3b7d35c1ed6bd7cc4e0dc24+ 1;
assign flogtanh_00013_00002 = ~I2d9632ae6a0f3ba44c3da8f56ba3fedf+ 1;
assign flogtanh_00013_00003 = ~I38cc7b117c0bcd5e3060cd370d710d7e+ 1;
assign flogtanh_00013_00004 = ~I793ddbf6a5d026a57ab72984ca19deac+ 1;
assign flogtanh_00014_00000 = ~I79458089b042e181e37cc44c06d08681+ 1;
assign flogtanh_00014_00001 = ~I42460fae0acff25fa2b829e39ddcc4fd+ 1;
assign flogtanh_00014_00002 = ~Id3670a6f05d40ab69624544de92b9c64+ 1;
assign flogtanh_00014_00003 = ~I81800fb49855a4fd2737faa07ff15d29+ 1;
assign flogtanh_00014_00004 = ~Ibfe325e48511372569e0d98d9c4e70e3+ 1;
assign flogtanh_00015_00000 = ~I326660e98f61bb2ced4c23c7bcc9324a+ 1;
assign flogtanh_00015_00001 = ~Ic6fa98631d742b27f252fe7c95caef55+ 1;
assign flogtanh_00015_00002 = ~Iab6d0f72579687407e029c630b107f7d+ 1;
assign flogtanh_00015_00003 = ~I19eae741ef89baa1a64c403fb29f14f4+ 1;
assign flogtanh_00015_00004 = ~I749b9c345f23aae03c595a2c76126ecb+ 1;
assign flogtanh_00016_00000 = ~Idc77c7d5123717fc2596a51d904c6d82+ 1;
assign flogtanh_00016_00001 = ~I779da979707d9712c1626d6025f97599+ 1;
assign flogtanh_00016_00002 = ~I97aede8502e443f98938487a5a5c072c+ 1;
assign flogtanh_00016_00003 = ~Ie7820d1a242bc28c19ec32d2c91e47b7+ 1;
assign flogtanh_00016_00004 = ~I82a14e1ee4723e7d9a13c1f2b8b13691+ 1;
assign flogtanh_00017_00000 = ~I77a94cd9186ca546ca9664942ea3537f+ 1;
assign flogtanh_00017_00001 = ~I3c0ddec25c53c166d30eb78d4518840e+ 1;
assign flogtanh_00017_00002 = ~I98bbe3b75958f10195dee6460cf2aca6+ 1;
assign flogtanh_00017_00003 = ~If6d436031f68ef587750c5c1dfcfffc2+ 1;
assign flogtanh_00017_00004 = ~I461398638cb8280f1779915298540b00+ 1;
assign flogtanh_00018_00000 = ~I20c65000bbc10299168af7390776a03c+ 1;
assign flogtanh_00018_00001 = ~Ia840e19ca36795a50ab1a6e6a1729edb+ 1;
assign flogtanh_00018_00002 = ~I7d98d1e5f07fccff5f20eaca6363c700+ 1;
assign flogtanh_00018_00003 = ~I97a75b8625ae2a143cf364790ae77753+ 1;
assign flogtanh_00018_00004 = ~Idbea892c8109117f90b453efe8ae25af+ 1;
assign flogtanh_00019_00000 = ~Icfc1c6d96a3598af73e99a350c387d72+ 1;
assign flogtanh_00019_00001 = ~I523e9b6f828ec7f166750112f8a3f676+ 1;
assign flogtanh_00019_00002 = ~I79259217f63b2f6263552c434d0e5c93+ 1;
assign flogtanh_00019_00003 = ~Ice6db5ba70d3c7499df6723a2df56bfe+ 1;
assign flogtanh_00019_00004 = ~I28aa517220bf597cf898660f698ef19d+ 1;
assign flogtanh_00020_00000 = ~I07048dc5cbe24ff72d24902d572face0+ 1;
assign flogtanh_00020_00001 = ~Iab3876e5107e3a56b1fafe41e16d9482+ 1;
assign flogtanh_00020_00002 = ~I511a55c2f4d6d3727dff5825597f55a9+ 1;
assign flogtanh_00020_00003 = ~I2493237a24acdcab8b5bda10e804a5cf+ 1;
assign flogtanh_00020_00004 = ~I03829256e357ac17c7ca7cae2f980f41+ 1;
assign flogtanh_00020_00005 = ~Iae32c44b88fe7ddb5d4f19cf8fff3ba6+ 1;
assign flogtanh_00020_00006 = ~I3bdc5ba374f85dc61346e4868c41a6bf+ 1;
assign flogtanh_00020_00007 = ~I557ef77ce931535467a07a8d70145f55+ 1;
assign flogtanh_00020_00008 = ~Ib4695d4389db72c5ac7e31809072c290+ 1;
assign flogtanh_00020_00009 = ~Ie81315a3a14a5ef879d8e3f405936365+ 1;
assign flogtanh_00020_00010 = ~Ia7520053a7c4a94437c6a780b03a28a5+ 1;
assign flogtanh_00020_00011 = ~Ic308a5413f38b96d244cac3b0bc9462c+ 1;
assign flogtanh_00020_00012 = ~I034fb3850485fae2d1358041a1c41888+ 1;
assign flogtanh_00020_00013 = ~I0e7079db66c15210046b997f319ece89+ 1;
assign flogtanh_00021_00000 = ~I9a5388f8aa6e9924a309aa8db4c1983b+ 1;
assign flogtanh_00021_00001 = ~Ief76663994991118b1899ea4ddf4527d+ 1;
assign flogtanh_00021_00002 = ~I6fb63ea54e492bdbc6d1145affc683e9+ 1;
assign flogtanh_00021_00003 = ~If83ce1cbe3a73472419520c225b288a6+ 1;
assign flogtanh_00021_00004 = ~Id1df78ab32daf524b77c0431c782f2bf+ 1;
assign flogtanh_00021_00005 = ~Iff142b88493149045fc0de355b767c16+ 1;
assign flogtanh_00021_00006 = ~I28c3818247c7c6de11790f6692882b5a+ 1;
assign flogtanh_00021_00007 = ~Ib451127b69a0a800332a712af77c6d29+ 1;
assign flogtanh_00021_00008 = ~I3d601db540da359ae4d22f960d3d5af8+ 1;
assign flogtanh_00021_00009 = ~I2c1f2476efe593829ade470fe8ec2526+ 1;
assign flogtanh_00021_00010 = ~I7e685b06df8a8c2ac351fa9f9b76a81d+ 1;
assign flogtanh_00021_00011 = ~I1338d211b5d2d409bfe0df76d2ca2701+ 1;
assign flogtanh_00021_00012 = ~Ia40dad546d9c852e2fa8942c62a1c1f8+ 1;
assign flogtanh_00021_00013 = ~I0b0dd019d8bd24684403a29aed668b6d+ 1;
assign flogtanh_00022_00000 = ~I66a304016a9adfd85a2abb6f8fd39afc+ 1;
assign flogtanh_00022_00001 = ~I177be24718c59688752097fe2a4085c4+ 1;
assign flogtanh_00022_00002 = ~I7e66a42eb7cdb820cd1297c39f0625e8+ 1;
assign flogtanh_00022_00003 = ~If2021f0735c6c5649ebac0d230fda87c+ 1;
assign flogtanh_00022_00004 = ~Ie1bf5d97b8f679095d2442bbf9f95608+ 1;
assign flogtanh_00022_00005 = ~I632469889d6bb1c268b45fb805467ebd+ 1;
assign flogtanh_00022_00006 = ~Ie230ba3c73808e102eee9e5868595e7c+ 1;
assign flogtanh_00022_00007 = ~Ie1e9326e4eee006ec07abb6bb7d269a5+ 1;
assign flogtanh_00022_00008 = ~Ica4ec1647bdb5a3aad6db6b447bd7995+ 1;
assign flogtanh_00022_00009 = ~Ia17295aec0a40c2b46a595dacfede2d5+ 1;
assign flogtanh_00022_00010 = ~I4c6d3d6fc2d10066a744fdd9405a7902+ 1;
assign flogtanh_00022_00011 = ~Ia9c043c5e8873fd13e39cf6bd8136c51+ 1;
assign flogtanh_00022_00012 = ~I2e802c75c6ce34b05943b678ecbfacb1+ 1;
assign flogtanh_00022_00013 = ~Ieb3f28762410fb40a0c8a8556b4b3ca0+ 1;
assign flogtanh_00023_00000 = ~Ie3e0c0e40c7a67ce7f957e74bd2a895d+ 1;
assign flogtanh_00023_00001 = ~I491f2373b2df19a4c22e1787ef034179+ 1;
assign flogtanh_00023_00002 = ~Ief96603d41b4f670d2bbfa3d3875c903+ 1;
assign flogtanh_00023_00003 = ~I7a029c27d92754041eb6d605837238dd+ 1;
assign flogtanh_00023_00004 = ~I00dad36628d2fa923120fdaa79bf0045+ 1;
assign flogtanh_00023_00005 = ~I3707f68de059df0af5c652fc0478e543+ 1;
assign flogtanh_00023_00006 = ~I94af4b6b9dc11935db54ba872889392d+ 1;
assign flogtanh_00023_00007 = ~I38e2dbba093928b874d447362d89b291+ 1;
assign flogtanh_00023_00008 = ~Ia48f0029e9e76386f3dd70aacd9adbfa+ 1;
assign flogtanh_00023_00009 = ~Ic2b20168744fafbe15037ed7fa83da72+ 1;
assign flogtanh_00023_00010 = ~I62fdc8936121a2707d94cf3bd6e660ac+ 1;
assign flogtanh_00023_00011 = ~Ia0932b3fd6a5ae6da2bacd2b86ba3a43+ 1;
assign flogtanh_00023_00012 = ~I9fce6091885f1bb97d29fb1f543b1a38+ 1;
assign flogtanh_00023_00013 = ~Ib402cdbfaa9900820b85bd625415c547+ 1;
assign flogtanh_00024_00000 = ~I518a2736384c14c02f27bfa3d8ea7aff+ 1;
assign flogtanh_00024_00001 = ~I847cf7ff866f8a666872c12d6b67b1b1+ 1;
assign flogtanh_00024_00002 = ~I9e45e3d7117ce48cdbfc5db8c0ccfcf4+ 1;
assign flogtanh_00024_00003 = ~I380ff8528cdba4026fac3c4eda8b2c52+ 1;
assign flogtanh_00024_00004 = ~Iee8f9b0654f6f6797f11cae0947e454e+ 1;
assign flogtanh_00024_00005 = ~Ie3e54a4700d8d0f6478187e06cb6f85d+ 1;
assign flogtanh_00024_00006 = ~I8c0069e8756bcff203ce21ae3170aa42+ 1;
assign flogtanh_00025_00000 = ~I856eada207c5006beb8f83f01d5d74c9+ 1;
assign flogtanh_00025_00001 = ~I79a46279070c53678a5af54f661c5821+ 1;
assign flogtanh_00025_00002 = ~Ica807adc510a2e32580ca77c18ea0b45+ 1;
assign flogtanh_00025_00003 = ~Ia8094903aed8dd0ce8e9ff459a5287b0+ 1;
assign flogtanh_00025_00004 = ~Ie018f3003c5f124bddd13c359257bf35+ 1;
assign flogtanh_00025_00005 = ~Ice18bceb10fec484ffc96155e14c4974+ 1;
assign flogtanh_00025_00006 = ~Ib484aa64b795f7e36198b800f302164f+ 1;
assign flogtanh_00026_00000 = ~Icdb143a4ce96029c2441758bf2edd7b0+ 1;
assign flogtanh_00026_00001 = ~I3a76f70ca3bfbcacc6f3342aa71f1912+ 1;
assign flogtanh_00026_00002 = ~I9470c7ab9634c01bb832c9e4ff5496bf+ 1;
assign flogtanh_00026_00003 = ~I218ee96418a4f5d734d3d71685bc09c7+ 1;
assign flogtanh_00026_00004 = ~I924514226fdb5bac110a2650bcb2e85f+ 1;
assign flogtanh_00026_00005 = ~Idc57f37015a48393608e2b026bc7065c+ 1;
assign flogtanh_00026_00006 = ~I41af7e4c97fc04154fe6de66b82499f5+ 1;
assign flogtanh_00027_00000 = ~I972bee4216f8e532e8fa4bd25fbb9c57+ 1;
assign flogtanh_00027_00001 = ~Ib303ea0240e7ab5f000dd10e975b2274+ 1;
assign flogtanh_00027_00002 = ~I5971253546899e9a82f387d5eabcc7b3+ 1;
assign flogtanh_00027_00003 = ~I1fc36e6f738fab96df356979e1e3a612+ 1;
assign flogtanh_00027_00004 = ~Ie2d8c84d8c9a4c8f637068a2ae39fdde+ 1;
assign flogtanh_00027_00005 = ~I114c595caa67a3f777f087a634130a6d+ 1;
assign flogtanh_00027_00006 = ~Idad14b6383b9af54eb35e72ff3d10035+ 1;
assign flogtanh_00028_00000 = ~I46e9c76b19ed1ff21f102efe6ee5c732+ 1;
assign flogtanh_00028_00001 = ~Ic75b8bbb1b80001ec188a0cd25623420+ 1;
assign flogtanh_00028_00002 = ~Idc7df6877bdb7e7d392307d78183d31c+ 1;
assign flogtanh_00028_00003 = ~Ib8b95ece5da3877b261a06e6d0571921+ 1;
assign flogtanh_00028_00004 = ~Ic99654bf4833c9132912eeb4c0dc92fa+ 1;
assign flogtanh_00028_00005 = ~I2461055ef9b1aa2ffca0f5cac3300e71+ 1;
assign flogtanh_00028_00006 = ~I2bc3ffbe5b42b0833206437d3863278e+ 1;
assign flogtanh_00028_00007 = ~Id5e02d4c48fa6c3b0d45a9e66f09448f+ 1;
assign flogtanh_00028_00008 = ~I40e99289d5762e77a3766eb8251eef00+ 1;
assign flogtanh_00028_00009 = ~I20beb3fdbe91936f74a200cd8ec9817b+ 1;
assign flogtanh_00028_00010 = ~Id435b68afb53bef4afc7b70a9512e955+ 1;
assign flogtanh_00028_00011 = ~I0cf5cb4cd472502b84dbf6fe1af0be78+ 1;
assign flogtanh_00028_00012 = ~Iacf6340a29a5592b61ea875304a2de48+ 1;
assign flogtanh_00029_00000 = ~I5dfc71255cba279420b7545df4d35c40+ 1;
assign flogtanh_00029_00001 = ~Ibadcb205c7e9a0f3345cac7eb41b5985+ 1;
assign flogtanh_00029_00002 = ~I762b2abb876381eff6de97cef0798405+ 1;
assign flogtanh_00029_00003 = ~Ib3e7633767b6e09e4ee54f6feaddd31e+ 1;
assign flogtanh_00029_00004 = ~I3f193e9c265c1dfaeada63d59db5b79f+ 1;
assign flogtanh_00029_00005 = ~Ie72268e979cf069b88f6eadde789e5ab+ 1;
assign flogtanh_00029_00006 = ~I5732fdb805258fc13c8ba4aaf56574ca+ 1;
assign flogtanh_00029_00007 = ~I3afe987d8f2c93cc19534a3221d1939c+ 1;
assign flogtanh_00029_00008 = ~Ic66af6c3c0268cfb0e9f0776c4f4e961+ 1;
assign flogtanh_00029_00009 = ~Ia605d14205926b3edc6d1c2f69f70ac0+ 1;
assign flogtanh_00029_00010 = ~I0071f2168787bd42ab7f2370aed9d0f5+ 1;
assign flogtanh_00029_00011 = ~I4936f823841b0ffe32f801f5134c0211+ 1;
assign flogtanh_00029_00012 = ~I5975ef8f6cf53cf2132cdd9d707e7912+ 1;
assign flogtanh_00030_00000 = ~I954ff0f9ee871a31774a3d786128fa13+ 1;
assign flogtanh_00030_00001 = ~I31f6bbfbbbd4c20d0c5c71663da1d4c1+ 1;
assign flogtanh_00030_00002 = ~I1898bc3cc6a8b6f71d65c758d1f08366+ 1;
assign flogtanh_00030_00003 = ~If86532f849bd392dbf599eeb2fae0545+ 1;
assign flogtanh_00030_00004 = ~Ia344734d285ac29b53cf401c08a0f987+ 1;
assign flogtanh_00030_00005 = ~I502a8e382aa0881dc86f3c13e0566ca3+ 1;
assign flogtanh_00030_00006 = ~Ic462cebbfc39190b22d20013259e39eb+ 1;
assign flogtanh_00030_00007 = ~I385d03def4cfb49f54867687ebd710ed+ 1;
assign flogtanh_00030_00008 = ~If8aa3ec1b5a4a3c122da82467be917da+ 1;
assign flogtanh_00030_00009 = ~I8daf79a0a2ee1bac7f055af441539fa4+ 1;
assign flogtanh_00030_00010 = ~I6261e0d339762cb2364421e6b87086cb+ 1;
assign flogtanh_00030_00011 = ~I0e2f746715b901feb69f6b3c94f3a828+ 1;
assign flogtanh_00030_00012 = ~I7b8da162c08f8aa2ae90522ee1526cf6+ 1;
assign flogtanh_00031_00000 = ~I5e8ecdbb018402b2fbc0049ee44bae8c+ 1;
assign flogtanh_00031_00001 = ~I06d859184884c07a14c83d2f06587ad5+ 1;
assign flogtanh_00031_00002 = ~I79e3e49f57d47231c0fe6aaafdbc57f1+ 1;
assign flogtanh_00031_00003 = ~I12c07042202f66db926861c9ce7c2b25+ 1;
assign flogtanh_00031_00004 = ~I9d0fdb45b9e86bd409740e538a690320+ 1;
assign flogtanh_00031_00005 = ~Id5fd6f25dc3df22a322434ae3c90dea6+ 1;
assign flogtanh_00031_00006 = ~Id812a8ea2a3b4a912d151be582833fcf+ 1;
assign flogtanh_00031_00007 = ~Ifd3638d44e1ba2285891fac152dee327+ 1;
assign flogtanh_00031_00008 = ~Idd1b6014de2f053554ed09c29bf3e640+ 1;
assign flogtanh_00031_00009 = ~I0d96336eb4d5071d7e1d350e86513b25+ 1;
assign flogtanh_00031_00010 = ~I31e5b2cdc3dc571eafa37510076bcc64+ 1;
assign flogtanh_00031_00011 = ~Ia8849f78971a45ed0daa2489e7d27dd7+ 1;
assign flogtanh_00031_00012 = ~Ie4749f8e9ad2b370f9f9814b5a463c43+ 1;
assign flogtanh_00032_00000 = ~I3096d11098113da669ee0a94686e600d+ 1;
assign flogtanh_00032_00001 = ~I09a1d04c307fcb8a0e30925d86df3fe9+ 1;
assign flogtanh_00032_00002 = ~Idb0a98cea3ee6cd4308bfc2414a003e1+ 1;
assign flogtanh_00032_00003 = ~Id4788855f9a503e8b506d012aaeea445+ 1;
assign flogtanh_00032_00004 = ~I5b937934e7aae1f916c2848889f12685+ 1;
assign flogtanh_00032_00005 = ~I9275bb36e58e0f17964e13ee7f027ab7+ 1;
assign flogtanh_00033_00000 = ~I02330ade2eed926076cc071e45eed82c+ 1;
assign flogtanh_00033_00001 = ~I296bc392d4223cbdd6f77be6523df819+ 1;
assign flogtanh_00033_00002 = ~I31b0f2fe98cfddbc05dbd14be8be394b+ 1;
assign flogtanh_00033_00003 = ~Ia71663e8f563041c27cd21a0c9c27a28+ 1;
assign flogtanh_00033_00004 = ~Ib46b13498ec14ceaa56719f26f18febb+ 1;
assign flogtanh_00033_00005 = ~I9bc2d5692474b8368c570d92835191b3+ 1;
assign flogtanh_00034_00000 = ~If8b0b96a659183e3651c691a2848b86b+ 1;
assign flogtanh_00034_00001 = ~I87d958c00fc6209d901147831b0c951c+ 1;
assign flogtanh_00034_00002 = ~Ie4e4eaf3e5d2f581210af8054df71c6c+ 1;
assign flogtanh_00034_00003 = ~I0b557cf102da41afd26936cbdb64b6e8+ 1;
assign flogtanh_00034_00004 = ~I49eb064043f91112c854e31e4eb9b885+ 1;
assign flogtanh_00034_00005 = ~I1039bc43e88eee527d2ed6adb8c7d1ba+ 1;
assign flogtanh_00035_00000 = ~I9aab16e89f1b64117caece8ca8af5940+ 1;
assign flogtanh_00035_00001 = ~I343df614f97cf732e57cf2ad3f95dc9e+ 1;
assign flogtanh_00035_00002 = ~Ie02de90d8eb06b16314946d21299500c+ 1;
assign flogtanh_00035_00003 = ~I3353a7916b569f2c0ca122180608dccc+ 1;
assign flogtanh_00035_00004 = ~Ibfe760474fcac99f1e5ffa2e008fef99+ 1;
assign flogtanh_00035_00005 = ~I3caf1211dcbcdc746a3e4c7fbbdae4a8+ 1;
assign flogtanh_00036_00000 = ~I2dcc0d17b9fcac35693bf32b5c5540fd+ 1;
assign flogtanh_00036_00001 = ~Ie6764a631310e312ba5c2c1e601d828f+ 1;
assign flogtanh_00036_00002 = ~I220f8e45e5fe6e69f02cded87f12e1e5+ 1;
assign flogtanh_00036_00003 = ~I896cd566a3d078b0f697a788efd223f2+ 1;
assign flogtanh_00036_00004 = ~I7caa41076a293edf18c7c4309fdcfc91+ 1;
assign flogtanh_00036_00005 = ~I928a0e4951208aab170656596f456209+ 1;
assign flogtanh_00036_00006 = ~Ia3d129fd297905bee180293c0c39d9ef+ 1;
assign flogtanh_00036_00007 = ~Id555c88cf7f0904db74d45cc75c8f5d6+ 1;
assign flogtanh_00037_00000 = ~I1ddfd31bbf062aa5c3c71d61e492e3a2+ 1;
assign flogtanh_00037_00001 = ~Iae9e023628eb6686708b2656f15616cc+ 1;
assign flogtanh_00037_00002 = ~If4b100d26126e460c41b8c1bc8fbbb96+ 1;
assign flogtanh_00037_00003 = ~I85a7fede715578be0634d71e9c7951cd+ 1;
assign flogtanh_00037_00004 = ~I2d7715a3af03d9664729fa6df85034a2+ 1;
assign flogtanh_00037_00005 = ~I571ddcb0a10938e4c0816c965214b4a8+ 1;
assign flogtanh_00037_00006 = ~I8bf8b0cf27a2654a0e7fdf3255945b67+ 1;
assign flogtanh_00037_00007 = ~I63f82f075d53205b5b556c0054f1a0b8+ 1;
assign flogtanh_00038_00000 = ~I3c6fb0df5846a19228a4e6cf9f9106ac+ 1;
assign flogtanh_00038_00001 = ~I7168b0efdd2fae57292379c9d15c62eb+ 1;
assign flogtanh_00038_00002 = ~Ibe502ebbb366f54a8f8fda4e361308e3+ 1;
assign flogtanh_00038_00003 = ~Ifce70fefde8f5ea4d2c1857236f66d65+ 1;
assign flogtanh_00038_00004 = ~Ice2c390d296e09b117d60905343e9098+ 1;
assign flogtanh_00038_00005 = ~I4b94402a53d981e953c21ef316c709b7+ 1;
assign flogtanh_00038_00006 = ~I450c0d6ad5d3b1f18bb28e3a432b5442+ 1;
assign flogtanh_00038_00007 = ~I2587a5800a5a9ffeabc4dca503e3d964+ 1;
assign flogtanh_00039_00000 = ~I1182655739d7ab5bbe4a6546a5ca36fd+ 1;
assign flogtanh_00039_00001 = ~I8110a5a62607093b21b7cd088b1d9ee0+ 1;
assign flogtanh_00039_00002 = ~I8b611f7c12ddd81de403ba74e212857f+ 1;
assign flogtanh_00039_00003 = ~I84a62a133dbceb5a32a7c907f371663d+ 1;
assign flogtanh_00039_00004 = ~Ia2fc8a1bbc3cb0dd7d89a7f05b04909c+ 1;
assign flogtanh_00039_00005 = ~I2a3eb42a4402e873d081f94a14a99c20+ 1;
assign flogtanh_00039_00006 = ~I58447d6ae49a6be2d043477a06f83df0+ 1;
assign flogtanh_00039_00007 = ~I83292bcda4645233d8e8a1dfe8e5f60b+ 1;
assign flogtanh_00040_00000 = ~Ic5e0a84cf1a2ef907b2456559ea26c75+ 1;
assign flogtanh_00040_00001 = ~I2cefbf897bb7f6f67ca500727e85c683+ 1;
assign flogtanh_00040_00002 = ~If47be2ca4617a426258c51f8d977ba3f+ 1;
assign flogtanh_00040_00003 = ~I7c68e0ae30efc4ca4d68b6047119c6c3+ 1;
assign flogtanh_00040_00004 = ~Iccca1936f4c1c9496205e77b588e9985+ 1;
assign flogtanh_00040_00005 = ~I59d4567d3355fdae5660a1364d1b8d00+ 1;
assign flogtanh_00040_00006 = ~I4600963866dcb9bbea2515c805f885cb+ 1;
assign flogtanh_00040_00007 = ~If26d90629e70c5a871e6f5b14471b8cf+ 1;
assign flogtanh_00040_00008 = ~Iedb9bb14951bf67bc8865b0983490c14+ 1;
assign flogtanh_00041_00000 = ~I6a3854ed571e8c262aa3ec377c247778+ 1;
assign flogtanh_00041_00001 = ~I05028975b49ec0c089bd981696f85a8b+ 1;
assign flogtanh_00041_00002 = ~Ife732309efcc740cfff5c747aab2e3d6+ 1;
assign flogtanh_00041_00003 = ~Idcef10a0465614cf38e0d6f503b5174a+ 1;
assign flogtanh_00041_00004 = ~Ibd4aaf02982068ffbfd1b8b3795d9217+ 1;
assign flogtanh_00041_00005 = ~I788c64785b992c675fe348a1fa181525+ 1;
assign flogtanh_00041_00006 = ~Ib235af5b28d56f24372d3f0af816f2c2+ 1;
assign flogtanh_00041_00007 = ~I4c03a6569d1b954d088053e38827e811+ 1;
assign flogtanh_00041_00008 = ~Idda26504e422367082caeafbb29871f9+ 1;
assign flogtanh_00042_00000 = ~I195c3a82123142d509886ee37dc6fc98+ 1;
assign flogtanh_00042_00001 = ~I1abb512ca0383c9e7104418e07281841+ 1;
assign flogtanh_00042_00002 = ~I00ff1331b1900bb031ee81d2a58c1bd5+ 1;
assign flogtanh_00042_00003 = ~If65eb5e743a7b1878fb232ef2fe13cb0+ 1;
assign flogtanh_00042_00004 = ~I24ae7de3549a84f4f88f561b6017b7a8+ 1;
assign flogtanh_00042_00005 = ~I449c77140475475b138d839a74078337+ 1;
assign flogtanh_00042_00006 = ~Ia9e102d8679943c079f16c0228f0f0d1+ 1;
assign flogtanh_00042_00007 = ~Ibf1c9d86665f696d91c554db748ff42b+ 1;
assign flogtanh_00042_00008 = ~Ieb0336a1974a2aec0966f4f59f460802+ 1;
assign flogtanh_00043_00000 = ~Ic0819ccefe784a6379716b3633ae0196+ 1;
assign flogtanh_00043_00001 = ~I0c4bbd1827b1859caabb067e864ce4b3+ 1;
assign flogtanh_00043_00002 = ~I004c98da87996b77b5761d366210f782+ 1;
assign flogtanh_00043_00003 = ~Ia457938da4efe847cb06f645f2a54a52+ 1;
assign flogtanh_00043_00004 = ~I7e0474089ebc1c34747be1bc17a81d72+ 1;
assign flogtanh_00043_00005 = ~Ib0b46b99e61d724ae664d9d1fec1e29f+ 1;
assign flogtanh_00043_00006 = ~I56d1025271f1f7704a40dd7f0df02b0b+ 1;
assign flogtanh_00043_00007 = ~I72c2256ba47cf03f95143df8f741fd83+ 1;
assign flogtanh_00043_00008 = ~I733c3fa4d84e5680792b16a70bb1a51d+ 1;
assign flogtanh_00044_00000 = ~If367d63311c96726517240de13bd2a4b+ 1;
assign flogtanh_00044_00001 = ~Icc6d895d943e14f2801c22e79ce190e8+ 1;
assign flogtanh_00044_00002 = ~Ieb664ac9be65fba2e25960141f7fb4b6+ 1;
assign flogtanh_00044_00003 = ~I66071f20991b414140869a2e3b750471+ 1;
assign flogtanh_00044_00004 = ~Iffeefa89a2ba7d032db5db64cbf05e20+ 1;
assign flogtanh_00044_00005 = ~I9ab3cea6ee8d8473221da21bae06066b+ 1;
assign flogtanh_00044_00006 = ~I3403ce6e697b523a9f441d8fd5e2d420+ 1;
assign flogtanh_00044_00007 = ~Ia98a70144e466b356d2998948dc4b602+ 1;
assign flogtanh_00044_00008 = ~Ie4ca0836695d951ee09622892ee35928+ 1;
assign flogtanh_00044_00009 = ~I485a48b4ff4da08f977425fd10e6d392+ 1;
assign flogtanh_00044_00010 = ~Ie8c79e6a5378808c0ead5a4b24319ce9+ 1;
assign flogtanh_00044_00011 = ~I9ca81c841a75a9ac242835956509e0fe+ 1;
assign flogtanh_00044_00012 = ~Id50f18f642f3b00ffa34986f78a0eae6+ 1;
assign flogtanh_00044_00013 = ~I75838ca09e301b8e1301cbf603a1f8c2+ 1;
assign flogtanh_00044_00014 = ~Id968b34075e351ab01d65abcb4ed8cca+ 1;
assign flogtanh_00044_00015 = ~I84da4ce7441e132e775167c1cd81dbe5+ 1;
assign flogtanh_00045_00000 = ~If19dc22d45cc4664c85a043ec4c00617+ 1;
assign flogtanh_00045_00001 = ~Ibf482db0f5058be72061267c42ebc292+ 1;
assign flogtanh_00045_00002 = ~I6d2dbb953a58b91dafa7f0d34d41bdc3+ 1;
assign flogtanh_00045_00003 = ~Ib393146d81d3cf031466543311cee2ad+ 1;
assign flogtanh_00045_00004 = ~I42564ec6a794ea803795f0b5b3523a93+ 1;
assign flogtanh_00045_00005 = ~I4a0033a180d7edce81fcfef603532e28+ 1;
assign flogtanh_00045_00006 = ~Ic7a21921e2716fba55aad2e351f4498a+ 1;
assign flogtanh_00045_00007 = ~I9a3f0b4867087790c78f674b719dbf7b+ 1;
assign flogtanh_00045_00008 = ~I138f008a6206a1067bb0e22ce3d90990+ 1;
assign flogtanh_00045_00009 = ~I48ad9b737892d7c49340ed679f46e034+ 1;
assign flogtanh_00045_00010 = ~I04a9c9765fd468a7e841577f09fc287b+ 1;
assign flogtanh_00045_00011 = ~I7b929c228c865112f00bc6b4dcc95b52+ 1;
assign flogtanh_00045_00012 = ~I2b54a135e59945901e9c11580a29ee3d+ 1;
assign flogtanh_00045_00013 = ~I566221060f06e724676ec9bec861d7de+ 1;
assign flogtanh_00045_00014 = ~Icd9a876a0feb16ea62bcad5be2004dac+ 1;
assign flogtanh_00045_00015 = ~I8f8273c4cb2a9ace8a09847efd4bdec7+ 1;
assign flogtanh_00046_00000 = ~I96ef4b631a7f63e19f67f3920685f0e6+ 1;
assign flogtanh_00046_00001 = ~I9e2de71442b8f504358e582087a6d19f+ 1;
assign flogtanh_00046_00002 = ~I1fb13d7500f5ac3821c424bd3688cf4e+ 1;
assign flogtanh_00046_00003 = ~I2aabda12ff89e708d04b4399472b5203+ 1;
assign flogtanh_00046_00004 = ~I8c733a5d394e6b8d045eede5cc7451f6+ 1;
assign flogtanh_00046_00005 = ~I4f45dd50d2825ab338b8a2a8264096c0+ 1;
assign flogtanh_00046_00006 = ~Ib45caf6b563d22144be3e9225a99a1cd+ 1;
assign flogtanh_00046_00007 = ~I9d6730140c690037b5ca58aa30103f5b+ 1;
assign flogtanh_00046_00008 = ~I9df5b63f66c162d517daa69f5d0e6095+ 1;
assign flogtanh_00046_00009 = ~I1b40adfd6fa6c943dfa8d230d9e65514+ 1;
assign flogtanh_00046_00010 = ~I0eb3df4d4094e09e6c4b3c788baed61f+ 1;
assign flogtanh_00046_00011 = ~Id6f7923a16cc5adc96a730083153ca6d+ 1;
assign flogtanh_00046_00012 = ~Idf8ebc0d747ae143aa61866e33d458c0+ 1;
assign flogtanh_00046_00013 = ~Id682e531735437bc24abbf3d3d51e18b+ 1;
assign flogtanh_00046_00014 = ~I05ecce409cca00ea5b0df25de5a50cf2+ 1;
assign flogtanh_00046_00015 = ~I831d214dcb4f8d534b5ddaaeaeeb81ce+ 1;
assign flogtanh_00047_00000 = ~Ia540866403683bc30504bace19bdda7b+ 1;
assign flogtanh_00047_00001 = ~I05fb1982415bd3fa78dd9a00af7a3d4a+ 1;
assign flogtanh_00047_00002 = ~I977864efb0d94149cce7dc4d165f11de+ 1;
assign flogtanh_00047_00003 = ~I9362b615a612599239e3b752a9334e8c+ 1;
assign flogtanh_00047_00004 = ~I5d4fb4b5a5ad3dc48beebfa0e0cebbed+ 1;
assign flogtanh_00047_00005 = ~Ifb9b29c43f435452cc761218c509f5df+ 1;
assign flogtanh_00047_00006 = ~If2143db72bf9a02b64eb45b3a4faa39d+ 1;
assign flogtanh_00047_00007 = ~Ice780b1695a8e80607a03dee3c426ffe+ 1;
assign flogtanh_00047_00008 = ~I90b0296f5ef87dfaa6110fc2e9d6ed9d+ 1;
assign flogtanh_00047_00009 = ~Icd37da8ea84a606529e32b2db4eb7f5f+ 1;
assign flogtanh_00047_00010 = ~Ie626a24e3680f7d3995dd0c2ce60cbcc+ 1;
assign flogtanh_00047_00011 = ~Iebee55168fb47664095b11c9f6641124+ 1;
assign flogtanh_00047_00012 = ~Ic0954671eb1dc893c3932e456800fadf+ 1;
assign flogtanh_00047_00013 = ~Ia4131464996aabab8aae1db85f6a50e4+ 1;
assign flogtanh_00047_00014 = ~I2de1ca2c390bdd3011fff4a359bb5332+ 1;
assign flogtanh_00047_00015 = ~I6fb55222b69475b7168874423226ec9c+ 1;
assign flogtanh_00048_00000 = ~I9b09b800a9dcd8ac36f25cb0324e748d+ 1;
assign flogtanh_00048_00001 = ~I74ac0327175f50f508a5013df298df02+ 1;
assign flogtanh_00048_00002 = ~Ica26f542586d50c56ce0f3c00f36b388+ 1;
assign flogtanh_00048_00003 = ~I7c6862830daffc98cb2c1fc121d82c38+ 1;
assign flogtanh_00048_00004 = ~Icf19dd665616a8c96146b3ab9f46c741+ 1;
assign flogtanh_00048_00005 = ~I97f2813ec39bbf1513faf66b3e38838a+ 1;
assign flogtanh_00048_00006 = ~I716ee53e79883f69aa045380a357e913+ 1;
assign flogtanh_00048_00007 = ~I25c324feaca84e80f58075597e8c448f+ 1;
assign flogtanh_00048_00008 = ~I7fc190647082a3d71614f46f670167bc+ 1;
assign flogtanh_00049_00000 = ~Iebdf938a28594624f4d4a337356485cb+ 1;
assign flogtanh_00049_00001 = ~I3fd068d55154441ffd005999ea823fd0+ 1;
assign flogtanh_00049_00002 = ~Ic5ca74b66763c6e5591c7c2bfeeb0663+ 1;
assign flogtanh_00049_00003 = ~I5ab556386d2973354a5551ba9823e4ba+ 1;
assign flogtanh_00049_00004 = ~I64f65df774d29696425ba460dda09b68+ 1;
assign flogtanh_00049_00005 = ~I9e09c25be9f877c1e1aaf79bf12c7943+ 1;
assign flogtanh_00049_00006 = ~I42c1d469ff97913cbf15e3ebee6fdfa8+ 1;
assign flogtanh_00049_00007 = ~If9f2a53dbf6e9b9a335a7657b7a2b468+ 1;
assign flogtanh_00049_00008 = ~I495f8be463b15db906474c518e0741e2+ 1;
assign flogtanh_00050_00000 = ~I3e265a7dcf29687248b9275df49771fb+ 1;
assign flogtanh_00050_00001 = ~Iffd94cf3a8a4681ff3327c90bf89bd8b+ 1;
assign flogtanh_00050_00002 = ~Iea71417e738c6ca54c50aa014cc38627+ 1;
assign flogtanh_00050_00003 = ~Ic8df04756f67e6dd29f3374c5f86d451+ 1;
assign flogtanh_00050_00004 = ~I546122346a22ad64a6ab2b4978cde095+ 1;
assign flogtanh_00050_00005 = ~Icaae0fb0f460f68d690ab00697355a49+ 1;
assign flogtanh_00050_00006 = ~I42455e7e4d0c63f97702d204d18a446e+ 1;
assign flogtanh_00050_00007 = ~Iaec2f15665e83416bc140890f3cdde9a+ 1;
assign flogtanh_00050_00008 = ~I487391402b6aa27bf212724a37ea9c33+ 1;
assign flogtanh_00051_00000 = ~Ia9f375709014a9d553d46cff2799b59f+ 1;
assign flogtanh_00051_00001 = ~I34d428a56bd0142a9be9f627f1c3c87f+ 1;
assign flogtanh_00051_00002 = ~I57db98eb439d59a895dabe029c6a3a8b+ 1;
assign flogtanh_00051_00003 = ~I9937af6fcf9d834f308bc3683d524981+ 1;
assign flogtanh_00051_00004 = ~I463f4f370e1ecad71de44780eff10df4+ 1;
assign flogtanh_00051_00005 = ~I53309409a6059c3bd39f037c23ec3458+ 1;
assign flogtanh_00051_00006 = ~I2603e0b8b93f6680e44c9c8883f6512c+ 1;
assign flogtanh_00051_00007 = ~Iab354cc9ac1173335c0efeef694f3567+ 1;
assign flogtanh_00051_00008 = ~I6c19936ca2edeb0e261e880a1055e964+ 1;
assign flogtanh_00052_00000 = ~Ifebfa58419ecd22a334ed4b67f5c3581+ 1;
assign flogtanh_00052_00001 = ~I71a28e8525f07dabeabe4b4f45f353d0+ 1;
assign flogtanh_00052_00002 = ~I514830acdad20c4ff3d078477e939b4b+ 1;
assign flogtanh_00052_00003 = ~I036342f6be0f2e2f1f4927099a5c4a78+ 1;
assign flogtanh_00052_00004 = ~Iedb655aa25e5f0e35137ec6c3acdc527+ 1;
assign flogtanh_00052_00005 = ~I0c59e8c82a31aacbf5977ff778a7ff49+ 1;
assign flogtanh_00052_00006 = ~I1b6d20c64b9f23fb6c30f723546aa285+ 1;
assign flogtanh_00052_00007 = ~I0d66aa55747362354aa81d96057bc4c2+ 1;
assign flogtanh_00052_00008 = ~I1ea33707e40a2e41513fdb3118371437+ 1;
assign flogtanh_00052_00009 = ~I68c85727adecde0aa8aa66ed08c4b502+ 1;
assign flogtanh_00052_00010 = ~Iebd050e29044153d5881ef80b2db8c28+ 1;
assign flogtanh_00052_00011 = ~I3c057d64cf4fca0238a874f0ced99c76+ 1;
assign flogtanh_00053_00000 = ~I066cd52173ec5dbce9a3f470d73325af+ 1;
assign flogtanh_00053_00001 = ~Ic7ad59f6a232a997706d17b4098e0324+ 1;
assign flogtanh_00053_00002 = ~Icf8cfc800f0a2aa5140a7f83f035b0cc+ 1;
assign flogtanh_00053_00003 = ~I6bfbf7ff79ff0a6facc9ba5031239644+ 1;
assign flogtanh_00053_00004 = ~I78ade92efd265027807c861be44a10af+ 1;
assign flogtanh_00053_00005 = ~I2bc5a10c587d89d10021aa5eaafb490a+ 1;
assign flogtanh_00053_00006 = ~I30080cc6c03bbe933165d266558a822c+ 1;
assign flogtanh_00053_00007 = ~I7e28234bdf66ab5489d36d15678db797+ 1;
assign flogtanh_00053_00008 = ~I74b3c9dd3a8168aacd4369b9ff68fdfd+ 1;
assign flogtanh_00053_00009 = ~Ia7046faae1ab05978e4b32bd44049fb9+ 1;
assign flogtanh_00053_00010 = ~I0c5250aaca86185fed5978438c8861b6+ 1;
assign flogtanh_00053_00011 = ~Ic78949e07e643f571f23df7e8f15d9fb+ 1;
assign flogtanh_00054_00000 = ~Ifb8b3586a5b69b20cf03eabf51344ab6+ 1;
assign flogtanh_00054_00001 = ~I9ea09f27ce4484f2e7fc3a6b6d6ecb7c+ 1;
assign flogtanh_00054_00002 = ~If0b9225e759438be175c4128c78605ea+ 1;
assign flogtanh_00054_00003 = ~I33d941ad9d4858fcfb77f0f6cf99d2ec+ 1;
assign flogtanh_00054_00004 = ~Ia0868eee7e7e0640ce1a4d3ca9c001cb+ 1;
assign flogtanh_00054_00005 = ~Icb3ab2c67a87b2ee158e0021b72fc186+ 1;
assign flogtanh_00054_00006 = ~I5b64997d083769666741c794dd92fb7f+ 1;
assign flogtanh_00054_00007 = ~I0a3323aac825506435068f6746aee974+ 1;
assign flogtanh_00054_00008 = ~Ibec442c099da091afcf75a7c970bf8ea+ 1;
assign flogtanh_00054_00009 = ~If3a79ede332c39a8d2a276de833242f6+ 1;
assign flogtanh_00054_00010 = ~I49ccb3e14fe61618806e791ecb4f4eae+ 1;
assign flogtanh_00054_00011 = ~I461ebbf3a02ae63e2eb27531b1370f24+ 1;
assign flogtanh_00055_00000 = ~Ice66c108aa66981051df71e226cb0e4d+ 1;
assign flogtanh_00055_00001 = ~I645ff0d8c0a87ba7f792fc83f342b958+ 1;
assign flogtanh_00055_00002 = ~Ica94017f26e96fb22a47add326ee126e+ 1;
assign flogtanh_00055_00003 = ~Id32e7ad5b1aa825732d9b26d0fa02ca1+ 1;
assign flogtanh_00055_00004 = ~I51b5e641856239367cf43f9b5679b268+ 1;
assign flogtanh_00055_00005 = ~I2d1a5645b126761fc7fb70d24e37189a+ 1;
assign flogtanh_00055_00006 = ~I49f5f87662fbb540d72c94bfd1acd060+ 1;
assign flogtanh_00055_00007 = ~I30253dc91301ca27b5732312c01145e0+ 1;
assign flogtanh_00055_00008 = ~I143f5e324716a94d24ada126886bf895+ 1;
assign flogtanh_00055_00009 = ~If64aa8c220b9ab6652e081da7e404e80+ 1;
assign flogtanh_00055_00010 = ~I1092325b801600fa7ec85fa640167da9+ 1;
assign flogtanh_00055_00011 = ~Ib028686da9c849e827cf249a744b7db3+ 1;
assign flogtanh_00056_00000 = ~I5f3ff7fa8686f7a380302d71b88cfb4b+ 1;
assign flogtanh_00057_00000 = ~Ic01904f7c518990eff2dc1de127676c4+ 1;
assign flogtanh_00058_00000 = ~I43f2ddd9780f86af489f8deae51168ec+ 1;
assign flogtanh_00059_00000 = ~I0a013fff6c792363bd7feb03d9691db8+ 1;
assign flogtanh_00060_00000 = ~I7cf8401bf6893eab0b9f33a0f91ddd05+ 1;
assign flogtanh_00061_00000 = ~Ic7ccbeaf4ab94d0660eb7a0533723e24+ 1;
assign flogtanh_00062_00000 = ~I08043393cb7f2558c145a698ea6652c9+ 1;
assign flogtanh_00063_00000 = ~I84865c4f872c0845124b78fabf695c2c+ 1;
assign flogtanh_00064_00000 = ~I57b9dd7a7deea6695dcd03439c9723cf+ 1;
assign flogtanh_00065_00000 = ~I1cd6b35bcdfd461db69a4c1bdb1d387f+ 1;
assign flogtanh_00066_00000 = ~I40a1ecabded8add5bffe316f2d8beda9+ 1;
assign flogtanh_00067_00000 = ~I7c52ae4af926267b5e27a530202fcce0+ 1;
assign flogtanh_00068_00000 = ~I1a5c6c50817db8bde279d5f0b5095d76+ 1;
assign flogtanh_00069_00000 = ~Idf0c1b85712fcbbbcc12915158ebff62+ 1;
assign flogtanh_00070_00000 = ~I6b32298e8c61e75d0a38bca3084c0528+ 1;
assign flogtanh_00071_00000 = ~I5b0d72cedc120406402076148e2d30b0+ 1;
assign flogtanh_00072_00000 = ~Iaf624549f73b0d13c1a73c850b99f810+ 1;
assign flogtanh_00073_00000 = ~Iaaf7efeae9f6dc9e8222dc2b10122000+ 1;
assign flogtanh_00074_00000 = ~Iea1cd2321d2ac9b891b344e2ba2363d3+ 1;
assign flogtanh_00075_00000 = ~Ia544fa24b953fe91800978895e3e610e+ 1;
assign flogtanh_00076_00000 = ~I7fa710c37f5f96c3cdc35612a702a71c+ 1;
assign flogtanh_00077_00000 = ~I98fd105696fca11c1075f9bd30013747+ 1;
assign flogtanh_00078_00000 = ~I61345963ceabdaa0f25f8a463fc9fe5d+ 1;
assign flogtanh_00079_00000 = ~I9e8375af6af10f4bac3e87e416d430ee+ 1;
assign flogtanh_00080_00000 = ~Ida1cd844022bbf1b8431225e66b2b78f+ 1;
assign flogtanh_00081_00000 = ~I30e9ab592e97dbc5fb6ab58d2ffbf8d4+ 1;
assign flogtanh_00082_00000 = ~I2ec2a6de2be39b1bc259b0be72e35a0f+ 1;
assign flogtanh_00083_00000 = ~Ic32e349efae2ca419e095ee5e15a501d+ 1;
assign flogtanh_00084_00000 = ~I1befb935ee9cb871c9a7476c1fc0da3f+ 1;
assign flogtanh_00085_00000 = ~I01c57f697f2af7d2c6ae904319f10725+ 1;
assign flogtanh_00086_00000 = ~Id580f8a2748efff9b6b747c497c16e9c+ 1;
assign flogtanh_00087_00000 = ~I77b54488bd26318f14b4364035cd1836+ 1;
assign flogtanh_00088_00000 = ~I786338397f55073dce91e1c8c5f8e298+ 1;
assign flogtanh_00089_00000 = ~I0e5931219d94c8e8e1f4af081404dcab+ 1;
assign flogtanh_00090_00000 = ~I8d96b419b010f8076311420d7b9c8a18+ 1;
assign flogtanh_00091_00000 = ~Ife13f962c7a8df3845cde104a959f678+ 1;
assign flogtanh_00092_00000 = ~I7f701ff37ad3fc34d2f4efafe5ff5351+ 1;
assign flogtanh_00093_00000 = ~I43c815a8ce0b2df9744a525328969691+ 1;
assign flogtanh_00094_00000 = ~I6c4a1ded9bf39091cf302ebe0103e2f0+ 1;
assign flogtanh_00095_00000 = ~Icd4ff8d14af2699db2b5168027894ebb+ 1;
assign flogtanh_00096_00000 = ~Ia79d52fe2130426c07890fcaa50137db+ 1;
assign flogtanh_00097_00000 = ~I308aaa8ac500b5589aa4af533a9062bf+ 1;
assign flogtanh_00098_00000 = ~Iac91f4037e542d9fda30fadafe7e79ac+ 1;
assign flogtanh_00099_00000 = ~I8cd5970682bc84881489c12ff073212c+ 1;
assign flogtanh_00100_00000 = ~I1ee27be7e1a38aff0039b21c45f406d1+ 1;
assign flogtanh_00101_00000 = ~Idf90f01353ad1057e11fd060442f4e53+ 1;
assign flogtanh_00102_00000 = ~Id45f4e0f142b6c3925f24a37dcf7c0ae+ 1;
assign flogtanh_00103_00000 = ~I52a9bcfbd2d3a763671f19cfeaf7bb8b+ 1;
assign flogtanh_00104_00000 = ~Ia3cc6acf2cae41e560e09993007ffd2b+ 1;
assign flogtanh_00105_00000 = ~Iba0d2f08788f2208a648ae7b5414195d+ 1;
assign flogtanh_00106_00000 = ~I9f7df6ad60284c812aeb522974578e0b+ 1;
assign flogtanh_00107_00000 = ~Iab1fb7006598181bd8749ed90c519b13+ 1;
assign flogtanh_00108_00000 = ~Ieef3b299ec35075c71ef9fb10525bfc4+ 1;
assign flogtanh_00109_00000 = ~I58a7c08adf48d0737c5803e2a818c045+ 1;
assign flogtanh_00110_00000 = ~I30a1c8fcd9a510a6ed559f07dd809b90+ 1;
assign flogtanh_00111_00000 = ~Ic4f5e9d49419e1c57cfa387761ab643d+ 1;
assign flogtanh_00112_00000 = ~Id3dd71ea0bf0f2996fbe42b8c3318762+ 1;
assign flogtanh_00113_00000 = ~Ib834b91bf81067e8efa9d470023e8b9d+ 1;
assign flogtanh_00114_00000 = ~Ic6ead78ed741442f17a15a157cd6ef9c+ 1;
assign flogtanh_00115_00000 = ~I4e257dbd6f196a02dc0f5a2e5f6047d7+ 1;
assign flogtanh_00116_00000 = ~I3dbfbd34d1fdfd4f422d900154123b6b+ 1;
assign flogtanh_00117_00000 = ~I529b763dace1924613d184c6c70c2708+ 1;
assign flogtanh_00118_00000 = ~I7a600aeb6cf8c3311c10afa4d82767a1+ 1;
assign flogtanh_00119_00000 = ~I8c7aab31f8cb705ea13a41a5bd349303+ 1;
assign flogtanh_00120_00000 = ~I171149dcaab2c0f0e2a10547ad95084d+ 1;
assign flogtanh_00121_00000 = ~I23b60ca4da2df0ec40c1df62d058deef+ 1;
assign flogtanh_00122_00000 = ~I7978d2d800b4438d0644ae3df6bcac9c+ 1;
assign flogtanh_00123_00000 = ~Ibc4eddc0f1768e9ec7e38e951a28ec42+ 1;
assign flogtanh_00124_00000 = ~I1c97fd1d21a31af8b5498a79b1a3e7b6+ 1;
assign flogtanh_00125_00000 = ~Ie4f063eeaf7ee3f033e2a01ffaca623e+ 1;
assign flogtanh_00126_00000 = ~Ibb3d57d510cad00064a331f61f6400a2+ 1;
assign flogtanh_00127_00000 = ~I9485ae915474a31562ce358666d66245+ 1;
assign flogtanh_00128_00000 = ~Ia54b6f7044a831020e49f1bf48bc063a+ 1;
assign flogtanh_00129_00000 = ~Ie71c7babb5d17378d40444b6bbd4e7a6+ 1;
assign flogtanh_00130_00000 = ~Ia0977b79857bdbf058535c30e338c38a+ 1;
assign flogtanh_00131_00000 = ~I600ea1371a2be66430ac9534583b512b+ 1;
assign flogtanh_00132_00000 = ~Ife5b9afdbb30c122b84d5378f9cb366d+ 1;
assign flogtanh_00133_00000 = ~I27556d599dd1a27ee8f49e819ccbf29a+ 1;
assign flogtanh_00134_00000 = ~Icce595233ce089eafcca3eae5e71e5f8+ 1;
assign flogtanh_00135_00000 = ~Icc3cadf40c09be1a8c2847caf0e3e63c+ 1;
assign flogtanh_00136_00000 = ~Ib43886d923b8c683004713ff25b2f90d+ 1;
assign flogtanh_00137_00000 = ~I132d9671c582876568c0f7f5335f5227+ 1;
assign flogtanh_00138_00000 = ~I0859c80b42a8c60dade8f05d58ee3701+ 1;
assign flogtanh_00139_00000 = ~Ib3690ec149adde94343d3e617931a287+ 1;
assign flogtanh_00140_00000 = ~I41f2bf9ff00f983ad1298c8c83b041cb+ 1;
assign flogtanh_00141_00000 = ~Ib5414585cd6976cfce42e42190cc08d7+ 1;
assign flogtanh_00142_00000 = ~I1ca59325ff30db83df5bf0a2cd9706b6+ 1;
assign flogtanh_00143_00000 = ~Ie2f5b03f3b136e651b8aba92a30d298a+ 1;
assign flogtanh_00144_00000 = ~I312ce79a8dd2ce3d37c930d42640509b+ 1;
assign flogtanh_00145_00000 = ~I467d5e2554ef25873e0b44e947ee0011+ 1;
assign flogtanh_00146_00000 = ~Ice73b514709469fd21cd254bf4ceadd9+ 1;
assign flogtanh_00147_00000 = ~I45ba06a6d6f00c174b1439a6f226a085+ 1;
assign flogtanh_00148_00000 = ~Ic8a272f82736fd599fb3250e970edf9b+ 1;
assign flogtanh_00149_00000 = ~I5b9710b16effc8bf0695517c6e651836+ 1;
assign flogtanh_00150_00000 = ~I038b42a83025f5eaebf45799d1ebe7b0+ 1;
assign flogtanh_00151_00000 = ~I73ddd7cf9272ceab5a663e2244e72d7e+ 1;
assign flogtanh_00152_00000 = ~I16507fab8f9076bfeb419896fa7cdc1d+ 1;
assign flogtanh_00153_00000 = ~I3dd1f28cf199299aba54e47a429c9b11+ 1;
assign flogtanh_00154_00000 = ~I49d9203dc6f8c17f17383e8f7e01f005+ 1;
assign flogtanh_00155_00000 = ~Ibeec86c75d950ee00dd63a2930f08a24+ 1;
assign flogtanh_00156_00000 = ~I47b2438c3680b2d816168df37d7c491c+ 1;
assign flogtanh_00157_00000 = ~I5983bf2c6c90b872ee6cf58b5e520311+ 1;
assign flogtanh_00158_00000 = ~I6745cacecb7ee86cf3c7ad7eeee6048f+ 1;
assign flogtanh_00159_00000 = ~Ib9672d20643d856ff31905ab14c0ac87+ 1;
assign flogtanh_00160_00000 = ~Ib9dfea1f34a120eda30d5bd919365a6a+ 1;
assign flogtanh_00161_00000 = ~Ia7bf82c9e5ca4467b5e50beeaeb975e9+ 1;
assign flogtanh_00162_00000 = ~I327c9acb8934729b4ea5486787afa2e8+ 1;
assign flogtanh_00163_00000 = ~Ieddef08050c38d07e5d38f5bb7b099c0+ 1;
assign flogtanh_00164_00000 = ~I39f9e8430db114991bfb27cc46ef3e39+ 1;
assign flogtanh_00165_00000 = ~I56aa548618a4a15e9a35e04f5eeb823f+ 1;
assign flogtanh_00166_00000 = ~I1908897b529ca04df7e7da395be4a8ce+ 1;
assign flogtanh_00167_00000 = ~Ib2bbd59cd6098608ed53ac556036534f+ 1;
assign flogtanh_00168_00000 = ~If004552b2047ab1cf23bb50375460b01+ 1;
assign flogtanh_00169_00000 = ~If97092e1e2147de199c94a23831cf6b9+ 1;
assign flogtanh_00170_00000 = ~Ibf74a4dfaab7f7f538d2b5fac7394b63+ 1;
assign flogtanh_00171_00000 = ~I991a7a7d562eb0a8b4b8d8f008ef2225+ 1;
assign flogtanh_00172_00000 = ~I64c3d7be41abaa17d6992f9af8e72789+ 1;
assign flogtanh_00173_00000 = ~Icb91e63ebabc7a75a54eb7c731df4fa0+ 1;
assign flogtanh_00174_00000 = ~I673d1d0d0daab99bd940c46cc14ef55a+ 1;
assign flogtanh_00175_00000 = ~I62cadbd70b07a6a7a2974c7c392696b3+ 1;
assign flogtanh_00176_00000 = ~Icd8257d7f53d93db989eb56eaeb7e593+ 1;
assign flogtanh_00177_00000 = ~I05931ceae6eff26e5a66a44a54d628ae+ 1;
assign flogtanh_00178_00000 = ~I306fec0aa68a0396053a6e0fa1cda38f+ 1;
assign flogtanh_00179_00000 = ~Idee8c8144207d676d1f2f9064bbdff45+ 1;
assign flogtanh_00180_00000 = ~I5855124d566af739caa6511f8598f2c5+ 1;
assign flogtanh_00181_00000 = ~I50729db4a8e04f18979707df14cb2419+ 1;
assign flogtanh_00182_00000 = ~Ia3cb3ea64576a3e7332e1fb55953aa3e+ 1;
assign flogtanh_00183_00000 = ~I3cb1f233951d49f985b0deac6e052bfd+ 1;
assign flogtanh_00184_00000 = ~I7015def91103398e54f446ce3e43af01+ 1;
assign flogtanh_00185_00000 = ~I04874bd1bf257f205b5189c8c20e5a12+ 1;
assign flogtanh_00186_00000 = ~I937e3a8ede2305ea7c1750283224a870+ 1;
assign flogtanh_00187_00000 = ~Ia7206430a739a11af4d860096eedd6c3+ 1;
assign flogtanh_00188_00000 = ~Ibf4c2c00f8e012e9498361bfd3c5b06e+ 1;
assign flogtanh_00189_00000 = ~I899e5f03cd1d52d11f898959559aaeea+ 1;
assign flogtanh_00190_00000 = ~I59c80c7ec26f43308b1a646c47160568+ 1;
assign flogtanh_00191_00000 = ~I8a954a331d36266465a0813d2e8b319b+ 1;
assign flogtanh_00192_00000 = ~Ib49e53ca8efd9564ee9572eb3089bb51+ 1;
assign flogtanh_00193_00000 = ~Icbde2c6230e9cc67ef12031e38bb344f+ 1;
assign flogtanh_00194_00000 = ~I2e22e867f6f84a7807b82f64a147022e+ 1;
assign flogtanh_00195_00000 = ~Id9704e1d8096cd28577c5c357d30b7a4+ 1;
assign flogtanh_00196_00000 = ~I4b8554cab486a4fc1e14884a6495016e+ 1;
assign flogtanh_00197_00000 = ~Iaa235d085a5916a3b0814c3ed2a9026f+ 1;
assign flogtanh_00198_00000 = ~I5d86ce0b58c0b281d747116a9069ef33+ 1;
assign flogtanh_00199_00000 = ~Id20394136fb036435bb4680aac64581f+ 1;
assign flogtanh_00200_00000 = ~I8a16afac6e470ca69634d7fe9656387a+ 1;
assign flogtanh_00201_00000 = ~Ic4e7f690bc050f1d1f84eae7ca193e1c+ 1;
assign flogtanh_00202_00000 = ~Ia60421aa427236540b4d0d08d52ff507+ 1;
assign flogtanh_00203_00000 = ~Icace650ee3865bd7bbddd2d9435c5561+ 1;
assign flogtanh_00204_00000 = ~I7d27d070b96b7810f667e1d1845342d3+ 1;
assign flogtanh_00205_00000 = ~Ida7ec09c913caa0e78a2c4cbaae517c8+ 1;
assign flogtanh_00206_00000 = ~Ic5eba898858be1f768841ead792d6d86+ 1;
assign flogtanh_00207_00000 = ~I72197797a307c611fa8952533e63d7bf+ 1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00000_U (
.flogtanh_sel( Ic93835a022c46b7aa00a465c407d7da2[flogtanh_SEL-1:0]),
.flogtanh( Ia67805b59c3011bc4fc5cb1d2996f90d),
.start_in(start_d3),
.start_out(start_d4),
.rstn(rstn),
.clk(clk)
);

assign I0313213a8c479f77e683ce3fa232450c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia67805b59c3011bc4fc5cb1d2996f90d };
assign I5f68368511b59d2e365cc91b806b334e = (Ic93835a022c46b7aa00a465c407d7da2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0313213a8c479f77e683ce3fa232450c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00001_U (
.flogtanh_sel( I2e30088bf29cedd7debc15b1e6ec4ada[flogtanh_SEL-1:0]),
.flogtanh( I61fb47b07547e09c746b1fb5d7c8710d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iad493302f9a77b86d5db79901fcf4a49  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I61fb47b07547e09c746b1fb5d7c8710d };
assign I71e4d98dca37256fcc84248a26d703e2 = (I2e30088bf29cedd7debc15b1e6ec4ada[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iad493302f9a77b86d5db79901fcf4a49;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00002_U (
.flogtanh_sel( I38f512bfb84094d1e92a10a345d5505f[flogtanh_SEL-1:0]),
.flogtanh( Ib2220549c84e87683ccf85798b2bb22f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If50382087360c9884aa683e4e94bcab8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib2220549c84e87683ccf85798b2bb22f };
assign Ib8380902ac4082f834744ddef6d0cc6a = (I38f512bfb84094d1e92a10a345d5505f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If50382087360c9884aa683e4e94bcab8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00003_U (
.flogtanh_sel( I1e878f00f056f637625cb013a93325a8[flogtanh_SEL-1:0]),
.flogtanh( I12f063ad18938c2ca008e1165f9119e9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I549ce8de585aa301a4e144342ed29fc6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I12f063ad18938c2ca008e1165f9119e9 };
assign I9570f8498d95bee230bb3c5e720bb857 = (I1e878f00f056f637625cb013a93325a8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I549ce8de585aa301a4e144342ed29fc6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00004_U (
.flogtanh_sel( I25db27464b31fee41ccd7a3cfe4d403e[flogtanh_SEL-1:0]),
.flogtanh( Iae6b4023f9f2641ca00636181f4fb028),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8af1960c06a98594d58b64b42421b21b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iae6b4023f9f2641ca00636181f4fb028 };
assign I55c425102db0a6838012a165c0597680 = (I25db27464b31fee41ccd7a3cfe4d403e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8af1960c06a98594d58b64b42421b21b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00005_U (
.flogtanh_sel( I19417a224c5cdf1211e9790aa29c4c5c[flogtanh_SEL-1:0]),
.flogtanh( Id11b7d1aeb413fd4920ef0e0097fc6c4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I76b14b396d6e5193cc059e68cbd400bd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id11b7d1aeb413fd4920ef0e0097fc6c4 };
assign Ic970a88c435a85d21ed71c6060b8a8e4 = (I19417a224c5cdf1211e9790aa29c4c5c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I76b14b396d6e5193cc059e68cbd400bd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00006_U (
.flogtanh_sel( I16dcafa854ea9c67d8a080feb2ba9166[flogtanh_SEL-1:0]),
.flogtanh( I3af03d3e0bb7e0e73e034dceda70ff3a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8c0c834150ae5da887ab265f0f5b2982  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3af03d3e0bb7e0e73e034dceda70ff3a };
assign Iec8dc328edd6cbaa2d697e05ed222746 = (I16dcafa854ea9c67d8a080feb2ba9166[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8c0c834150ae5da887ab265f0f5b2982;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00007_U (
.flogtanh_sel( I7f63338eee2663fbe61fffd248433310[flogtanh_SEL-1:0]),
.flogtanh( Iba30a494dc1b66bd2862f82c16017a99),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I79934362360a11c365095cfa70a112a1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iba30a494dc1b66bd2862f82c16017a99 };
assign I16d2084ccfb102c3bafc701872f5ef2d = (I7f63338eee2663fbe61fffd248433310[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I79934362360a11c365095cfa70a112a1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00008_U (
.flogtanh_sel( Icb1e3c56c8729c32d43c69710e345db2[flogtanh_SEL-1:0]),
.flogtanh( Iefa075dc743d616eca65f76d2c03371c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I65d0cff1828f6d8ba153cadd058a8672  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iefa075dc743d616eca65f76d2c03371c };
assign Id680a9affed622577164b3a8380494f5 = (Icb1e3c56c8729c32d43c69710e345db2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I65d0cff1828f6d8ba153cadd058a8672;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00009_U (
.flogtanh_sel( I6ece8e3c1e89613879336936f77d732f[flogtanh_SEL-1:0]),
.flogtanh( Icc7a632da404a9cda7b8247706391f85),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8a4669217f831b4e42875fea28da24fd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icc7a632da404a9cda7b8247706391f85 };
assign Ifcd68be4bea38622d2d57d3a4e6fc5bb = (I6ece8e3c1e89613879336936f77d732f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8a4669217f831b4e42875fea28da24fd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00010_U (
.flogtanh_sel( I72a646ae7e32a16af0f5930a6e95b36a[flogtanh_SEL-1:0]),
.flogtanh( I708c5d8d6d8f7f16c2f348c3b97b906d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ife6c86fee255f30215fca193d9288a8e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I708c5d8d6d8f7f16c2f348c3b97b906d };
assign I16deb9107193a3536979e4b5e5654b9c = (I72a646ae7e32a16af0f5930a6e95b36a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ife6c86fee255f30215fca193d9288a8e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00011_U (
.flogtanh_sel( I7e72d119dd93a6ab05a23fde0a865866[flogtanh_SEL-1:0]),
.flogtanh( I51ba1e25e01c39a77559089626bafa09),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id8e7f39e4cdcd6d7e1ee2c8f6cce1e46  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I51ba1e25e01c39a77559089626bafa09 };
assign I28cac65a4db3f708cc90a1b023bfe894 = (I7e72d119dd93a6ab05a23fde0a865866[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id8e7f39e4cdcd6d7e1ee2c8f6cce1e46;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00012_U (
.flogtanh_sel( Ied4fdf5805039cd2fcd042fd13755fdc[flogtanh_SEL-1:0]),
.flogtanh( I2217e483aaf5124d9beb9baf5037326b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8c394ac9f9f7e5d96afde79240c0744f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2217e483aaf5124d9beb9baf5037326b };
assign Ie763738b7faf253837e1c45de255cb5e = (Ied4fdf5805039cd2fcd042fd13755fdc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8c394ac9f9f7e5d96afde79240c0744f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00013_U (
.flogtanh_sel( Id44c2293b765cff450dd1d747c47c1f3[flogtanh_SEL-1:0]),
.flogtanh( Ib47f8220e7a319e690649f9d6cc9f0cc),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4ab5a06a58aa9b4d293e73712d7a21e7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib47f8220e7a319e690649f9d6cc9f0cc };
assign Icfef12499b53cd84f0aae067f30c17d0 = (Id44c2293b765cff450dd1d747c47c1f3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4ab5a06a58aa9b4d293e73712d7a21e7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00014_U (
.flogtanh_sel( I8f4ed02f7aeb823b745040f7f3f43ac7[flogtanh_SEL-1:0]),
.flogtanh( Iffc502b536d88d080c59eb3aedd55bd1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib09e4bab1aeb88aa15f375adc930c9c8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iffc502b536d88d080c59eb3aedd55bd1 };
assign I0982b8d7f99aceb8871c9c10448f54c5 = (I8f4ed02f7aeb823b745040f7f3f43ac7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib09e4bab1aeb88aa15f375adc930c9c8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00015_U (
.flogtanh_sel( I6488b9b8f405d7d81a4874fab2678102[flogtanh_SEL-1:0]),
.flogtanh( Iaa823b6b13acb376f979dd52683a2231),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifd56f5082b3fb8406b4c07761d1d61b9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iaa823b6b13acb376f979dd52683a2231 };
assign I6c661048307c23c699d4b3636564de0f = (I6488b9b8f405d7d81a4874fab2678102[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifd56f5082b3fb8406b4c07761d1d61b9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00016_U (
.flogtanh_sel( Ifff612d16828ec907a348479e19ddf31[flogtanh_SEL-1:0]),
.flogtanh( Ic5f3f371b1ebfe733404b4165fe746dc),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1a7d739018ade49afeb6fbbf0315070d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic5f3f371b1ebfe733404b4165fe746dc };
assign I786dfcaa131b99c254aaff15bd2c2b6d = (Ifff612d16828ec907a348479e19ddf31[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1a7d739018ade49afeb6fbbf0315070d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00017_U (
.flogtanh_sel( I268262076f22bc6b1507bc8f91b98a0a[flogtanh_SEL-1:0]),
.flogtanh( I021d991730d154218106f00e74bf9d4c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I25c7e7936b9c7b257e5766618159b29d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I021d991730d154218106f00e74bf9d4c };
assign I2b49d74cb130542f2ca99534e2c513b1 = (I268262076f22bc6b1507bc8f91b98a0a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I25c7e7936b9c7b257e5766618159b29d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00018_U (
.flogtanh_sel( If1f732841adb7c0cad1ba37c0f5fd517[flogtanh_SEL-1:0]),
.flogtanh( I688e5b6520508178afdf85bb2194186d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie96ab4759efe3dc122ef44bfc6a90d57  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I688e5b6520508178afdf85bb2194186d };
assign I0f6cb7a5a31d6f2f6178632c0c898bc6 = (If1f732841adb7c0cad1ba37c0f5fd517[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie96ab4759efe3dc122ef44bfc6a90d57;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00019_U (
.flogtanh_sel( I0df8a24f31c027756d248c3bd1b9bf7b[flogtanh_SEL-1:0]),
.flogtanh( I658630f3cf0e86ea86c5fb78b025b0a5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I04dc248d1a638da8d295d8061c0c05af  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I658630f3cf0e86ea86c5fb78b025b0a5 };
assign I03bea609a189246a2375b355df47cf81 = (I0df8a24f31c027756d248c3bd1b9bf7b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I04dc248d1a638da8d295d8061c0c05af;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00020_U (
.flogtanh_sel( I8ef901e733b12e76412eb36684e2b575[flogtanh_SEL-1:0]),
.flogtanh( I8b17f8bae259d829b52aba173bf10b4f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1260e022c28d8a62d5d93d3d79ddb362  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8b17f8bae259d829b52aba173bf10b4f };
assign If56555b7cf539750706cf678030ccdb2 = (I8ef901e733b12e76412eb36684e2b575[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1260e022c28d8a62d5d93d3d79ddb362;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00000_00021_U (
.flogtanh_sel( Ia48916a02f68b1b8f5fc7fece04677bb[flogtanh_SEL-1:0]),
.flogtanh( I944da8181119550916eaf431c7b04c50),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic77c9c3db51f43825807763f215fd048  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I944da8181119550916eaf431c7b04c50 };
assign I94e89b3a841f9760e3967c97e86d7160 = (Ia48916a02f68b1b8f5fc7fece04677bb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic77c9c3db51f43825807763f215fd048;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00000_U (
.flogtanh_sel( Ia37409944d9fdd3b16e7007e13d82a79[flogtanh_SEL-1:0]),
.flogtanh( I3aa615fa11ad382432ca658ec233f094),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ied24350a62d144813a9469693b4ebdf9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3aa615fa11ad382432ca658ec233f094 };
assign I8cab6f6faf0758f26d1a8851fae43896 = (Ia37409944d9fdd3b16e7007e13d82a79[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ied24350a62d144813a9469693b4ebdf9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00001_U (
.flogtanh_sel( Idd65f149afe9d5f63ddaf34b82b11e95[flogtanh_SEL-1:0]),
.flogtanh( Ib7c4f77c160ec436e93ca9de75b9fe42),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I167e15d8d78007dec518f69156f35a5a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib7c4f77c160ec436e93ca9de75b9fe42 };
assign I6ecf7249e6151477fe74a79d0b126b21 = (Idd65f149afe9d5f63ddaf34b82b11e95[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I167e15d8d78007dec518f69156f35a5a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00002_U (
.flogtanh_sel( If2886d560854faed32ebd8e33d868973[flogtanh_SEL-1:0]),
.flogtanh( Ic1e06942b276ee0933dc8b85dec58756),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If253f429b0dfc533c619ae813c74142b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic1e06942b276ee0933dc8b85dec58756 };
assign I3753b2c4ba8f1bee70def390a96586b0 = (If2886d560854faed32ebd8e33d868973[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If253f429b0dfc533c619ae813c74142b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00003_U (
.flogtanh_sel( I77778118bb3ea900c080754ff4c49c26[flogtanh_SEL-1:0]),
.flogtanh( Idd96d8b4e7be386203ec3ed3a81391d9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2921abdedb74a12af95c937ddaa1b8f4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idd96d8b4e7be386203ec3ed3a81391d9 };
assign I9b919f3d4ee3f33506b87bcdaf2d43a3 = (I77778118bb3ea900c080754ff4c49c26[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2921abdedb74a12af95c937ddaa1b8f4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00004_U (
.flogtanh_sel( I7292ed752d8741594d757730950feea4[flogtanh_SEL-1:0]),
.flogtanh( I7df43eec4d78baa1e0680be2715c4495),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia79f124f8610ca14d7c94a6bcbae2fbc  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7df43eec4d78baa1e0680be2715c4495 };
assign Ib3be128b6704cc04c61e0fc9814dcf20 = (I7292ed752d8741594d757730950feea4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia79f124f8610ca14d7c94a6bcbae2fbc;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00005_U (
.flogtanh_sel( I68cfd7868e061793ee8a41e69e80219b[flogtanh_SEL-1:0]),
.flogtanh( Ief08536c38479e6bc7fe786cfaf9a10f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3eb57d0d824ddfa6c789f4bee8a31bc9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ief08536c38479e6bc7fe786cfaf9a10f };
assign If365a3c3ef86dca7c7315b91298c2db8 = (I68cfd7868e061793ee8a41e69e80219b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3eb57d0d824ddfa6c789f4bee8a31bc9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00006_U (
.flogtanh_sel( I667ead814b303fca64ef047bb8246b19[flogtanh_SEL-1:0]),
.flogtanh( I6ef440b2077563ebbe50dde593c3875a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic6b78f30df38e245b28bc68cf70c2ae7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6ef440b2077563ebbe50dde593c3875a };
assign I83560e8d0f8cd37815cca6336fb2208d = (I667ead814b303fca64ef047bb8246b19[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic6b78f30df38e245b28bc68cf70c2ae7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00007_U (
.flogtanh_sel( I4f25c7edb12e868cb5532e42b4ba5133[flogtanh_SEL-1:0]),
.flogtanh( I20cfad172f0a614687d72d2337ef1003),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I68c4a1f713673e5cfd7d40fa2bafb2ec  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I20cfad172f0a614687d72d2337ef1003 };
assign I099441ae3d3dffe49b18bc578af54dc7 = (I4f25c7edb12e868cb5532e42b4ba5133[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I68c4a1f713673e5cfd7d40fa2bafb2ec;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00008_U (
.flogtanh_sel( I5aed2d82717f359bb5ac5a0ab91b7beb[flogtanh_SEL-1:0]),
.flogtanh( Icc6a92285959b25d53b452aed0718c8e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I740a82b22b7a0952639a5d85216e21a3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icc6a92285959b25d53b452aed0718c8e };
assign I58f89947eead94b5054a0fea3520ae33 = (I5aed2d82717f359bb5ac5a0ab91b7beb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I740a82b22b7a0952639a5d85216e21a3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00009_U (
.flogtanh_sel( I92835fd54631deaefa7b214e2c4b9bff[flogtanh_SEL-1:0]),
.flogtanh( I132c12f1eafbe34bca7b070354bd5f43),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I09eae10c74bf18420f829c7f7370e37f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I132c12f1eafbe34bca7b070354bd5f43 };
assign Ibf565bf1803ed43120fa54b80f6f1f29 = (I92835fd54631deaefa7b214e2c4b9bff[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I09eae10c74bf18420f829c7f7370e37f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00010_U (
.flogtanh_sel( I67e067da565635fcff166e3a7d0c446b[flogtanh_SEL-1:0]),
.flogtanh( I0f327225758bc82a67a65b8714949a91),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I939101803b39bb81310da5f0e6c4a0cb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0f327225758bc82a67a65b8714949a91 };
assign I619957528c630e7f64924a25127c93fb = (I67e067da565635fcff166e3a7d0c446b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I939101803b39bb81310da5f0e6c4a0cb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00011_U (
.flogtanh_sel( Ifdb0f307b1b9458c0487a1574ccc094b[flogtanh_SEL-1:0]),
.flogtanh( Ia90d4bc44d3687e912b59e4b6ca02718),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifea9a62f7fd17b6084afeb9d8ea50e91  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia90d4bc44d3687e912b59e4b6ca02718 };
assign If3cc31fd16469339470702045fc6d0da = (Ifdb0f307b1b9458c0487a1574ccc094b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifea9a62f7fd17b6084afeb9d8ea50e91;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00012_U (
.flogtanh_sel( I5c6b7d143e42fd3b8bcdb7d7ed4da2c2[flogtanh_SEL-1:0]),
.flogtanh( I21c1757545cc2732445c7f978f7247c4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1b740d99a82724a4bf44d320c0327ad9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I21c1757545cc2732445c7f978f7247c4 };
assign I338ccc17dc6158aec0129c8b0c02c429 = (I5c6b7d143e42fd3b8bcdb7d7ed4da2c2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1b740d99a82724a4bf44d320c0327ad9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00013_U (
.flogtanh_sel( Ie679a21d0136a08cc5e6526e9f8d1843[flogtanh_SEL-1:0]),
.flogtanh( I096fb1aff9431ed667e5d85a6f3726a4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2f8f6138bbd0bde03c51eafca516e891  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I096fb1aff9431ed667e5d85a6f3726a4 };
assign I83d71a89f35eb73265ee3e54184e1277 = (Ie679a21d0136a08cc5e6526e9f8d1843[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2f8f6138bbd0bde03c51eafca516e891;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00014_U (
.flogtanh_sel( I611942a72a5e12f6afaea6bde6699ef6[flogtanh_SEL-1:0]),
.flogtanh( Ia69d80cc1f2957ccd79cbd466dea987e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I685c70ac0a2f3404b34c778e92ed5cc7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia69d80cc1f2957ccd79cbd466dea987e };
assign I7362f08ed4e4ae309dfbfda112c56ad6 = (I611942a72a5e12f6afaea6bde6699ef6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I685c70ac0a2f3404b34c778e92ed5cc7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00015_U (
.flogtanh_sel( Ica9883c97f823a4491cbee5b45c43590[flogtanh_SEL-1:0]),
.flogtanh( I2243822bb5cdbca7f2ea942c7b720da8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I759d865a49afde724f226924f73a05eb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2243822bb5cdbca7f2ea942c7b720da8 };
assign I8be4be8471625db0749e6385f87d2dcc = (Ica9883c97f823a4491cbee5b45c43590[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I759d865a49afde724f226924f73a05eb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00016_U (
.flogtanh_sel( I8e6addfc61f5bfb7af74fc2993639565[flogtanh_SEL-1:0]),
.flogtanh( Ia77953e90a0cb40984d138c2c209db01),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1917af731dc6b46486e61cf077527e99  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia77953e90a0cb40984d138c2c209db01 };
assign I3d6a685a1913bd8be01fddbce1edec2e = (I8e6addfc61f5bfb7af74fc2993639565[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1917af731dc6b46486e61cf077527e99;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00017_U (
.flogtanh_sel( I9d53619f10e2a426f7297bbf7c81158a[flogtanh_SEL-1:0]),
.flogtanh( Id0b03e6dafabbe570f2626f51c9b7121),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3a0a357e2a3b16010a236fa1390680bb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id0b03e6dafabbe570f2626f51c9b7121 };
assign Ifd77e040c5f82790b1d5636a42fca602 = (I9d53619f10e2a426f7297bbf7c81158a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3a0a357e2a3b16010a236fa1390680bb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00018_U (
.flogtanh_sel( I8a055c27778913287ad951183fa0d4d6[flogtanh_SEL-1:0]),
.flogtanh( I5bfac7858439b218179c95c8d8669f17),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8fc051eb8bedd8d14a81345e7f7914c1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5bfac7858439b218179c95c8d8669f17 };
assign Ifbe479e5cab3cba43444bec1e12e72a0 = (I8a055c27778913287ad951183fa0d4d6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8fc051eb8bedd8d14a81345e7f7914c1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00019_U (
.flogtanh_sel( I8f6ae5c80bb2f50084b5f5ee5ab0ffc3[flogtanh_SEL-1:0]),
.flogtanh( I52497c500164c2417f928196ddcdbf84),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9fb6f6ed170f2e914c07ca1973723f74  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I52497c500164c2417f928196ddcdbf84 };
assign Ia784f35a5a46837b69eb048dabf84052 = (I8f6ae5c80bb2f50084b5f5ee5ab0ffc3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9fb6f6ed170f2e914c07ca1973723f74;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00020_U (
.flogtanh_sel( I3db8b3a342e8e2f13a448246aa001c2f[flogtanh_SEL-1:0]),
.flogtanh( Ib499dd504da7e433bc1caa258d7e7101),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib061c8e0e8a973cd42a1861b6f27af43  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib499dd504da7e433bc1caa258d7e7101 };
assign I8d0f440df332ea96e2d56eec490fbd51 = (I3db8b3a342e8e2f13a448246aa001c2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib061c8e0e8a973cd42a1861b6f27af43;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00001_00021_U (
.flogtanh_sel( Ibbee0996ea0f5e16b1f711345be7f2ae[flogtanh_SEL-1:0]),
.flogtanh( I7af88e2be096e488d7269479f935d185),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If746d7ebe9868d7bdf6b1884d933fbf8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7af88e2be096e488d7269479f935d185 };
assign I8d431a0524241fa54cf6dd1e79de4c74 = (Ibbee0996ea0f5e16b1f711345be7f2ae[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If746d7ebe9868d7bdf6b1884d933fbf8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00000_U (
.flogtanh_sel( Idb777f1eb4c3cbba103b9b43f948ccf9[flogtanh_SEL-1:0]),
.flogtanh( Ief51cc849e0034a9a6b3ff061064ad64),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4c999268e31b807c7ebf1fcb6d0e92e0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ief51cc849e0034a9a6b3ff061064ad64 };
assign If49f97cc0c42b23ce393b534015559a0 = (Idb777f1eb4c3cbba103b9b43f948ccf9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4c999268e31b807c7ebf1fcb6d0e92e0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00001_U (
.flogtanh_sel( Id5e46b1f8844c7587f99d22170581a24[flogtanh_SEL-1:0]),
.flogtanh( Ic5f096a42ae6fec933dcaf85faeeda49),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If3b89280e3fb4b1526d886740bfcafa4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic5f096a42ae6fec933dcaf85faeeda49 };
assign Ie932a22a7f1fa37087cbc9e8d73efef4 = (Id5e46b1f8844c7587f99d22170581a24[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If3b89280e3fb4b1526d886740bfcafa4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00002_U (
.flogtanh_sel( I67aadabd3cf49456cace7392a1e7a35a[flogtanh_SEL-1:0]),
.flogtanh( Ic9c0a2ce51d641ba7896c2c6911d0f96),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I608cd3a092bac42c3f31cea0545ba5b1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic9c0a2ce51d641ba7896c2c6911d0f96 };
assign I2956687a5fc2fba7149889624ef85647 = (I67aadabd3cf49456cace7392a1e7a35a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I608cd3a092bac42c3f31cea0545ba5b1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00003_U (
.flogtanh_sel( Id5635595d6b7b6dd7e6d510a27ad6702[flogtanh_SEL-1:0]),
.flogtanh( Ia96b3ea2e8395671b3ac674f5a956771),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6c65ea90fb08a2fc85cd61ef7db74ad1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia96b3ea2e8395671b3ac674f5a956771 };
assign Iebf28886bd39c2540c90e808a9c20d3d = (Id5635595d6b7b6dd7e6d510a27ad6702[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6c65ea90fb08a2fc85cd61ef7db74ad1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00004_U (
.flogtanh_sel( Ice783314a4868f0bba8bc3c5e3b65ae4[flogtanh_SEL-1:0]),
.flogtanh( Ib81d241e073c97c8c8d1d0abd9a9a64f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iac77fb31885852fa8f837806ffc0f7b5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib81d241e073c97c8c8d1d0abd9a9a64f };
assign I8d4f3e64c8e3b0710a4a6b30d27c8be8 = (Ice783314a4868f0bba8bc3c5e3b65ae4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iac77fb31885852fa8f837806ffc0f7b5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00005_U (
.flogtanh_sel( Ib2d9b7f58cf571b904be02e6073f9b94[flogtanh_SEL-1:0]),
.flogtanh( I0fc5e49719d7132c7724ee0d406ff93e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9b000348cc0f46026065aa4af2e5411c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0fc5e49719d7132c7724ee0d406ff93e };
assign I16e3f3a6802fd206654bb622fa1393fe = (Ib2d9b7f58cf571b904be02e6073f9b94[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9b000348cc0f46026065aa4af2e5411c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00006_U (
.flogtanh_sel( I61b6effae91ae4bdcce4550eb5cf0796[flogtanh_SEL-1:0]),
.flogtanh( I4479a0c26d4fa67dee328ecae12d14a4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9ed46b5dfd0052a65799266c17e3a6e2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4479a0c26d4fa67dee328ecae12d14a4 };
assign I4b5713aee09999592256c407d4b8a95a = (I61b6effae91ae4bdcce4550eb5cf0796[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9ed46b5dfd0052a65799266c17e3a6e2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00007_U (
.flogtanh_sel( If5cf6e81b0e3b77f6a45f2555201acc2[flogtanh_SEL-1:0]),
.flogtanh( If5693e079544d04478ec3da9a0ba28d7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie1cc391df396e85d4eb86799697a10f5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If5693e079544d04478ec3da9a0ba28d7 };
assign Ieb1dbb98d5e5bda5b9ce803857f2ca26 = (If5cf6e81b0e3b77f6a45f2555201acc2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie1cc391df396e85d4eb86799697a10f5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00008_U (
.flogtanh_sel( I62fae5bf51588f28c3521715b834909d[flogtanh_SEL-1:0]),
.flogtanh( I701a0ec899c88feef97aeb45fe19e639),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4d60c396c543011e7df7eeb9c9a97137  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I701a0ec899c88feef97aeb45fe19e639 };
assign Ife1c8d014675240a94f1133a78703ed5 = (I62fae5bf51588f28c3521715b834909d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4d60c396c543011e7df7eeb9c9a97137;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00009_U (
.flogtanh_sel( If5cbdab78a4cf86b6285a400d0e0ac90[flogtanh_SEL-1:0]),
.flogtanh( I6e9d61b111a45e4ea92ff12d33801755),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2ceb0debcadefafcbf0243be5f88f1a0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6e9d61b111a45e4ea92ff12d33801755 };
assign I94d9412a7b43fa0bd4b9a6d32d313fc7 = (If5cbdab78a4cf86b6285a400d0e0ac90[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2ceb0debcadefafcbf0243be5f88f1a0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00010_U (
.flogtanh_sel( I6e481cc49441c08bcd9fdcabbe90a000[flogtanh_SEL-1:0]),
.flogtanh( Ief65b0dab6ce1c2fc23cd297a21ac8de),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieeb8646e8e988cd3e9af56d6aeb23bc1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ief65b0dab6ce1c2fc23cd297a21ac8de };
assign If13e359e530823319046ce20027445dd = (I6e481cc49441c08bcd9fdcabbe90a000[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieeb8646e8e988cd3e9af56d6aeb23bc1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00011_U (
.flogtanh_sel( I3aa663be3dd604564ef68b9a2b9d7319[flogtanh_SEL-1:0]),
.flogtanh( Ibb843c4198a06c8e46bc954663c52a28),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibcadabc2f0ee0f0666a36571bf34a329  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibb843c4198a06c8e46bc954663c52a28 };
assign I221777352b48c4e228c6637410113854 = (I3aa663be3dd604564ef68b9a2b9d7319[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibcadabc2f0ee0f0666a36571bf34a329;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00012_U (
.flogtanh_sel( I8031632ee8700c63c207e2d6a6bdb630[flogtanh_SEL-1:0]),
.flogtanh( I0c043ef5daa388e93fb3cf6465c217b5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic762049ed90ead4c601316c55b05f9fc  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0c043ef5daa388e93fb3cf6465c217b5 };
assign I1ee46fec2b82cf8e5142f8e2ac5d9d8a = (I8031632ee8700c63c207e2d6a6bdb630[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic762049ed90ead4c601316c55b05f9fc;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00013_U (
.flogtanh_sel( If9be2701858da0bdffbf2dff7bcfd7e1[flogtanh_SEL-1:0]),
.flogtanh( Ife3f07ad3ad5228f10da7020a01e7069),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8c490934df0e2ca56338854686dec05d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ife3f07ad3ad5228f10da7020a01e7069 };
assign Ie45aaf966aa0a94803050b5f43d69e6c = (If9be2701858da0bdffbf2dff7bcfd7e1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8c490934df0e2ca56338854686dec05d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00014_U (
.flogtanh_sel( Ief209532f4cbf1c6a41bea414577f825[flogtanh_SEL-1:0]),
.flogtanh( I2dacd37cecd93c6e9134cb55ed917d78),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I16d19d1f42cf6f0bb1a4f67256aa2d75  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2dacd37cecd93c6e9134cb55ed917d78 };
assign I88aedd7f52399f5fd435c3415f2218ca = (Ief209532f4cbf1c6a41bea414577f825[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I16d19d1f42cf6f0bb1a4f67256aa2d75;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00015_U (
.flogtanh_sel( I1c8953ad3f64f3c3cc506808aad29dab[flogtanh_SEL-1:0]),
.flogtanh( I2419bc316181acd41e29ad005241d812),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5f703ca84e25e921f2d39aae0e1ce236  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2419bc316181acd41e29ad005241d812 };
assign I7651176b0a74846108fbaabc5cc4900a = (I1c8953ad3f64f3c3cc506808aad29dab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5f703ca84e25e921f2d39aae0e1ce236;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00016_U (
.flogtanh_sel( I1b519d88bbf86cfb080a50ea0480a128[flogtanh_SEL-1:0]),
.flogtanh( I35faf0af91f4972ae843883993fc84f4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib9de52ec38d9894c339f0d2222da3392  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I35faf0af91f4972ae843883993fc84f4 };
assign I57ac487adc18165136e9b3c7c50f95ad = (I1b519d88bbf86cfb080a50ea0480a128[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib9de52ec38d9894c339f0d2222da3392;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00017_U (
.flogtanh_sel( I5b8258f35d889071109216b464abb2a4[flogtanh_SEL-1:0]),
.flogtanh( I4dd2e7b6a685958d7aac77a38354e05f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ida9dc9ab7922a658c11f40e95543380e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4dd2e7b6a685958d7aac77a38354e05f };
assign Ic95668328a2121027436f682bac50b9c = (I5b8258f35d889071109216b464abb2a4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ida9dc9ab7922a658c11f40e95543380e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00018_U (
.flogtanh_sel( Id9681d4e0e4d375f9279de115a4337a3[flogtanh_SEL-1:0]),
.flogtanh( Ib27460a2e2b13abc54f5ba37f32c8653),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I37405a9f44d2155c4e3ecbb317d4b460  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib27460a2e2b13abc54f5ba37f32c8653 };
assign I118726375ca9381e45f001965fcefc5b = (Id9681d4e0e4d375f9279de115a4337a3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I37405a9f44d2155c4e3ecbb317d4b460;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00019_U (
.flogtanh_sel( Ib42144ece00b82debd70011724a29c91[flogtanh_SEL-1:0]),
.flogtanh( Ia3fa91387788798672eb6199a2eaa389),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I47527b41185c39cf18b85e38e3b870de  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia3fa91387788798672eb6199a2eaa389 };
assign Ic8d47ff5d6c31601a57df868da78c2d4 = (Ib42144ece00b82debd70011724a29c91[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I47527b41185c39cf18b85e38e3b870de;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00020_U (
.flogtanh_sel( Ic5717058a1815f63f164de1b1defe8cb[flogtanh_SEL-1:0]),
.flogtanh( Ieecd194ccc5698a2ba16efd969cfd621),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I995e084dd500652af249f8362d318a97  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ieecd194ccc5698a2ba16efd969cfd621 };
assign I7cdc5ada6fc68ee31fd4062e2ff004d3 = (Ic5717058a1815f63f164de1b1defe8cb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I995e084dd500652af249f8362d318a97;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00002_00021_U (
.flogtanh_sel( Iea41672f012f225d64d9c75b198c812f[flogtanh_SEL-1:0]),
.flogtanh( Ifb09fa1840c5a1ddbfc81cda21c11f1e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id844e291780b20b6e8fd26f9e45fa605  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifb09fa1840c5a1ddbfc81cda21c11f1e };
assign I59547aacdcfde31dc016ec2acbb2f4b4 = (Iea41672f012f225d64d9c75b198c812f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id844e291780b20b6e8fd26f9e45fa605;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00000_U (
.flogtanh_sel( I7a070bd014e1d2c5e55e5fcba88a5664[flogtanh_SEL-1:0]),
.flogtanh( I4ce505ae2025bab3abcf5a44e0ed5034),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If47a892c09147f3013077bf8ecf88619  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4ce505ae2025bab3abcf5a44e0ed5034 };
assign Ia7f53f0cd86055da72c13ac474f052a1 = (I7a070bd014e1d2c5e55e5fcba88a5664[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If47a892c09147f3013077bf8ecf88619;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00001_U (
.flogtanh_sel( I4a0a8b28429b708363458c74230b0fc2[flogtanh_SEL-1:0]),
.flogtanh( Id40a7ca1cde7a70cc13e752e19132808),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I41d2ac3db0c604f72f048017b3e8c5cb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id40a7ca1cde7a70cc13e752e19132808 };
assign I915054f2fbb8b93516d8748a3e3e29e2 = (I4a0a8b28429b708363458c74230b0fc2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I41d2ac3db0c604f72f048017b3e8c5cb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00002_U (
.flogtanh_sel( If585e4075ac1740f3b141ae6a50200f7[flogtanh_SEL-1:0]),
.flogtanh( If7274be2bcc8b2a235c3538db5506d90),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9a54d4d4c2c34cc7807874b016d7c4e2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If7274be2bcc8b2a235c3538db5506d90 };
assign If257757fa31c2f4cc9ec322e4ecccf83 = (If585e4075ac1740f3b141ae6a50200f7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9a54d4d4c2c34cc7807874b016d7c4e2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00003_U (
.flogtanh_sel( Ie1a68cf09bb21a1629369fde87f51bea[flogtanh_SEL-1:0]),
.flogtanh( I3e611982ec9ff6437f22e11b2552693a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ica6b595e3f7d1227e3e90d111d4d7585  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3e611982ec9ff6437f22e11b2552693a };
assign If91268e2b84df18785cd6a53e53eb4e9 = (Ie1a68cf09bb21a1629369fde87f51bea[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ica6b595e3f7d1227e3e90d111d4d7585;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00004_U (
.flogtanh_sel( I72b8547125d0ad6c1ad39a68b55c818c[flogtanh_SEL-1:0]),
.flogtanh( I8fcf0a468234f365c33059e26b9f5821),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icb87e0bd4997398dfb11b851e85e5d50  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8fcf0a468234f365c33059e26b9f5821 };
assign Ia072f1d679429d3c3180f8eb67fc7dd7 = (I72b8547125d0ad6c1ad39a68b55c818c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icb87e0bd4997398dfb11b851e85e5d50;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00005_U (
.flogtanh_sel( Ie14ba4a8657740f9a8d057258db2cb09[flogtanh_SEL-1:0]),
.flogtanh( I3f80250ee19e8250898f2bcc055c2e5b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia1d6b8a34f2f4b6b3495ae760183f9b3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3f80250ee19e8250898f2bcc055c2e5b };
assign I91a8168d3b087ab3891cd6d479427b95 = (Ie14ba4a8657740f9a8d057258db2cb09[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia1d6b8a34f2f4b6b3495ae760183f9b3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00006_U (
.flogtanh_sel( I27490a69fb2a1f6f298639254c37cf9e[flogtanh_SEL-1:0]),
.flogtanh( I06b3652935db14aaa057f0cf3cffef66),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib74566da453368c9846342fdeafcee15  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I06b3652935db14aaa057f0cf3cffef66 };
assign Id1dce8c1542f1279badb381aca3c9b51 = (I27490a69fb2a1f6f298639254c37cf9e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib74566da453368c9846342fdeafcee15;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00007_U (
.flogtanh_sel( I49b9c212fbe74a5dd8b087e417296186[flogtanh_SEL-1:0]),
.flogtanh( Ib01d30e88a3a1fcb204246baafeb47c8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If2cfb11905db55514942ab73b9db82aa  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib01d30e88a3a1fcb204246baafeb47c8 };
assign I8983f003c30a218543f39f5bbcd9a25c = (I49b9c212fbe74a5dd8b087e417296186[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If2cfb11905db55514942ab73b9db82aa;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00008_U (
.flogtanh_sel( I0a8e6f5cc8b6ea599b7605abe6479bec[flogtanh_SEL-1:0]),
.flogtanh( I9f688c58878405d1d2865ddc40659c2b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I60da6c145c6e2723bf4ff550f857a977  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9f688c58878405d1d2865ddc40659c2b };
assign Id1b5c33bc63f75561b7cce6fc0981c69 = (I0a8e6f5cc8b6ea599b7605abe6479bec[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I60da6c145c6e2723bf4ff550f857a977;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00009_U (
.flogtanh_sel( Ib6d94b34d3886717e4016fec196f277f[flogtanh_SEL-1:0]),
.flogtanh( Ic9c77123914f831cee5bc4586b6a2a8b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0f3219717265b7d82d487dea1a63cb62  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic9c77123914f831cee5bc4586b6a2a8b };
assign I003f95fb8f2027efa41a1936e8b53986 = (Ib6d94b34d3886717e4016fec196f277f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0f3219717265b7d82d487dea1a63cb62;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00010_U (
.flogtanh_sel( Id7e53d36da7171e036ebfc984dbcea6e[flogtanh_SEL-1:0]),
.flogtanh( Ifd42760504e0f106eb9061d9b9a2d18a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9a4db851c1d6935ab3dfdae9fb85680e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifd42760504e0f106eb9061d9b9a2d18a };
assign Ie16dc913f571ae73ce03d755077345a9 = (Id7e53d36da7171e036ebfc984dbcea6e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9a4db851c1d6935ab3dfdae9fb85680e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00011_U (
.flogtanh_sel( I2ec254d80fd0683d782302cf3839559b[flogtanh_SEL-1:0]),
.flogtanh( I452794105cca79653f5509dac3794327),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I00b3675542777a857263214ae2fa08cd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I452794105cca79653f5509dac3794327 };
assign I86e53eed5b857c439039238bb486067c = (I2ec254d80fd0683d782302cf3839559b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I00b3675542777a857263214ae2fa08cd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00012_U (
.flogtanh_sel( Ibbedaef61051d5df82cd6d55e05c80da[flogtanh_SEL-1:0]),
.flogtanh( I33431ed9c549f5525adfa5d45fbc7653),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I695c8725ab88beb04f4eeb9d1ec5cbab  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I33431ed9c549f5525adfa5d45fbc7653 };
assign I89433799cfa534afd66e8d6b9f1b62b9 = (Ibbedaef61051d5df82cd6d55e05c80da[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I695c8725ab88beb04f4eeb9d1ec5cbab;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00013_U (
.flogtanh_sel( I501336bb7ba172c05dd5840036e6228c[flogtanh_SEL-1:0]),
.flogtanh( I4b8b4fd334b176cb449ad0296ebff4c8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3317b620629d4ed1162708dd76c7fea0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4b8b4fd334b176cb449ad0296ebff4c8 };
assign I80f2e8f6743e28e86e4d85b295e2f768 = (I501336bb7ba172c05dd5840036e6228c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3317b620629d4ed1162708dd76c7fea0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00014_U (
.flogtanh_sel( I8e5c4c6c63e42054359cee697cc0d026[flogtanh_SEL-1:0]),
.flogtanh( I66e7dacba9dbfb14e9a71b9d57229880),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I13a81876edd15dc11e22d573b5a33e83  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I66e7dacba9dbfb14e9a71b9d57229880 };
assign I1391018fb93372ccc2fcc08700e38b65 = (I8e5c4c6c63e42054359cee697cc0d026[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I13a81876edd15dc11e22d573b5a33e83;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00015_U (
.flogtanh_sel( Id3daa6db921871b752bf92366446afcc[flogtanh_SEL-1:0]),
.flogtanh( If3a842c52c8c0b2fd24ef265e8cfe330),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I64528d9704c63c85bdf41fb3bd66587d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If3a842c52c8c0b2fd24ef265e8cfe330 };
assign I8fd26d47ecd4cdd08294cf6133468d17 = (Id3daa6db921871b752bf92366446afcc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I64528d9704c63c85bdf41fb3bd66587d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00016_U (
.flogtanh_sel( Id8367ec60787bfad0da8aa76c6ed8ddb[flogtanh_SEL-1:0]),
.flogtanh( I0f3aea4265966e7bc673d3a08ad1c2e4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I38228bcb39eb9ea57aa0bd811e6976a2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0f3aea4265966e7bc673d3a08ad1c2e4 };
assign I7097c9518bb3351818b96f31ed49c6d3 = (Id8367ec60787bfad0da8aa76c6ed8ddb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I38228bcb39eb9ea57aa0bd811e6976a2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00017_U (
.flogtanh_sel( I533649312ec995f1f9e514c59a8675b1[flogtanh_SEL-1:0]),
.flogtanh( Ia9de78211d220e68835ff757eb75d919),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6ddd4fd20c147c6dff337057753a4ec2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia9de78211d220e68835ff757eb75d919 };
assign Id683d693cd50645c3d6d657aa1c8bdb2 = (I533649312ec995f1f9e514c59a8675b1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6ddd4fd20c147c6dff337057753a4ec2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00018_U (
.flogtanh_sel( I0621d0b2c83e70b4afd65eb9dca4b514[flogtanh_SEL-1:0]),
.flogtanh( I2c1c31b8bda73b145cdf74b18bc46a4d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I73f34929e9a61c1a6b95107e277fb254  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2c1c31b8bda73b145cdf74b18bc46a4d };
assign I88bd8012c93dd9e2ed52ea5e9b8b0004 = (I0621d0b2c83e70b4afd65eb9dca4b514[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I73f34929e9a61c1a6b95107e277fb254;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00019_U (
.flogtanh_sel( I2ae01892a3cd0432618d7280b31daddb[flogtanh_SEL-1:0]),
.flogtanh( I300a84deada851e18835d6af55c5e2a3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib078dd08f08128d55534715ee61ea4b8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I300a84deada851e18835d6af55c5e2a3 };
assign Ia8d3667adc34b2b50acf7edb970538d8 = (I2ae01892a3cd0432618d7280b31daddb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib078dd08f08128d55534715ee61ea4b8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00020_U (
.flogtanh_sel( I5ed8a2f30bd2ea269341c2267ae3fe83[flogtanh_SEL-1:0]),
.flogtanh( I1fc6745ba86be641dc9bdac044c19519),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3f723dfd62f8ae0057a07480d74562db  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1fc6745ba86be641dc9bdac044c19519 };
assign I3f0bba472e912f11dea8e788fbc1cb63 = (I5ed8a2f30bd2ea269341c2267ae3fe83[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3f723dfd62f8ae0057a07480d74562db;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00003_00021_U (
.flogtanh_sel( I2c819e7f62c0dc0aac650074b203163b[flogtanh_SEL-1:0]),
.flogtanh( I2791cc5f69dd0e7f306760048c759af7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iff7040b14913e56cdf2b36168dcd751e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2791cc5f69dd0e7f306760048c759af7 };
assign I6dc671e73b4e9c70cabfdeaac2e5c40b = (I2c819e7f62c0dc0aac650074b203163b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iff7040b14913e56cdf2b36168dcd751e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00000_U (
.flogtanh_sel( I30e20b58913d6fbe5817e1956ba8e570[flogtanh_SEL-1:0]),
.flogtanh( Ie8157cde860052619820431f87e13c83),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I72540f5da4495184c7ae5ecc11a96939  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie8157cde860052619820431f87e13c83 };
assign Ia6255a136d5f36ea6cba654bd5823850 = (I30e20b58913d6fbe5817e1956ba8e570[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I72540f5da4495184c7ae5ecc11a96939;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00001_U (
.flogtanh_sel( I1b922bed7f3c4a6705f3ce7a885a68cd[flogtanh_SEL-1:0]),
.flogtanh( I9059b74a8f3cf2e4905756cc9c71597f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6174d9699747eed0b49d44974bfb21b0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9059b74a8f3cf2e4905756cc9c71597f };
assign I2b9584392ef9a7828ff57bd4c522a302 = (I1b922bed7f3c4a6705f3ce7a885a68cd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6174d9699747eed0b49d44974bfb21b0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00002_U (
.flogtanh_sel( I2f65f0917713ecc8585392d3b557c1bf[flogtanh_SEL-1:0]),
.flogtanh( I99584eabd3cbd2546c85f474afa6fabb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iadc74d3274cb3d595c39a8118b2410aa  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I99584eabd3cbd2546c85f474afa6fabb };
assign I6c1235e88ae444a96ea64fd1bfd04d8f = (I2f65f0917713ecc8585392d3b557c1bf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iadc74d3274cb3d595c39a8118b2410aa;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00003_U (
.flogtanh_sel( I3301533e7d9e527118a67c462f1b4357[flogtanh_SEL-1:0]),
.flogtanh( I047abade6abf10a65a5b835ac725fa7c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I27493e743da259f4886f63a08165560e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I047abade6abf10a65a5b835ac725fa7c };
assign Id09b8242c22851fb960d55222fe733d4 = (I3301533e7d9e527118a67c462f1b4357[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I27493e743da259f4886f63a08165560e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00004_U (
.flogtanh_sel( I52a88bdb1f03da82730f7579b7b5305d[flogtanh_SEL-1:0]),
.flogtanh( Icf7ab1d1113bc44358c56a56fca7caf9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I834b01b9c0bdcbe8cd616ab7dc5e2b91  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icf7ab1d1113bc44358c56a56fca7caf9 };
assign Ie355fa27abbc41291eaf08f2cf9a6ff7 = (I52a88bdb1f03da82730f7579b7b5305d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I834b01b9c0bdcbe8cd616ab7dc5e2b91;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00005_U (
.flogtanh_sel( I644c730662b3725d26cd46fb46106104[flogtanh_SEL-1:0]),
.flogtanh( I4d24650be7a1088c2310d93000d6392a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id69fd2756995da4325484ac912de043a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4d24650be7a1088c2310d93000d6392a };
assign I566224393f6bb27bfd8b0b0d6b8e53d6 = (I644c730662b3725d26cd46fb46106104[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id69fd2756995da4325484ac912de043a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00006_U (
.flogtanh_sel( I3da3e36c76c4123bec6879bccb39e933[flogtanh_SEL-1:0]),
.flogtanh( Ic3aea8ebb8eab44a92e7d7d950e1a917),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia23d77f7fcff89e09068364cf3de713a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic3aea8ebb8eab44a92e7d7d950e1a917 };
assign I8fcad6e7d5ffc9f79eaaf634f6fe8cda = (I3da3e36c76c4123bec6879bccb39e933[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia23d77f7fcff89e09068364cf3de713a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00007_U (
.flogtanh_sel( Iebde55cddc8170f7dd8855ea55eff0ce[flogtanh_SEL-1:0]),
.flogtanh( I82af0956870500474eac2505bbf15e35),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I781d4698facda706103ef8265810eaf6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I82af0956870500474eac2505bbf15e35 };
assign I6f0f74dcc830fdcb0af9df75a2b722f7 = (Iebde55cddc8170f7dd8855ea55eff0ce[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I781d4698facda706103ef8265810eaf6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00008_U (
.flogtanh_sel( Ie673e2d92a7090b2fa1c5e14a2e03be3[flogtanh_SEL-1:0]),
.flogtanh( I2d8a8efaa0179340bf5d3ebbd4c11831),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia92f18f2e26ec8ad3578f230d2201274  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2d8a8efaa0179340bf5d3ebbd4c11831 };
assign Idd95fd099dd2b53c46d02f09575b8032 = (Ie673e2d92a7090b2fa1c5e14a2e03be3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia92f18f2e26ec8ad3578f230d2201274;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00009_U (
.flogtanh_sel( If90afe75714f8660ad0eb9f9ea06cd6b[flogtanh_SEL-1:0]),
.flogtanh( I32ff895ff659ec448270067f76e97a90),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1b1a08cc28279b3ffdd544d38704c1ec  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I32ff895ff659ec448270067f76e97a90 };
assign I0f277bc88d46a4e6e9f1f2c410b503fd = (If90afe75714f8660ad0eb9f9ea06cd6b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1b1a08cc28279b3ffdd544d38704c1ec;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00010_U (
.flogtanh_sel( Ifd96e3a6e0050c30a4308328cfecb21f[flogtanh_SEL-1:0]),
.flogtanh( I15a7fd79aeb5eed24b1c7be3d48296e0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie12755a265f6a32154b88d22f2037962  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I15a7fd79aeb5eed24b1c7be3d48296e0 };
assign I66b92f1de2cf408c3af53b161a6ffa60 = (Ifd96e3a6e0050c30a4308328cfecb21f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie12755a265f6a32154b88d22f2037962;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00011_U (
.flogtanh_sel( I68b92cc2d83e9a718edd2aea82314016[flogtanh_SEL-1:0]),
.flogtanh( I12f311f2311e26320a178d6fec95d9d0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7c27744991b38f3eb69eb9ba2aeb0907  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I12f311f2311e26320a178d6fec95d9d0 };
assign Id28d9545e8d20ac080fbac5e345692da = (I68b92cc2d83e9a718edd2aea82314016[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7c27744991b38f3eb69eb9ba2aeb0907;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00012_U (
.flogtanh_sel( I6bdbb92363f0e072ed04654e9aad17a5[flogtanh_SEL-1:0]),
.flogtanh( I2b8ce30d1338ad506e4996d2dd1dc11a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0bbd6f8a9e1e7489421d3b744005b6e6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2b8ce30d1338ad506e4996d2dd1dc11a };
assign I4a5cfd6ebd47cda4fa2e06ba9ad6e5b2 = (I6bdbb92363f0e072ed04654e9aad17a5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0bbd6f8a9e1e7489421d3b744005b6e6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00013_U (
.flogtanh_sel( I87a4267db59b97ef1b9bca8743cb0322[flogtanh_SEL-1:0]),
.flogtanh( Ic2b65e7bd42e94f2ad8b6506a6fce7af),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib9f20533ee570afdeffb0f5279b51d9d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic2b65e7bd42e94f2ad8b6506a6fce7af };
assign I62bda8dc70e0b5eb38abe094bbe92fc6 = (I87a4267db59b97ef1b9bca8743cb0322[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib9f20533ee570afdeffb0f5279b51d9d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00014_U (
.flogtanh_sel( I44eacb2bea725efab7c0dd560279f0f8[flogtanh_SEL-1:0]),
.flogtanh( I0f54a697ea3e2bbf90354c9a6173fb80),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8edc9f2bff969700d0a7e735b533ee9f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0f54a697ea3e2bbf90354c9a6173fb80 };
assign I223b05d94c09b095d1988df121aa5e37 = (I44eacb2bea725efab7c0dd560279f0f8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8edc9f2bff969700d0a7e735b533ee9f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00015_U (
.flogtanh_sel( I87a2736466c5ee62b7cc55f17e715ffa[flogtanh_SEL-1:0]),
.flogtanh( I6a6c0f8e4399c21285d66ddc0f1f70c0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id97e6a4e20414f9a23afe284f3e492e3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6a6c0f8e4399c21285d66ddc0f1f70c0 };
assign I5f73e5faf1aca83ee0a415c9ac4a1b9a = (I87a2736466c5ee62b7cc55f17e715ffa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id97e6a4e20414f9a23afe284f3e492e3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00016_U (
.flogtanh_sel( I7a66c7713ba126fdc24940cd92f7e10b[flogtanh_SEL-1:0]),
.flogtanh( Ibfcdfc01f09bcff031e359394947efef),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If992b3a65059c6e5866c3a03828efb18  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibfcdfc01f09bcff031e359394947efef };
assign I75f9d3a41019dca3044a1c2cf7069662 = (I7a66c7713ba126fdc24940cd92f7e10b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If992b3a65059c6e5866c3a03828efb18;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00017_U (
.flogtanh_sel( I1f11c579f34c41aade41c53f53468057[flogtanh_SEL-1:0]),
.flogtanh( I8efd478f1ae2ea6090774e1ed3bd7b28),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie7448467fe54559f10316db6ad186b9e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8efd478f1ae2ea6090774e1ed3bd7b28 };
assign I820fa56328e3919970dd64adb1d4d8e7 = (I1f11c579f34c41aade41c53f53468057[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie7448467fe54559f10316db6ad186b9e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00018_U (
.flogtanh_sel( I651a438f70583d476ae10f066e035435[flogtanh_SEL-1:0]),
.flogtanh( I502d3210c60c82ca682d8e2168d54be0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3df80bf9e919f723f65f34362854119f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I502d3210c60c82ca682d8e2168d54be0 };
assign I05eadf11cdc6c2f2b021e33f2438fa49 = (I651a438f70583d476ae10f066e035435[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3df80bf9e919f723f65f34362854119f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00019_U (
.flogtanh_sel( Ibdf17fa73794c846e15fe0a915b071e5[flogtanh_SEL-1:0]),
.flogtanh( I337d74c3c773a358a936806f751c1117),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iefe3ca0afaed4b8f7d63ec54591c6cec  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I337d74c3c773a358a936806f751c1117 };
assign I2c487770d606451440eecf358202db32 = (Ibdf17fa73794c846e15fe0a915b071e5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iefe3ca0afaed4b8f7d63ec54591c6cec;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00020_U (
.flogtanh_sel( I76d3221fbcefc0ee08655f7ba4919f3c[flogtanh_SEL-1:0]),
.flogtanh( Ia494fdbd70bff11510eb685f3b5d0aae),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1614bb17d0c7c14b07ac4dde98c1fb2a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia494fdbd70bff11510eb685f3b5d0aae };
assign I082aa8c413d7ef8f054b1c2857cbe39f = (I76d3221fbcefc0ee08655f7ba4919f3c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1614bb17d0c7c14b07ac4dde98c1fb2a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00021_U (
.flogtanh_sel( I3458f69c90ea8b20b3d1f67e9a13ec2e[flogtanh_SEL-1:0]),
.flogtanh( I547f7a4c3801c1caa4587c9aef397652),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib1672ae7e0ce15c6fc9eeabc17b8ee97  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I547f7a4c3801c1caa4587c9aef397652 };
assign I420e2c5a8745133f6263a71b458f1e2f = (I3458f69c90ea8b20b3d1f67e9a13ec2e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib1672ae7e0ce15c6fc9eeabc17b8ee97;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00004_00022_U (
.flogtanh_sel( Ia2d6e9e1e92a30c7028af50ddfbb9bf9[flogtanh_SEL-1:0]),
.flogtanh( I8009d84fd826dd21eb7091744792f4a7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5efb28aa360b27578d1bbda19162507c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8009d84fd826dd21eb7091744792f4a7 };
assign I4b8d520ee88fd39d83a16432e962f731 = (Ia2d6e9e1e92a30c7028af50ddfbb9bf9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5efb28aa360b27578d1bbda19162507c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00000_U (
.flogtanh_sel( I66c91b5133d9812a03daecc0b14211f8[flogtanh_SEL-1:0]),
.flogtanh( If724b1c92350989910925d275353e544),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic661342fb3f026ac5b7ca0d5712f572c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If724b1c92350989910925d275353e544 };
assign Ia3f7f07ddb09ea33218afe14281ac3c6 = (I66c91b5133d9812a03daecc0b14211f8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic661342fb3f026ac5b7ca0d5712f572c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00001_U (
.flogtanh_sel( Ifb5986949e88167526d9fcfe07b417ca[flogtanh_SEL-1:0]),
.flogtanh( I26f4a180e992f5de04bc047f539bcb48),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I84437247e54c9c225c1441622ec111c4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I26f4a180e992f5de04bc047f539bcb48 };
assign I25aefb53f59a00abe88b9dcf6be6907a = (Ifb5986949e88167526d9fcfe07b417ca[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I84437247e54c9c225c1441622ec111c4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00002_U (
.flogtanh_sel( Iedada801ca6cd173ee523ef335e91ff6[flogtanh_SEL-1:0]),
.flogtanh( I83ca10d71caf5ac98fef3d45d228be8e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9e0295a7fa30f62feb64d3b4ed2dd4d2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I83ca10d71caf5ac98fef3d45d228be8e };
assign I22c3140a8db02352d2e2a2a11eeba117 = (Iedada801ca6cd173ee523ef335e91ff6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9e0295a7fa30f62feb64d3b4ed2dd4d2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00003_U (
.flogtanh_sel( I4e2722e547586da7565b2d91a7fc91e7[flogtanh_SEL-1:0]),
.flogtanh( Ib8407faa17d1e96cd317c65459c4fa71),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1042cc8af315aa7120ea813ae2c5755a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib8407faa17d1e96cd317c65459c4fa71 };
assign I954dd66f60316803a8f13a39c460a39a = (I4e2722e547586da7565b2d91a7fc91e7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1042cc8af315aa7120ea813ae2c5755a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00004_U (
.flogtanh_sel( Ib321a8ceda62c64ab25dc1c718301bda[flogtanh_SEL-1:0]),
.flogtanh( I73829d98e5e2f368c4a2020e3d7814be),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1f64264a2c913aeaf4db38f4190cd2dd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I73829d98e5e2f368c4a2020e3d7814be };
assign I37b3988d699a1ed42923e3fd1584ecc0 = (Ib321a8ceda62c64ab25dc1c718301bda[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1f64264a2c913aeaf4db38f4190cd2dd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00005_U (
.flogtanh_sel( I58daeebec4873e6c1c07c090ff81235c[flogtanh_SEL-1:0]),
.flogtanh( I9a120c441f8d9ccb617057e042587ba1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7fa463286e319877ffc9682e696aae89  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9a120c441f8d9ccb617057e042587ba1 };
assign If79bc5a35cb55036a367efb88c7d5510 = (I58daeebec4873e6c1c07c090ff81235c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7fa463286e319877ffc9682e696aae89;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00006_U (
.flogtanh_sel( I3f103fbbe49c86c9db46129bd4632cab[flogtanh_SEL-1:0]),
.flogtanh( I8064df8bc33998ad58d460afae699e48),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I59c12008dc705cc23fb3093f2ace7c38  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8064df8bc33998ad58d460afae699e48 };
assign Ideab06dc2448a6950cd1a06a0c90c2c6 = (I3f103fbbe49c86c9db46129bd4632cab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I59c12008dc705cc23fb3093f2ace7c38;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00007_U (
.flogtanh_sel( Id6697ca17f1bd6ddd112951b9d89a8ea[flogtanh_SEL-1:0]),
.flogtanh( If016e079d3b453444558706ef9073233),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I63f19ffd1e2bf12ea726afc806340062  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If016e079d3b453444558706ef9073233 };
assign I1d7d7a68fc53b8be89c4637ac8f29380 = (Id6697ca17f1bd6ddd112951b9d89a8ea[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I63f19ffd1e2bf12ea726afc806340062;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00008_U (
.flogtanh_sel( I445ede2983c7470b4418a2ec0cbbd5e1[flogtanh_SEL-1:0]),
.flogtanh( I51cc187d91ee3c480a759104aed41b1b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib5408f87beae3f337dfb1e8a75a42a19  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I51cc187d91ee3c480a759104aed41b1b };
assign Ib34ad1d14978608d1440f59998a31672 = (I445ede2983c7470b4418a2ec0cbbd5e1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib5408f87beae3f337dfb1e8a75a42a19;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00009_U (
.flogtanh_sel( I034e56cd77ee400ed81b78177b202930[flogtanh_SEL-1:0]),
.flogtanh( I4b8068a6a866c2424439b2956245ac8d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I71c3e022d15f1fb4f7b8ffc67c61ab90  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4b8068a6a866c2424439b2956245ac8d };
assign Id081512cd113e4d09df0fb13e443d76b = (I034e56cd77ee400ed81b78177b202930[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I71c3e022d15f1fb4f7b8ffc67c61ab90;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00010_U (
.flogtanh_sel( I08edadbd9366786f96b44268d096b4aa[flogtanh_SEL-1:0]),
.flogtanh( I60513d924016bd300559b7a1bea7f521),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifd815e691b57a5d6f200b40f3953327c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I60513d924016bd300559b7a1bea7f521 };
assign I57a0f8c3710cf8e216d6dc2420f7621c = (I08edadbd9366786f96b44268d096b4aa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifd815e691b57a5d6f200b40f3953327c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00011_U (
.flogtanh_sel( I8f86a7af86eb04c5df18e09888cdce7b[flogtanh_SEL-1:0]),
.flogtanh( Iec98284ab12724bb63360f29d00f1ecb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I507e631ff186c6a13a989e3bf09dfda0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iec98284ab12724bb63360f29d00f1ecb };
assign Iaa164a078c8cdaad694a053c9c1e0313 = (I8f86a7af86eb04c5df18e09888cdce7b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I507e631ff186c6a13a989e3bf09dfda0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00012_U (
.flogtanh_sel( Ic00d037a11f8a27ab34e4daab8c9c2e6[flogtanh_SEL-1:0]),
.flogtanh( I3e3eba8135eb797d0a5e8ac1feefce0c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7b0ca33814446a75f820ed3983b8f806  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3e3eba8135eb797d0a5e8ac1feefce0c };
assign I7eb76b3d17296fdae702d8f820f1428d = (Ic00d037a11f8a27ab34e4daab8c9c2e6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7b0ca33814446a75f820ed3983b8f806;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00013_U (
.flogtanh_sel( I4d95ceccc6c3ad37f13c98339c59e5c4[flogtanh_SEL-1:0]),
.flogtanh( I6aa98bc7265b8b7c25181a06e75c24c0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic0dd354cd8b9e5eb33fffc13285f00e9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6aa98bc7265b8b7c25181a06e75c24c0 };
assign I00ecb5e329390023b318a2ceba0df231 = (I4d95ceccc6c3ad37f13c98339c59e5c4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic0dd354cd8b9e5eb33fffc13285f00e9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00014_U (
.flogtanh_sel( I1ea967d377f462a0e06d7d0d4d95b342[flogtanh_SEL-1:0]),
.flogtanh( I47f9c7018999e1cea25feddbe399e6b7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifa81b0a7df922d4d85e99dec97ca6c9a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I47f9c7018999e1cea25feddbe399e6b7 };
assign Iea32ebc385c6cfc9212ff37973a0a05d = (I1ea967d377f462a0e06d7d0d4d95b342[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifa81b0a7df922d4d85e99dec97ca6c9a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00015_U (
.flogtanh_sel( Ib0feec63123e66bd6ad6935e9b7fa6bf[flogtanh_SEL-1:0]),
.flogtanh( I7224803ba8f0a16a7b2e969fe727bfa1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I91549d4c802e94f6b0400b459b1b5f50  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7224803ba8f0a16a7b2e969fe727bfa1 };
assign If845af0d620024f04525244753ba5d18 = (Ib0feec63123e66bd6ad6935e9b7fa6bf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I91549d4c802e94f6b0400b459b1b5f50;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00016_U (
.flogtanh_sel( I7d120060ddae9ff8f7206b3ef63eda50[flogtanh_SEL-1:0]),
.flogtanh( I65bc4e0d837f94c4301cb2c87e24969c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id002cb5fd3d0c0a5c0f7ab1ad6cef723  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I65bc4e0d837f94c4301cb2c87e24969c };
assign I08e907b0619bec3ef2cf4cb3779e0794 = (I7d120060ddae9ff8f7206b3ef63eda50[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id002cb5fd3d0c0a5c0f7ab1ad6cef723;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00017_U (
.flogtanh_sel( Ib47f8f72386e2e65a88fbadd3a705225[flogtanh_SEL-1:0]),
.flogtanh( I444f8e61602b8994f7a01f3ebd4ac6ab),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4c6a3ad23b392e26c465731aa152c61c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I444f8e61602b8994f7a01f3ebd4ac6ab };
assign I68e5b12792a86dda0576742831d3b728 = (Ib47f8f72386e2e65a88fbadd3a705225[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4c6a3ad23b392e26c465731aa152c61c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00018_U (
.flogtanh_sel( I4e0efc35346e2934f5bb4c34a4bc5f90[flogtanh_SEL-1:0]),
.flogtanh( I86c51ec7ff965132e195835d21c24881),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iebf49da6d6689a63afa17717ce18e786  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I86c51ec7ff965132e195835d21c24881 };
assign I72db05084d30d7c59ba1cb06d3b09400 = (I4e0efc35346e2934f5bb4c34a4bc5f90[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iebf49da6d6689a63afa17717ce18e786;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00019_U (
.flogtanh_sel( I3ca1014802f58087e3434a1e0df19c01[flogtanh_SEL-1:0]),
.flogtanh( I07aa1b2db5dedc3230dff10534311a56),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id2f4466e93345d0e36e5d72ab56c495c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I07aa1b2db5dedc3230dff10534311a56 };
assign Ib1f1aef6c0a9291553b62fd555feb2e7 = (I3ca1014802f58087e3434a1e0df19c01[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id2f4466e93345d0e36e5d72ab56c495c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00020_U (
.flogtanh_sel( I688a3879b7be1544e6f94b4221c03213[flogtanh_SEL-1:0]),
.flogtanh( Ia8809cc89c377e8b4109cdc8976daa54),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I804df90e3a9f73c97b372fc4ecf3dcac  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia8809cc89c377e8b4109cdc8976daa54 };
assign Ib504b808f724ca6032e7c746517cd4fd = (I688a3879b7be1544e6f94b4221c03213[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I804df90e3a9f73c97b372fc4ecf3dcac;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00021_U (
.flogtanh_sel( Ic22988138610c8671ec342f65f34c7ae[flogtanh_SEL-1:0]),
.flogtanh( I7402dc21bfbc0af749dd8fb03c516a50),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I52aa4e2bc75f024d35a92ae35bf1b627  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7402dc21bfbc0af749dd8fb03c516a50 };
assign Ia47f7fb27f2d965cfd2989569c257356 = (Ic22988138610c8671ec342f65f34c7ae[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I52aa4e2bc75f024d35a92ae35bf1b627;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00005_00022_U (
.flogtanh_sel( I0b85fdd83569e5cbb7d71eed50cb32fd[flogtanh_SEL-1:0]),
.flogtanh( I8ca06f4250a69dde75889f7a6ba3f456),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iefe341800d7dacd81be0ab984ab16f9f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8ca06f4250a69dde75889f7a6ba3f456 };
assign If2b17f9e9186542117f43d0dd342326e = (I0b85fdd83569e5cbb7d71eed50cb32fd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iefe341800d7dacd81be0ab984ab16f9f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00000_U (
.flogtanh_sel( Idf55390c11e5b41ebc2a28e0af109913[flogtanh_SEL-1:0]),
.flogtanh( Ibab00faeaa6a7be99fa6a239193b92cb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic8a0166e91618bc4c689d8b1cb063fdd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibab00faeaa6a7be99fa6a239193b92cb };
assign I6c4ba0863ab4c8d1a56324a4d89ccbeb = (Idf55390c11e5b41ebc2a28e0af109913[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic8a0166e91618bc4c689d8b1cb063fdd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00001_U (
.flogtanh_sel( I6b48935ea25672ee9a42f49eae9e519f[flogtanh_SEL-1:0]),
.flogtanh( I8e44b109466e00487db9dfb7ae225f89),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5097124bb6e421210e0884fcac4f151a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8e44b109466e00487db9dfb7ae225f89 };
assign I4dbd1bb8f1641f15e3a4f1e309962811 = (I6b48935ea25672ee9a42f49eae9e519f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5097124bb6e421210e0884fcac4f151a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00002_U (
.flogtanh_sel( I6a9e6c39c20e45773dab7823a7ff9486[flogtanh_SEL-1:0]),
.flogtanh( Ib3e38e46bfa9e1bdc032918269223b32),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7334aa542e79be53450da08709732f13  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib3e38e46bfa9e1bdc032918269223b32 };
assign I26781ef851ed43c6f88ff1215cddca6b = (I6a9e6c39c20e45773dab7823a7ff9486[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7334aa542e79be53450da08709732f13;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00003_U (
.flogtanh_sel( I42907182010c5889ddb7a700ead16525[flogtanh_SEL-1:0]),
.flogtanh( I659fb1602b9d248940523c14c628ce86),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ice3479ba2aeeccb88630056b7ed6b114  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I659fb1602b9d248940523c14c628ce86 };
assign Ia349e1f7c10a63ddccb3f300c73b4572 = (I42907182010c5889ddb7a700ead16525[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ice3479ba2aeeccb88630056b7ed6b114;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00004_U (
.flogtanh_sel( Ib6c26f3e3358cc2ed6fbda83eabd4bd3[flogtanh_SEL-1:0]),
.flogtanh( I1a264a901911abed928628d819c162b2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I02dba95d878330150c37c8b9ff4475fe  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1a264a901911abed928628d819c162b2 };
assign I50c4e1d3a3f63b93bc36b5141226fb3c = (Ib6c26f3e3358cc2ed6fbda83eabd4bd3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I02dba95d878330150c37c8b9ff4475fe;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00005_U (
.flogtanh_sel( Ia50d85808790790450f87a5246874b3f[flogtanh_SEL-1:0]),
.flogtanh( I2a53bd293919bc846ab816144b42592a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iecdd6e6f19312081a8d1ecfdf064e85f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2a53bd293919bc846ab816144b42592a };
assign I12334038c2be8634c47869f397503019 = (Ia50d85808790790450f87a5246874b3f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iecdd6e6f19312081a8d1ecfdf064e85f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00006_U (
.flogtanh_sel( Id4a1744702d7808a80bc40697c864765[flogtanh_SEL-1:0]),
.flogtanh( I35ce9e616a3213f2b4ce0597a47f998c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iabe6eb7899a7a53e914f54167c877c95  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I35ce9e616a3213f2b4ce0597a47f998c };
assign I64692d5168554dfd7ce1c7a046aecf72 = (Id4a1744702d7808a80bc40697c864765[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iabe6eb7899a7a53e914f54167c877c95;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00007_U (
.flogtanh_sel( I0cf3d2f3e6793a2dcf15949da16ad28d[flogtanh_SEL-1:0]),
.flogtanh( Ic3f28aa77fc84cb8e2fe43bac7ede253),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifb841b166cfe3dc103d1cd92e990ea50  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic3f28aa77fc84cb8e2fe43bac7ede253 };
assign Ia4b438844530fff602ea04e72b07db8d = (I0cf3d2f3e6793a2dcf15949da16ad28d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifb841b166cfe3dc103d1cd92e990ea50;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00008_U (
.flogtanh_sel( I90bd9107f4c931fa1ccb92998ea8cdeb[flogtanh_SEL-1:0]),
.flogtanh( I7f91c0e606b4082c6aec2e1f111079c5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4f9506d81ccabb58d8a95431289c937b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7f91c0e606b4082c6aec2e1f111079c5 };
assign I9574759e112f27778f3645d5d49126b7 = (I90bd9107f4c931fa1ccb92998ea8cdeb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4f9506d81ccabb58d8a95431289c937b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00009_U (
.flogtanh_sel( Ida1c729e6bfcec2c31a92aa9002f2c68[flogtanh_SEL-1:0]),
.flogtanh( I8e0d66c2112193437146e0f503623559),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id02f4b88464b945a30c33049c759587f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8e0d66c2112193437146e0f503623559 };
assign I2ffb7c2ad09bac694ef13ec41e5de327 = (Ida1c729e6bfcec2c31a92aa9002f2c68[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id02f4b88464b945a30c33049c759587f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00010_U (
.flogtanh_sel( Ib848feeccd0ea78ebc8ba8368534c3d1[flogtanh_SEL-1:0]),
.flogtanh( Iabe6bf045784762fb6b97be3587fd68d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I66f957fcfe83e2474c7fbfa3f6ca7fb0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iabe6bf045784762fb6b97be3587fd68d };
assign Ib190f589f4d663dbc0a3c166a8dcf5fa = (Ib848feeccd0ea78ebc8ba8368534c3d1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I66f957fcfe83e2474c7fbfa3f6ca7fb0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00011_U (
.flogtanh_sel( Icc11970bbae3adcfa33a0e5dba3e78f4[flogtanh_SEL-1:0]),
.flogtanh( I11f0fd7033065e1695d846f08d11aed5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icdbc4ac0db607b9959380b85ca6f6a7c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I11f0fd7033065e1695d846f08d11aed5 };
assign I459c59ac61179d74170db53bf45ba89e = (Icc11970bbae3adcfa33a0e5dba3e78f4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icdbc4ac0db607b9959380b85ca6f6a7c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00012_U (
.flogtanh_sel( I86bb4ef4bdd7af8861280ef30fbeeeea[flogtanh_SEL-1:0]),
.flogtanh( Ife1589d99f0764e3757de2a7d8b43008),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I889d2418e278c2787154d3bf2a3b3b38  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ife1589d99f0764e3757de2a7d8b43008 };
assign Ie5e432a991aff25577639f1b4ffd594f = (I86bb4ef4bdd7af8861280ef30fbeeeea[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I889d2418e278c2787154d3bf2a3b3b38;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00013_U (
.flogtanh_sel( I7e0c259c6c7bacdff5edc44a22e005ba[flogtanh_SEL-1:0]),
.flogtanh( I7cb3f1f2e7f997b861d6c63d55c0f4ca),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I406358d104cee15dd2b7180a1227f7bc  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7cb3f1f2e7f997b861d6c63d55c0f4ca };
assign I72064a6a84ff956d76a5aa590bbc05a9 = (I7e0c259c6c7bacdff5edc44a22e005ba[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I406358d104cee15dd2b7180a1227f7bc;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00014_U (
.flogtanh_sel( I897ddba059b27f7ed009b0cb70cfb46f[flogtanh_SEL-1:0]),
.flogtanh( Iae2f185d6338026f3e37696327f214df),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I94aea1698b59b7a5bee244015bfec001  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iae2f185d6338026f3e37696327f214df };
assign Iea74ecbac92e1b8f2ec7ad68d10b8e7d = (I897ddba059b27f7ed009b0cb70cfb46f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I94aea1698b59b7a5bee244015bfec001;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00015_U (
.flogtanh_sel( I4496243eb0542a514b551b4d09bffd7d[flogtanh_SEL-1:0]),
.flogtanh( I4da8f5b31f5cf7c70bba0cf661d727d8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib871d01d3ccfcd49906cd631b4863880  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4da8f5b31f5cf7c70bba0cf661d727d8 };
assign I4f72d0db9fcc358c6fbec9964fbe0bbb = (I4496243eb0542a514b551b4d09bffd7d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib871d01d3ccfcd49906cd631b4863880;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00016_U (
.flogtanh_sel( Ic931fb08b2e8441321ebdeed84576a0d[flogtanh_SEL-1:0]),
.flogtanh( I46dd3a6d37d3df901689403a6215b65d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3e891af010063eeb5059e18c38ca1a9f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I46dd3a6d37d3df901689403a6215b65d };
assign Ifd958901d2ea2284f506e04a058012fa = (Ic931fb08b2e8441321ebdeed84576a0d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3e891af010063eeb5059e18c38ca1a9f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00017_U (
.flogtanh_sel( Ieb6af5390b98e893ee05a939c16d2ffd[flogtanh_SEL-1:0]),
.flogtanh( I84f43bb1814bdd83a682f7a859cfd611),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I58ea1ef4bc81f85225c8028171e8a161  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I84f43bb1814bdd83a682f7a859cfd611 };
assign Ie317bbd70b9092b840c0f2713204fb9d = (Ieb6af5390b98e893ee05a939c16d2ffd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I58ea1ef4bc81f85225c8028171e8a161;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00018_U (
.flogtanh_sel( Ic2a54bad4c5a8885dd24b8687c6db0de[flogtanh_SEL-1:0]),
.flogtanh( I476ea921894e07d3f1d2ff3e7c3b660a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9f78607e0bc87e0bc7d86de85ffa838a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I476ea921894e07d3f1d2ff3e7c3b660a };
assign I2f9e56d570e72714a06c59aa9e4334c0 = (Ic2a54bad4c5a8885dd24b8687c6db0de[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9f78607e0bc87e0bc7d86de85ffa838a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00019_U (
.flogtanh_sel( I6ecbad763d2b48b78a0584beaefc78ee[flogtanh_SEL-1:0]),
.flogtanh( I5cc52764eb8a9961469e1892559ed7ee),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9f1f04e7bc9539c7aa49815fe1515427  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5cc52764eb8a9961469e1892559ed7ee };
assign I5b53fd45210b92703cb10d583f471ab9 = (I6ecbad763d2b48b78a0584beaefc78ee[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9f1f04e7bc9539c7aa49815fe1515427;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00020_U (
.flogtanh_sel( I20556d23c873c71c7ebc8a961bf40251[flogtanh_SEL-1:0]),
.flogtanh( I76f68c50b69a7545c0077f5333bfa3e2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie07e94ec114e52df8086f86dc5fbc424  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I76f68c50b69a7545c0077f5333bfa3e2 };
assign I8edbe77bacf1975e014faeee6b861980 = (I20556d23c873c71c7ebc8a961bf40251[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie07e94ec114e52df8086f86dc5fbc424;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00021_U (
.flogtanh_sel( I79012e6351e6320c22437aa216ea4df1[flogtanh_SEL-1:0]),
.flogtanh( Id0bd4407ef72994435b3794096636553),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia048dc6a01575d1733276742fd45bdf5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id0bd4407ef72994435b3794096636553 };
assign I174fcbc2ee01fc55edbc8238e5da7f0c = (I79012e6351e6320c22437aa216ea4df1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia048dc6a01575d1733276742fd45bdf5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00006_00022_U (
.flogtanh_sel( Ibf74ab9af877d27c3a6f3881f00ddaf1[flogtanh_SEL-1:0]),
.flogtanh( I0879a96ba0ef5eb523ae807c40c66a63),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ice646ce92235cc21cb7fc0799053b50a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0879a96ba0ef5eb523ae807c40c66a63 };
assign Id4dc304aef5f35f6ceb91796c278e716 = (Ibf74ab9af877d27c3a6f3881f00ddaf1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ice646ce92235cc21cb7fc0799053b50a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00000_U (
.flogtanh_sel( I843d35db35d7b42a87ce78d3772cec2f[flogtanh_SEL-1:0]),
.flogtanh( I8304ab4dc851d69a7ad7db75ced3eb9e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6ea1aaf77ecc0369ff33b58439a99d1b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8304ab4dc851d69a7ad7db75ced3eb9e };
assign I0cbdfae6f75a639eb591d9c0022f5838 = (I843d35db35d7b42a87ce78d3772cec2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6ea1aaf77ecc0369ff33b58439a99d1b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00001_U (
.flogtanh_sel( I2b1398b4bfd374d7221b0a68da28e979[flogtanh_SEL-1:0]),
.flogtanh( I24d773b608ba1ee21855540ee84028da),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I93eed7c401e8f511efa112a82b9b9a4f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I24d773b608ba1ee21855540ee84028da };
assign I088898ee932a96c14f2f0f568f5455b6 = (I2b1398b4bfd374d7221b0a68da28e979[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I93eed7c401e8f511efa112a82b9b9a4f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00002_U (
.flogtanh_sel( I6f615d6e74b0c02f8e4265523ad16404[flogtanh_SEL-1:0]),
.flogtanh( I9458b9a213600ce0c8c1d54d31c8c5c2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9ef8088456f239e42f67e7b0ec062c35  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9458b9a213600ce0c8c1d54d31c8c5c2 };
assign Ide0abde3644a4fafb436aa59768d016e = (I6f615d6e74b0c02f8e4265523ad16404[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9ef8088456f239e42f67e7b0ec062c35;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00003_U (
.flogtanh_sel( Iae8a98dd4a7cbfbc56c1404b6a2020af[flogtanh_SEL-1:0]),
.flogtanh( Idb6b8e6f2df9b8d96efa93830df86a71),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5529826cbbfacc566e550b2fb6d34200  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idb6b8e6f2df9b8d96efa93830df86a71 };
assign I08581dc8d42be712cfb36d744f2786e0 = (Iae8a98dd4a7cbfbc56c1404b6a2020af[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5529826cbbfacc566e550b2fb6d34200;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00004_U (
.flogtanh_sel( Iad53375a54d01c559c74981bf279dfb5[flogtanh_SEL-1:0]),
.flogtanh( I0a8fb8a7a28b364bc8cf49b96fdc66a4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I71d41f3f13a20950a8f5e5dace0b9754  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0a8fb8a7a28b364bc8cf49b96fdc66a4 };
assign I29fb3830a5fc5922f1ec687a38941e97 = (Iad53375a54d01c559c74981bf279dfb5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I71d41f3f13a20950a8f5e5dace0b9754;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00005_U (
.flogtanh_sel( I5db1307f922e0c742d7d9f3a79a4a4f3[flogtanh_SEL-1:0]),
.flogtanh( I938f8896ddbf95751aea2b327f5d40f0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id031c3a3b6acda879451d8d73153bc49  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I938f8896ddbf95751aea2b327f5d40f0 };
assign I715d59fb27e519a9b76bdd8b5139a619 = (I5db1307f922e0c742d7d9f3a79a4a4f3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id031c3a3b6acda879451d8d73153bc49;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00006_U (
.flogtanh_sel( I9f78172ed5bf73752196f9a8810005f3[flogtanh_SEL-1:0]),
.flogtanh( Ib5b964583d3ef33b47643ca212bc0ada),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idf0dedc8613d3ebf20cfbbe7d4337be9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib5b964583d3ef33b47643ca212bc0ada };
assign Ibe6a876a041198a581c95457a7d1fcf8 = (I9f78172ed5bf73752196f9a8810005f3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idf0dedc8613d3ebf20cfbbe7d4337be9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00007_U (
.flogtanh_sel( If85a22d670d47f491dd7568d0453ba1d[flogtanh_SEL-1:0]),
.flogtanh( I4bae2a264af742ffe7be73f9a1129efe),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I034f9d302ce082349a9d812c9fe46411  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4bae2a264af742ffe7be73f9a1129efe };
assign Iec078a95a69b081cfb5e987ba9c5a613 = (If85a22d670d47f491dd7568d0453ba1d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I034f9d302ce082349a9d812c9fe46411;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00008_U (
.flogtanh_sel( Ib9e529170b2896e930a839295796fd31[flogtanh_SEL-1:0]),
.flogtanh( I041c1a7ef6128c7a1a8f8593d4401f1b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id1ad76a0501d9ea66134873e99cb211d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I041c1a7ef6128c7a1a8f8593d4401f1b };
assign I0e8f3f56bce3be1ee4d5f780a2f2a9fe = (Ib9e529170b2896e930a839295796fd31[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id1ad76a0501d9ea66134873e99cb211d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00009_U (
.flogtanh_sel( Ib7af536846bac40c1f221d1f72c6c25c[flogtanh_SEL-1:0]),
.flogtanh( I22c6d2c87ef183ef45805a7c99a7e473),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iec5b39a66a2fd9920c3bed36edb32f02  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I22c6d2c87ef183ef45805a7c99a7e473 };
assign Ia73cacadbf80c0701a5b5b430c0d5c98 = (Ib7af536846bac40c1f221d1f72c6c25c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iec5b39a66a2fd9920c3bed36edb32f02;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00010_U (
.flogtanh_sel( Ib0eb61a2cb831dd35ce9850994e7c2da[flogtanh_SEL-1:0]),
.flogtanh( I45fef5261954fc84be265f39eb8f9647),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iedeaa45a179ec994bce6b6cc6da0995c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I45fef5261954fc84be265f39eb8f9647 };
assign Ic634d26fc09589a29a160e4efb5613a8 = (Ib0eb61a2cb831dd35ce9850994e7c2da[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iedeaa45a179ec994bce6b6cc6da0995c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00011_U (
.flogtanh_sel( I89d338f59960af7a47595d6afa206abc[flogtanh_SEL-1:0]),
.flogtanh( I3b292cf842e3a7ca9e6d0c4ab345446f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I915031fb071f83ac6eb7357933151d20  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3b292cf842e3a7ca9e6d0c4ab345446f };
assign Ie1374cac341cf353b1863dae9f544e8b = (I89d338f59960af7a47595d6afa206abc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I915031fb071f83ac6eb7357933151d20;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00012_U (
.flogtanh_sel( Ib3c1176eb8991e3e85855a9fe845c303[flogtanh_SEL-1:0]),
.flogtanh( Ie7bff678d39738eb49b599772586210a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If7df947e519a3cd29b42434a9519fbb5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie7bff678d39738eb49b599772586210a };
assign Ia07447985347e9a7f3739bd98867cdfb = (Ib3c1176eb8991e3e85855a9fe845c303[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If7df947e519a3cd29b42434a9519fbb5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00013_U (
.flogtanh_sel( I93073d05d509b821a743998cf32c58ee[flogtanh_SEL-1:0]),
.flogtanh( Ib9d80aab3818d682b54122974fa3a424),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5bac22cea76db3326f60e45aa8ed14c1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib9d80aab3818d682b54122974fa3a424 };
assign I2121318f589878b4a9260625f97de518 = (I93073d05d509b821a743998cf32c58ee[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5bac22cea76db3326f60e45aa8ed14c1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00014_U (
.flogtanh_sel( Iab6dac1909c1564c3890ffecc13418df[flogtanh_SEL-1:0]),
.flogtanh( Iaa05186a94ba0559ab57ced9202ccefb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2e9180aad8498bc69a9c74af78238e6d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iaa05186a94ba0559ab57ced9202ccefb };
assign Ibd8424c228f87f85df3da6204edff2b5 = (Iab6dac1909c1564c3890ffecc13418df[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2e9180aad8498bc69a9c74af78238e6d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00015_U (
.flogtanh_sel( I1b75eeb29167a171d89f6e67039436d5[flogtanh_SEL-1:0]),
.flogtanh( I506f39735c3743b3705980c73295c035),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id965c3c3f0ab3fc022737b6b577ad6e0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I506f39735c3743b3705980c73295c035 };
assign I8a7fb51566bf215af214cd2fb5209974 = (I1b75eeb29167a171d89f6e67039436d5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id965c3c3f0ab3fc022737b6b577ad6e0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00016_U (
.flogtanh_sel( I3a31adc52a1405555017b2ddf219b407[flogtanh_SEL-1:0]),
.flogtanh( I8f16ead6735608b15b364b9af9b3a22a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0ecfcdb358eb5e5ed3eb9c5f3f137dd0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8f16ead6735608b15b364b9af9b3a22a };
assign I7c0f872988488ac69815d288885dfd2f = (I3a31adc52a1405555017b2ddf219b407[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0ecfcdb358eb5e5ed3eb9c5f3f137dd0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00017_U (
.flogtanh_sel( Iaadba89c6a370240fc0758029f7d8db0[flogtanh_SEL-1:0]),
.flogtanh( Id07af023803badc88c51b891cad1b7e5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I094f9bedec7e86f01b6f7e223d13b82f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id07af023803badc88c51b891cad1b7e5 };
assign I3521b10b97b0e74888ce385cfc772945 = (Iaadba89c6a370240fc0758029f7d8db0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I094f9bedec7e86f01b6f7e223d13b82f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00018_U (
.flogtanh_sel( I4f4a64fb3ced7d9f7ee4513178e9655a[flogtanh_SEL-1:0]),
.flogtanh( Iecb522fa10764b2c0c044be6c1ca807d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib67397a1a44a6cfd5ea04983f1847686  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iecb522fa10764b2c0c044be6c1ca807d };
assign I58f0b81a46549cab8e74ecbc285df23a = (I4f4a64fb3ced7d9f7ee4513178e9655a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib67397a1a44a6cfd5ea04983f1847686;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00019_U (
.flogtanh_sel( I0c76ca58f69c91758e755cd581241284[flogtanh_SEL-1:0]),
.flogtanh( I58b9a09be96353ba6c18f310e1987742),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2e49a1e612abcd98120c4528eda7c359  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I58b9a09be96353ba6c18f310e1987742 };
assign I7095040b38bf9d6b5229c11d2a0d7c57 = (I0c76ca58f69c91758e755cd581241284[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2e49a1e612abcd98120c4528eda7c359;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00020_U (
.flogtanh_sel( I2312bce18958346149c868846e04643b[flogtanh_SEL-1:0]),
.flogtanh( I86ced95bff4327e4ab07338663f82029),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id87382649fe91c747a380e2ec4e4cdcd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I86ced95bff4327e4ab07338663f82029 };
assign I675ab6c4fb93b006f3fcafc985fbc405 = (I2312bce18958346149c868846e04643b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id87382649fe91c747a380e2ec4e4cdcd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00021_U (
.flogtanh_sel( I3e154098cb0a48f1c23234f46613f406[flogtanh_SEL-1:0]),
.flogtanh( Ia802328754db2d72d6ec8e12a79b2341),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia29f77138da85cd201325cc411528c73  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia802328754db2d72d6ec8e12a79b2341 };
assign I239a992ebb62899120a74b1c9e6cc4b4 = (I3e154098cb0a48f1c23234f46613f406[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia29f77138da85cd201325cc411528c73;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00007_00022_U (
.flogtanh_sel( I1645c1c588bcbf15dd62d47e08b8e139[flogtanh_SEL-1:0]),
.flogtanh( I5b5a9fa50a6e4c7e07017249e5dee137),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I29ffc08244342190be5b2adcb968fbea  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5b5a9fa50a6e4c7e07017249e5dee137 };
assign I927c870d09285dcb47e6d399f319471e = (I1645c1c588bcbf15dd62d47e08b8e139[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I29ffc08244342190be5b2adcb968fbea;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00008_00000_U (
.flogtanh_sel( I4c25de66590e1745d37112e08d8c8e2c[flogtanh_SEL-1:0]),
.flogtanh( I73ef262450353dfcfabe3051ab0006f9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I58ea03377afb90bb2f408efebc0fe7eb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I73ef262450353dfcfabe3051ab0006f9 };
assign Ie23ed3ee61f468f59f2baf661cb7f85d = (I4c25de66590e1745d37112e08d8c8e2c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I58ea03377afb90bb2f408efebc0fe7eb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00008_00001_U (
.flogtanh_sel( Ia03092ac621b8dd1c206fea1e8b0215f[flogtanh_SEL-1:0]),
.flogtanh( I959c5d62629333d1d60766a6d935ae4a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5f7e827df9d731c1ffd418b1ad028b31  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I959c5d62629333d1d60766a6d935ae4a };
assign I68e58664be09261e5a80d6f8ecdd1b60 = (Ia03092ac621b8dd1c206fea1e8b0215f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5f7e827df9d731c1ffd418b1ad028b31;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00008_00002_U (
.flogtanh_sel( I5c9bdb033436dc9f6069baca31f24c2d[flogtanh_SEL-1:0]),
.flogtanh( I659d579ea5b5d24ef0ccbb8160dfe2ae),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6e5a9a96c90b19eb113510e4dc7fe113  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I659d579ea5b5d24ef0ccbb8160dfe2ae };
assign Id2808e0f40992c79ead4da7c734e5b79 = (I5c9bdb033436dc9f6069baca31f24c2d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6e5a9a96c90b19eb113510e4dc7fe113;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00008_00003_U (
.flogtanh_sel( I8f07cf4865480f18ad6945974ec2231c[flogtanh_SEL-1:0]),
.flogtanh( Icae3ba8a84ee6ee051a3caf210f47b51),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9a1438cdffb8de6db7d253106895fd6c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icae3ba8a84ee6ee051a3caf210f47b51 };
assign Icb2b390266bff241a688961136db0f51 = (I8f07cf4865480f18ad6945974ec2231c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9a1438cdffb8de6db7d253106895fd6c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00008_00004_U (
.flogtanh_sel( I4a7119e8862fe4a6a4100dd9ac67dd24[flogtanh_SEL-1:0]),
.flogtanh( I92a005abe2d27beb2949fe29c0d8bc65),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I972c89a3fa5af605d673f846c71f8f57  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I92a005abe2d27beb2949fe29c0d8bc65 };
assign I54cfd68212d97a2cc8241ef429429453 = (I4a7119e8862fe4a6a4100dd9ac67dd24[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I972c89a3fa5af605d673f846c71f8f57;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00008_00005_U (
.flogtanh_sel( Id78fcfc6724a05f46d44d7c3e7d0c756[flogtanh_SEL-1:0]),
.flogtanh( I28fb1164936618d653aa7bf06c03b38f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6cdde8c6984cc120c0f0a1a0472d50c5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I28fb1164936618d653aa7bf06c03b38f };
assign I8d4e3962525c424786ae822a6981a5e6 = (Id78fcfc6724a05f46d44d7c3e7d0c756[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6cdde8c6984cc120c0f0a1a0472d50c5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00008_00006_U (
.flogtanh_sel( I7cbd9d619623cbabf8ed6b1fece8f012[flogtanh_SEL-1:0]),
.flogtanh( I8720bdf2c91f113b39aa5b6f82421feb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id2f5757d8a8432506fbffa192a4e0c49  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8720bdf2c91f113b39aa5b6f82421feb };
assign I1a5f22b4e326d1684c0a8c7a7e754ab4 = (I7cbd9d619623cbabf8ed6b1fece8f012[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id2f5757d8a8432506fbffa192a4e0c49;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00008_00007_U (
.flogtanh_sel( I58951165d251e370b0f3b3fb537aed18[flogtanh_SEL-1:0]),
.flogtanh( I07320e5fb3beddb93ae325a98c5e3782),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iefdb7ed85a168a0fa2e5e93d1d67701e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I07320e5fb3beddb93ae325a98c5e3782 };
assign I8c2e0c83a8204d6b21e0e3e458d56f05 = (I58951165d251e370b0f3b3fb537aed18[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iefdb7ed85a168a0fa2e5e93d1d67701e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00008_00008_U (
.flogtanh_sel( I21daac106f526d84cb8fa5239c19499d[flogtanh_SEL-1:0]),
.flogtanh( Ib8b29bc86ad9c07d7ae5b358f66cb9ba),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If1f93a57723e97173a4289a0052945b8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib8b29bc86ad9c07d7ae5b358f66cb9ba };
assign Ie0622ff815747e4a9f368c74787026ec = (I21daac106f526d84cb8fa5239c19499d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If1f93a57723e97173a4289a0052945b8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00008_00009_U (
.flogtanh_sel( I178029cec3a5d6141abdfa91b91fdbf4[flogtanh_SEL-1:0]),
.flogtanh( I8e2ed2040f5bf8ea125e5b953cf89300),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia5ec300f6b8946d5e6ff0cfb22eba4ed  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8e2ed2040f5bf8ea125e5b953cf89300 };
assign I5ffed139764d90825b9f2eddacd0eddc = (I178029cec3a5d6141abdfa91b91fdbf4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia5ec300f6b8946d5e6ff0cfb22eba4ed;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00009_00000_U (
.flogtanh_sel( I96dfb2efbb55a644616e3474ed07c364[flogtanh_SEL-1:0]),
.flogtanh( I4ad3a5b591cd6b13de04897fbbd068ec),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0c27572b0776655756ce831c506bef53  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4ad3a5b591cd6b13de04897fbbd068ec };
assign I5a3297f48e1045273db6522744582b05 = (I96dfb2efbb55a644616e3474ed07c364[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0c27572b0776655756ce831c506bef53;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00009_00001_U (
.flogtanh_sel( I7a17d8f0e2d16c441044db68ee037731[flogtanh_SEL-1:0]),
.flogtanh( If5208f94e99b0e7ff353c048b55ad7ba),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I088d29bd92758302c48dabb469993251  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If5208f94e99b0e7ff353c048b55ad7ba };
assign I9858bb2a3cc458aca5bf7eb077ee55dd = (I7a17d8f0e2d16c441044db68ee037731[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I088d29bd92758302c48dabb469993251;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00009_00002_U (
.flogtanh_sel( I2ced9bb3ae6bdc5b5ef2865fb46abf07[flogtanh_SEL-1:0]),
.flogtanh( I66106fad536bb49418e7d09e3f4221ac),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iec3bf0eb952518b856f1596f964e3ae5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I66106fad536bb49418e7d09e3f4221ac };
assign I6e7e27bb176196e4493bf9c45ca19719 = (I2ced9bb3ae6bdc5b5ef2865fb46abf07[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iec3bf0eb952518b856f1596f964e3ae5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00009_00003_U (
.flogtanh_sel( I89a93384020d93cf4d26b3902e06cd9e[flogtanh_SEL-1:0]),
.flogtanh( I6af88c096ca3af849bbedb15b2ac7153),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I990ed4f7284e44d83197a4cc987c8ff1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6af88c096ca3af849bbedb15b2ac7153 };
assign I4cff1804df738cbf4f940c775236df9c = (I89a93384020d93cf4d26b3902e06cd9e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I990ed4f7284e44d83197a4cc987c8ff1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00009_00004_U (
.flogtanh_sel( Ibbb47d29b9a45559c13ffa3b046c66f5[flogtanh_SEL-1:0]),
.flogtanh( I15d6e1e431457b954b5f86cd4fb16a77),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7d0dc027656ba91703f0ac89aae218d3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I15d6e1e431457b954b5f86cd4fb16a77 };
assign I0c1e22375d5e023c24519901b92eceb5 = (Ibbb47d29b9a45559c13ffa3b046c66f5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7d0dc027656ba91703f0ac89aae218d3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00009_00005_U (
.flogtanh_sel( I0034177eb1049577a3578b371527f34b[flogtanh_SEL-1:0]),
.flogtanh( Ifd67d6dec292171610a805560d7cb9a0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I421d6fb792792366ca3d3bf8f8520f56  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifd67d6dec292171610a805560d7cb9a0 };
assign Ida5b16851dc06534844a0b037d74feb3 = (I0034177eb1049577a3578b371527f34b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I421d6fb792792366ca3d3bf8f8520f56;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00009_00006_U (
.flogtanh_sel( I22d9ea7bb5a1a3405bcd04b9af40fa62[flogtanh_SEL-1:0]),
.flogtanh( I681c4ec303ff366746d35234fe5a1ff4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If538078378e360ac004d4b122f75cb42  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I681c4ec303ff366746d35234fe5a1ff4 };
assign Iac3cb5b4481687fcf430c8bf52cfb74d = (I22d9ea7bb5a1a3405bcd04b9af40fa62[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If538078378e360ac004d4b122f75cb42;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00009_00007_U (
.flogtanh_sel( I8a632e7a911bf5726fee587189cb6f16[flogtanh_SEL-1:0]),
.flogtanh( I5df2eac3ace0bcef9e48b0850d975cce),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia144749f2f8b6f0e06f00dd3a6954616  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5df2eac3ace0bcef9e48b0850d975cce };
assign Ia1499972c4995268acd828c1289f353d = (I8a632e7a911bf5726fee587189cb6f16[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia144749f2f8b6f0e06f00dd3a6954616;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00009_00008_U (
.flogtanh_sel( I3765afc490b34e8a310998a4ebcff8cb[flogtanh_SEL-1:0]),
.flogtanh( Icf6f5254160a82036c4ba0367e8f0404),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8dff03248f37764bfe0c2c6b4fcc795f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icf6f5254160a82036c4ba0367e8f0404 };
assign Ie559401a3a913400dc5e3e5641297fa6 = (I3765afc490b34e8a310998a4ebcff8cb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8dff03248f37764bfe0c2c6b4fcc795f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00009_00009_U (
.flogtanh_sel( I7607e800ae46a96e016b303120da4247[flogtanh_SEL-1:0]),
.flogtanh( If1de12bbb90e49cc1b28eafc2aa551e5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5d98e3e3fbce58307f7df7fc7d580ac8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If1de12bbb90e49cc1b28eafc2aa551e5 };
assign Ie0667fbe76244eaec0b155d69dcc9447 = (I7607e800ae46a96e016b303120da4247[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5d98e3e3fbce58307f7df7fc7d580ac8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00010_00000_U (
.flogtanh_sel( I29b2f1fddee5e32f217d25410bcfce4f[flogtanh_SEL-1:0]),
.flogtanh( Ibf9f7f1f6a759af21ac82d6e6ff7df43),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia47119d76cf6a40b200cd5ecfd4b1409  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibf9f7f1f6a759af21ac82d6e6ff7df43 };
assign I1d0f031e8ae9c0335d501d1565118220 = (I29b2f1fddee5e32f217d25410bcfce4f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia47119d76cf6a40b200cd5ecfd4b1409;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00010_00001_U (
.flogtanh_sel( Iba5f8a31a81f6aa06f5e38c03dc6db54[flogtanh_SEL-1:0]),
.flogtanh( Ie44bc9632854c4c2077bcec5f46d29ad),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia10ec5bac071d9ad1941489d7457e0ef  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie44bc9632854c4c2077bcec5f46d29ad };
assign Ie2c801b2de066c3218d7312615b7bfda = (Iba5f8a31a81f6aa06f5e38c03dc6db54[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia10ec5bac071d9ad1941489d7457e0ef;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00010_00002_U (
.flogtanh_sel( Ifcb5c907ad503331317599e4e0ce7be8[flogtanh_SEL-1:0]),
.flogtanh( I97ae894cd928e17cad4c4631aec2c7a0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I048bdd98d2fdac75bdae08d64fa7ef22  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I97ae894cd928e17cad4c4631aec2c7a0 };
assign I64c4bb0d40d80ec52aab61ce46954f43 = (Ifcb5c907ad503331317599e4e0ce7be8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I048bdd98d2fdac75bdae08d64fa7ef22;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00010_00003_U (
.flogtanh_sel( I62d6f2ab4ec8b6ecfa544ad4d90eb30b[flogtanh_SEL-1:0]),
.flogtanh( I500a903104b4b532b3c07d1640e80b55),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie8075a19a463a00c303aea3814991070  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I500a903104b4b532b3c07d1640e80b55 };
assign I512f57a40c7c8cb2f040bdde73e44ca3 = (I62d6f2ab4ec8b6ecfa544ad4d90eb30b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie8075a19a463a00c303aea3814991070;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00010_00004_U (
.flogtanh_sel( Ide65414c51b3cb182c0f2f238903d60a[flogtanh_SEL-1:0]),
.flogtanh( I1d3ae54c8fa3d87a39e3a51018a20727),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaa6e4f7efa27d63fff2fae677e914cdb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1d3ae54c8fa3d87a39e3a51018a20727 };
assign Id60cbf534604e5dba988050ef5abe625 = (Ide65414c51b3cb182c0f2f238903d60a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaa6e4f7efa27d63fff2fae677e914cdb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00010_00005_U (
.flogtanh_sel( I03a8dc2288eaeb619e746990e20cc868[flogtanh_SEL-1:0]),
.flogtanh( I23d3b6da58b66185ddb3c5eae0f68dae),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3eb15cc35c68ee4a5f5294eb5b993259  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I23d3b6da58b66185ddb3c5eae0f68dae };
assign I37998a91d20db2248ebdd8e661d42f70 = (I03a8dc2288eaeb619e746990e20cc868[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3eb15cc35c68ee4a5f5294eb5b993259;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00010_00006_U (
.flogtanh_sel( Id81c1b44d16ddbcd466382c60fe84986[flogtanh_SEL-1:0]),
.flogtanh( I88b1352db9aa35be019bc0f345c7131e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I094201803df7b2720fd55ca7a7d870c4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I88b1352db9aa35be019bc0f345c7131e };
assign Ib65ff82aff398f6ff7ba711a36f41ee4 = (Id81c1b44d16ddbcd466382c60fe84986[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I094201803df7b2720fd55ca7a7d870c4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00010_00007_U (
.flogtanh_sel( I503d72f4a2fd20dbf35aa27321d2ede7[flogtanh_SEL-1:0]),
.flogtanh( I1115071c073981f4db4917844fb12a73),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3831fdb5ff3d1597900808314bfa0fd5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1115071c073981f4db4917844fb12a73 };
assign I3d1dd8b9c7c6d3913f7ac369ad7e625c = (I503d72f4a2fd20dbf35aa27321d2ede7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3831fdb5ff3d1597900808314bfa0fd5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00010_00008_U (
.flogtanh_sel( Id6595a4cf33062d1f05cbcee2d0685f1[flogtanh_SEL-1:0]),
.flogtanh( Ia9e4e593fd82657c81aeea8fbcd1194b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I092c808c76ddb6c2dc97a552d1f903cf  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia9e4e593fd82657c81aeea8fbcd1194b };
assign I097722547450582dc5776bdaff914741 = (Id6595a4cf33062d1f05cbcee2d0685f1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I092c808c76ddb6c2dc97a552d1f903cf;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00010_00009_U (
.flogtanh_sel( I83ebdd7331ca8fbcf5250851b346c0b0[flogtanh_SEL-1:0]),
.flogtanh( I22300986ed621a97a6dac1f3b4d59b8e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I21dc24999451f1e4d8f14813d7d0e58d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I22300986ed621a97a6dac1f3b4d59b8e };
assign Id4a213e494f9c9be0fd1a307e87c756a = (I83ebdd7331ca8fbcf5250851b346c0b0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I21dc24999451f1e4d8f14813d7d0e58d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00011_00000_U (
.flogtanh_sel( I7f6ea26cdfe5986065e7b5aa6842cc1c[flogtanh_SEL-1:0]),
.flogtanh( Icc08ab7c64b40e53278a93f4ae0f9209),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I779162012544d75b0d1559145dd29468  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icc08ab7c64b40e53278a93f4ae0f9209 };
assign I21594c8b0169efd7c2aa6cbc31f4a901 = (I7f6ea26cdfe5986065e7b5aa6842cc1c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I779162012544d75b0d1559145dd29468;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00011_00001_U (
.flogtanh_sel( Idab1ec32c20f93c4cc1acb38158f92d5[flogtanh_SEL-1:0]),
.flogtanh( I8cc9f5531f2675b3058df110912551b6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0c0f66943d6470070aeddf77435e28f7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8cc9f5531f2675b3058df110912551b6 };
assign I15022e1b349eee259d3567837283dbf6 = (Idab1ec32c20f93c4cc1acb38158f92d5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0c0f66943d6470070aeddf77435e28f7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00011_00002_U (
.flogtanh_sel( I0738add83419502e73674ded2f1ad6c7[flogtanh_SEL-1:0]),
.flogtanh( Icdba6332ba9ea91ffefd690150fba09f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I30faa261a877ce65b3a057bae448bf7f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icdba6332ba9ea91ffefd690150fba09f };
assign I1070940dc2ef6e8ee3d1227ec9ff3162 = (I0738add83419502e73674ded2f1ad6c7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I30faa261a877ce65b3a057bae448bf7f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00011_00003_U (
.flogtanh_sel( I6c93e63a8e5a2dbd598f1565c7323b39[flogtanh_SEL-1:0]),
.flogtanh( Idaef789d04cd5c6291dae88f616460e6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia0f7dfeea453a44869ad21670b100db5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idaef789d04cd5c6291dae88f616460e6 };
assign I8922cc37cde6ba132f632743113e42af = (I6c93e63a8e5a2dbd598f1565c7323b39[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia0f7dfeea453a44869ad21670b100db5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00011_00004_U (
.flogtanh_sel( I4aa57a9d46371f1680d5f95596f60b5d[flogtanh_SEL-1:0]),
.flogtanh( I016cb9c8307b28a7cabf9a91e8da03d6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I32165a54dc2b00d05357e4512ff40ae3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I016cb9c8307b28a7cabf9a91e8da03d6 };
assign Ia66c399023e500ed67197dcf236f5d42 = (I4aa57a9d46371f1680d5f95596f60b5d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I32165a54dc2b00d05357e4512ff40ae3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00011_00005_U (
.flogtanh_sel( I5369a7203b78951a3c006c2d3b22507c[flogtanh_SEL-1:0]),
.flogtanh( I54517f62dd6f2e7de7d522dfc506383e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I94df0a38de39d37156cb5d84f3c360fc  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I54517f62dd6f2e7de7d522dfc506383e };
assign I1171dc208d5db1024dc3f09a90c78ca0 = (I5369a7203b78951a3c006c2d3b22507c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I94df0a38de39d37156cb5d84f3c360fc;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00011_00006_U (
.flogtanh_sel( Ie72a79a6966cf198687b7c8a8bcdeb13[flogtanh_SEL-1:0]),
.flogtanh( I6b0c1ef6f0a94adaf62425829edf28dd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I85c46907cc9da850a5123a2140d7d75c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6b0c1ef6f0a94adaf62425829edf28dd };
assign Ic28b148967a5b3d05409976fa9001ac8 = (Ie72a79a6966cf198687b7c8a8bcdeb13[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I85c46907cc9da850a5123a2140d7d75c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00011_00007_U (
.flogtanh_sel( Ie917ae4c44ab0f9c2f1747ff0d2a754e[flogtanh_SEL-1:0]),
.flogtanh( I067ce754b1084de762c33b295f2f47b2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib09c12fe109a9604c5877b84c0d09874  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I067ce754b1084de762c33b295f2f47b2 };
assign I79fe46308b93fbb24245fe1c75edf4a5 = (Ie917ae4c44ab0f9c2f1747ff0d2a754e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib09c12fe109a9604c5877b84c0d09874;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00011_00008_U (
.flogtanh_sel( I0b1a31ccb34a742552c11b1945e23dd8[flogtanh_SEL-1:0]),
.flogtanh( Ib2fe88cfe23c363993dfcb7722c4fef0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4e8f05ec6bda855c0625055f7d7d015e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib2fe88cfe23c363993dfcb7722c4fef0 };
assign I3bfcd63e92f1949234ab1d2701dbb499 = (I0b1a31ccb34a742552c11b1945e23dd8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4e8f05ec6bda855c0625055f7d7d015e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00011_00009_U (
.flogtanh_sel( I9a65a845cf2eced39050e8481665f557[flogtanh_SEL-1:0]),
.flogtanh( I71f836227a1f7f81500a6c980c06f1f7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If3e09ed5717deb2229298308143c32ce  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I71f836227a1f7f81500a6c980c06f1f7 };
assign I5e2331edf6e881e9f3a8c47eebda0ac4 = (I9a65a845cf2eced39050e8481665f557[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If3e09ed5717deb2229298308143c32ce;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00012_00000_U (
.flogtanh_sel( I3b402b35d38a9fde312c89b82297c1a5[flogtanh_SEL-1:0]),
.flogtanh( I6faf34757a61a0b64e61ba059aca33fa),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6cf5a36287d132e0eb71d9006b816cf9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6faf34757a61a0b64e61ba059aca33fa };
assign I4b66c202450986ef0df05e979cc8bc7f = (I3b402b35d38a9fde312c89b82297c1a5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6cf5a36287d132e0eb71d9006b816cf9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00012_00001_U (
.flogtanh_sel( I309fa33562370e339c19e2377e6a6a7a[flogtanh_SEL-1:0]),
.flogtanh( Ib1821b79b79aadf1486fe1e2df2f297c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If651c14f270904442ab9c299d25a4c16  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib1821b79b79aadf1486fe1e2df2f297c };
assign I737daf208eccf95feb3192897586cdce = (I309fa33562370e339c19e2377e6a6a7a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If651c14f270904442ab9c299d25a4c16;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00012_00002_U (
.flogtanh_sel( I7d06aed81222a030837cad2074c68e19[flogtanh_SEL-1:0]),
.flogtanh( I84daf07d3f3790c691b9192f7e2018c1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iebc916f489d40512cab9ad4494fe3405  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I84daf07d3f3790c691b9192f7e2018c1 };
assign I29c8133231cfda17668bbe7b692bdfe2 = (I7d06aed81222a030837cad2074c68e19[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iebc916f489d40512cab9ad4494fe3405;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00012_00003_U (
.flogtanh_sel( I835cc6af0cd8189035f2441c2e0d3100[flogtanh_SEL-1:0]),
.flogtanh( Ib4b3ed1f9d1dee96a3ec846424412e2f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5a0259d2bf5c8a842f607743dcff5851  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib4b3ed1f9d1dee96a3ec846424412e2f };
assign Id9d56f09595e80d66c2ac300f7d1d972 = (I835cc6af0cd8189035f2441c2e0d3100[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5a0259d2bf5c8a842f607743dcff5851;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00012_00004_U (
.flogtanh_sel( If6f768d12f04087246a0d65de1aef99b[flogtanh_SEL-1:0]),
.flogtanh( Ibe73f00bb6f1494ede2e6f11f5e7d3f8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icac9d2c51408fe77883a998c48953a3a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibe73f00bb6f1494ede2e6f11f5e7d3f8 };
assign I97e89a2ee18d2688d7c1a640318a1e0d = (If6f768d12f04087246a0d65de1aef99b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icac9d2c51408fe77883a998c48953a3a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00013_00000_U (
.flogtanh_sel( Ie4b180e1e2cadb865b0eaf6509f99dbb[flogtanh_SEL-1:0]),
.flogtanh( I1542461b996a466d7d3d50bb48ebd690),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icaca84de45cecbfbbc4613ee6b1ebd78  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1542461b996a466d7d3d50bb48ebd690 };
assign Ife123bf57fe693dabe6aeaa236c4e058 = (Ie4b180e1e2cadb865b0eaf6509f99dbb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icaca84de45cecbfbbc4613ee6b1ebd78;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00013_00001_U (
.flogtanh_sel( Ie329a11fc3f6f59f6f1790612fde3250[flogtanh_SEL-1:0]),
.flogtanh( If97a5a2c523f51c5881496c5dc8ad11e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2dc2f2119d90018c1376658e22e66c56  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If97a5a2c523f51c5881496c5dc8ad11e };
assign I0c0d844fe3b7d35c1ed6bd7cc4e0dc24 = (Ie329a11fc3f6f59f6f1790612fde3250[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2dc2f2119d90018c1376658e22e66c56;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00013_00002_U (
.flogtanh_sel( Idb7ddbee4076f7bf49177e69f5e4d112[flogtanh_SEL-1:0]),
.flogtanh( Ie19ea558cf2a95ca0c8ae769a809d908),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If570315645da3ffaedc01b9bb830e1e5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie19ea558cf2a95ca0c8ae769a809d908 };
assign I2d9632ae6a0f3ba44c3da8f56ba3fedf = (Idb7ddbee4076f7bf49177e69f5e4d112[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If570315645da3ffaedc01b9bb830e1e5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00013_00003_U (
.flogtanh_sel( I614d66a7dca2d08efdfdc157ca803d5c[flogtanh_SEL-1:0]),
.flogtanh( I6532e6299b8c1fdf7f61b3a44b61c35c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id5083f0249f7b1bd62260a38e2ad71c9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6532e6299b8c1fdf7f61b3a44b61c35c };
assign I38cc7b117c0bcd5e3060cd370d710d7e = (I614d66a7dca2d08efdfdc157ca803d5c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id5083f0249f7b1bd62260a38e2ad71c9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00013_00004_U (
.flogtanh_sel( Iea16eb0ab70ebb1bc47ae55e11ced62d[flogtanh_SEL-1:0]),
.flogtanh( Ic7102fb8b5df222fff6151e8794bec3c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7b4308ad008be7a70f2d1d5d7a259479  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic7102fb8b5df222fff6151e8794bec3c };
assign I793ddbf6a5d026a57ab72984ca19deac = (Iea16eb0ab70ebb1bc47ae55e11ced62d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7b4308ad008be7a70f2d1d5d7a259479;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00014_00000_U (
.flogtanh_sel( Ifa8db43284d5bbebaed4f72d65cf9f92[flogtanh_SEL-1:0]),
.flogtanh( I1f97ea0e7bf46382824cbffc3e94e9df),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6b0d8c39fbd70231e5bf5c9b9690476b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1f97ea0e7bf46382824cbffc3e94e9df };
assign I79458089b042e181e37cc44c06d08681 = (Ifa8db43284d5bbebaed4f72d65cf9f92[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6b0d8c39fbd70231e5bf5c9b9690476b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00014_00001_U (
.flogtanh_sel( I365d9f3e8b2a9890427f07386deeb093[flogtanh_SEL-1:0]),
.flogtanh( I801dfe17655932ad8fe9702cbaad270f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie7241b933e5ad5520235b6af19caa8d5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I801dfe17655932ad8fe9702cbaad270f };
assign I42460fae0acff25fa2b829e39ddcc4fd = (I365d9f3e8b2a9890427f07386deeb093[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie7241b933e5ad5520235b6af19caa8d5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00014_00002_U (
.flogtanh_sel( I466aaa0b6cde2ade1901797b8c11e32c[flogtanh_SEL-1:0]),
.flogtanh( Idbd834f0c907b233a8eff58eaca28863),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2a3101f6f107fd42234971ee8ec79ad2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idbd834f0c907b233a8eff58eaca28863 };
assign Id3670a6f05d40ab69624544de92b9c64 = (I466aaa0b6cde2ade1901797b8c11e32c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2a3101f6f107fd42234971ee8ec79ad2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00014_00003_U (
.flogtanh_sel( I7057e329a65ab240ed6cfa824307af65[flogtanh_SEL-1:0]),
.flogtanh( Ic69e0c34630bde15f4172714bc3d92be),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibc273f3403da77770e246102b6aad94c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic69e0c34630bde15f4172714bc3d92be };
assign I81800fb49855a4fd2737faa07ff15d29 = (I7057e329a65ab240ed6cfa824307af65[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibc273f3403da77770e246102b6aad94c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00014_00004_U (
.flogtanh_sel( I624e50e3457d33d12680eaf8e7c34aa3[flogtanh_SEL-1:0]),
.flogtanh( I465a735c8e94ddbfdbaeb2a7652e481e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5a2febf5da7cbbb8bb0aee0830d8122e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I465a735c8e94ddbfdbaeb2a7652e481e };
assign Ibfe325e48511372569e0d98d9c4e70e3 = (I624e50e3457d33d12680eaf8e7c34aa3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5a2febf5da7cbbb8bb0aee0830d8122e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00015_00000_U (
.flogtanh_sel( I9f356fd6820c33fdb5baff05a781e192[flogtanh_SEL-1:0]),
.flogtanh( Id1c6a3f52dd7972f47cbd8103ace643f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I166fdc6588cbe080275b58ccae50fd80  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id1c6a3f52dd7972f47cbd8103ace643f };
assign I326660e98f61bb2ced4c23c7bcc9324a = (I9f356fd6820c33fdb5baff05a781e192[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I166fdc6588cbe080275b58ccae50fd80;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00015_00001_U (
.flogtanh_sel( I39b9c7c664fe7017731877d145d55b44[flogtanh_SEL-1:0]),
.flogtanh( I26b9e2d073b20376980662c249bf9d43),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifde315b0389f701a061b3f765cf35ce7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I26b9e2d073b20376980662c249bf9d43 };
assign Ic6fa98631d742b27f252fe7c95caef55 = (I39b9c7c664fe7017731877d145d55b44[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifde315b0389f701a061b3f765cf35ce7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00015_00002_U (
.flogtanh_sel( Ic62ffbb9e58e0d08b0dec24bba1dc6f2[flogtanh_SEL-1:0]),
.flogtanh( Id4cc1b15055941d401ded6ff8b777461),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0df682bffaf274789733b11506a1630f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id4cc1b15055941d401ded6ff8b777461 };
assign Iab6d0f72579687407e029c630b107f7d = (Ic62ffbb9e58e0d08b0dec24bba1dc6f2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0df682bffaf274789733b11506a1630f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00015_00003_U (
.flogtanh_sel( I8da2a532288fb817e7dc0cb7b4e3761c[flogtanh_SEL-1:0]),
.flogtanh( I064bd1f4b7fa40b2cae3ea361edf9167),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia39290e9e73e101284fb99f7aa472db4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I064bd1f4b7fa40b2cae3ea361edf9167 };
assign I19eae741ef89baa1a64c403fb29f14f4 = (I8da2a532288fb817e7dc0cb7b4e3761c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia39290e9e73e101284fb99f7aa472db4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00015_00004_U (
.flogtanh_sel( I6a6e559f5c98f846014e8107fea5a5d9[flogtanh_SEL-1:0]),
.flogtanh( I4b5aadc25b0ed6811a665b33d6c4ae2a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib4f9fe5e96247d914bbdcc12be4044a0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4b5aadc25b0ed6811a665b33d6c4ae2a };
assign I749b9c345f23aae03c595a2c76126ecb = (I6a6e559f5c98f846014e8107fea5a5d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib4f9fe5e96247d914bbdcc12be4044a0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00016_00000_U (
.flogtanh_sel( Ibef9219f577b1a62dfdd77296fbfb24d[flogtanh_SEL-1:0]),
.flogtanh( Ic883bcc70572a237ba0e3d465337bc59),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3b06a47b2157c79d4a63dc94865a43c8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic883bcc70572a237ba0e3d465337bc59 };
assign Idc77c7d5123717fc2596a51d904c6d82 = (Ibef9219f577b1a62dfdd77296fbfb24d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3b06a47b2157c79d4a63dc94865a43c8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00016_00001_U (
.flogtanh_sel( I52e6688b5bfff75529d18e20b22832ce[flogtanh_SEL-1:0]),
.flogtanh( I7181ab1d663b0cbe30861e29fc3f8532),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9f91a577741c480378c018f313c68030  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7181ab1d663b0cbe30861e29fc3f8532 };
assign I779da979707d9712c1626d6025f97599 = (I52e6688b5bfff75529d18e20b22832ce[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9f91a577741c480378c018f313c68030;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00016_00002_U (
.flogtanh_sel( Iff22c49354eefca0ea3c5959c14b782c[flogtanh_SEL-1:0]),
.flogtanh( Id3fbb6d083344684de89d99c040b2100),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9997a7033ca3806006f2706960325d6d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id3fbb6d083344684de89d99c040b2100 };
assign I97aede8502e443f98938487a5a5c072c = (Iff22c49354eefca0ea3c5959c14b782c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9997a7033ca3806006f2706960325d6d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00016_00003_U (
.flogtanh_sel( Ie5377bbdb4111ed00356d5b7737102f3[flogtanh_SEL-1:0]),
.flogtanh( Iee8d139aa5a8ae046f5019abecdbc3c4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0dea21c66fdec2b891938d4cfb4452cd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iee8d139aa5a8ae046f5019abecdbc3c4 };
assign Ie7820d1a242bc28c19ec32d2c91e47b7 = (Ie5377bbdb4111ed00356d5b7737102f3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0dea21c66fdec2b891938d4cfb4452cd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00016_00004_U (
.flogtanh_sel( I55bf0f3379a8c44634b8f0a3d06c049e[flogtanh_SEL-1:0]),
.flogtanh( Idc0bfe36a3a9b3006a04d5dfc31b8107),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia6e3665657bc28e92fa4ffb8ddcbc537  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idc0bfe36a3a9b3006a04d5dfc31b8107 };
assign I82a14e1ee4723e7d9a13c1f2b8b13691 = (I55bf0f3379a8c44634b8f0a3d06c049e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia6e3665657bc28e92fa4ffb8ddcbc537;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00017_00000_U (
.flogtanh_sel( I9bc9541607f4f6aedb686cdde297bcda[flogtanh_SEL-1:0]),
.flogtanh( Ia2462ec52aaccc97597d1dfc2e33b7e2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4097acfa6a9dbc9297745f4891286bd0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia2462ec52aaccc97597d1dfc2e33b7e2 };
assign I77a94cd9186ca546ca9664942ea3537f = (I9bc9541607f4f6aedb686cdde297bcda[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4097acfa6a9dbc9297745f4891286bd0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00017_00001_U (
.flogtanh_sel( Ia4620554fbb1d81a71a15a846e4be2f5[flogtanh_SEL-1:0]),
.flogtanh( I8048bbe27b49b9d248fee919be6dc977),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icef9faf2ee30e443183708bda55cf706  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8048bbe27b49b9d248fee919be6dc977 };
assign I3c0ddec25c53c166d30eb78d4518840e = (Ia4620554fbb1d81a71a15a846e4be2f5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icef9faf2ee30e443183708bda55cf706;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00017_00002_U (
.flogtanh_sel( Ibb31b35388ba8ba2ecf98449308ee67d[flogtanh_SEL-1:0]),
.flogtanh( I838d1cc5e9ca5058c25223ec53d9c34f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I68c9c1da797be9d6d1093884fef3ec3e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I838d1cc5e9ca5058c25223ec53d9c34f };
assign I98bbe3b75958f10195dee6460cf2aca6 = (Ibb31b35388ba8ba2ecf98449308ee67d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I68c9c1da797be9d6d1093884fef3ec3e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00017_00003_U (
.flogtanh_sel( Ia20410fb3d56587f89a54c00b943b305[flogtanh_SEL-1:0]),
.flogtanh( Id9e5147e089e6e52ef2a687d76534f16),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iff7f4a450dee1fe869764249a7a4e612  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id9e5147e089e6e52ef2a687d76534f16 };
assign If6d436031f68ef587750c5c1dfcfffc2 = (Ia20410fb3d56587f89a54c00b943b305[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iff7f4a450dee1fe869764249a7a4e612;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00017_00004_U (
.flogtanh_sel( I9d268f3da12e35b9a4229b7340c0f018[flogtanh_SEL-1:0]),
.flogtanh( Ia043941abbcf10c16f086fe8d61dd456),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I323b8c5e397420e5eb3c0872162dc013  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia043941abbcf10c16f086fe8d61dd456 };
assign I461398638cb8280f1779915298540b00 = (I9d268f3da12e35b9a4229b7340c0f018[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I323b8c5e397420e5eb3c0872162dc013;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00018_00000_U (
.flogtanh_sel( I2fce29bd666082eedb2fb3ec8b5ae4dd[flogtanh_SEL-1:0]),
.flogtanh( I625ab32380498dfbf9d3290c2053bf3d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib62e0c5c630f77706a8bc2ef1409214c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I625ab32380498dfbf9d3290c2053bf3d };
assign I20c65000bbc10299168af7390776a03c = (I2fce29bd666082eedb2fb3ec8b5ae4dd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib62e0c5c630f77706a8bc2ef1409214c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00018_00001_U (
.flogtanh_sel( Ia1e8b61e2579a90f5c88ded11c7322c2[flogtanh_SEL-1:0]),
.flogtanh( I903f7844e55d1cd6969352490c275c8e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id51115ce716fdb681e7d5d4cad1fa1c5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I903f7844e55d1cd6969352490c275c8e };
assign Ia840e19ca36795a50ab1a6e6a1729edb = (Ia1e8b61e2579a90f5c88ded11c7322c2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id51115ce716fdb681e7d5d4cad1fa1c5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00018_00002_U (
.flogtanh_sel( I8cf3718ba65b7fed72e3955f190e34d1[flogtanh_SEL-1:0]),
.flogtanh( Ie5951bc919195ba594fe87375ad41269),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifbb85fd268ca90f905cbe5587d34cbbb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie5951bc919195ba594fe87375ad41269 };
assign I7d98d1e5f07fccff5f20eaca6363c700 = (I8cf3718ba65b7fed72e3955f190e34d1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifbb85fd268ca90f905cbe5587d34cbbb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00018_00003_U (
.flogtanh_sel( I7e802d300af54d394b4ee041798c0513[flogtanh_SEL-1:0]),
.flogtanh( Ieeed8d4eebc0adea7ee0af6a5dbe045c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7e91bd3d8b70220941a7eb290852b898  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ieeed8d4eebc0adea7ee0af6a5dbe045c };
assign I97a75b8625ae2a143cf364790ae77753 = (I7e802d300af54d394b4ee041798c0513[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7e91bd3d8b70220941a7eb290852b898;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00018_00004_U (
.flogtanh_sel( Id4fd5a4b97cfa1e176a26f3a823c5516[flogtanh_SEL-1:0]),
.flogtanh( I266cd5f0a56cd5171da8d59df0042d5d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I366001777963d791fb7811c0fed5f268  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I266cd5f0a56cd5171da8d59df0042d5d };
assign Idbea892c8109117f90b453efe8ae25af = (Id4fd5a4b97cfa1e176a26f3a823c5516[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I366001777963d791fb7811c0fed5f268;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00019_00000_U (
.flogtanh_sel( Icbf8d4e75fc66c05eb49c5075696fb07[flogtanh_SEL-1:0]),
.flogtanh( Ie5a57c603ad520441bc5819c81fb877f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5db5b227fee3a0a53935d1fd86b1ec77  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie5a57c603ad520441bc5819c81fb877f };
assign Icfc1c6d96a3598af73e99a350c387d72 = (Icbf8d4e75fc66c05eb49c5075696fb07[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5db5b227fee3a0a53935d1fd86b1ec77;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00019_00001_U (
.flogtanh_sel( I746a7e90adb2f213b75ae12a161aca0d[flogtanh_SEL-1:0]),
.flogtanh( I17ac503f4f952f9e2fcdea3f955cc1a9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id9a0ece818dcc0a00e66ebc35c664c73  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I17ac503f4f952f9e2fcdea3f955cc1a9 };
assign I523e9b6f828ec7f166750112f8a3f676 = (I746a7e90adb2f213b75ae12a161aca0d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id9a0ece818dcc0a00e66ebc35c664c73;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00019_00002_U (
.flogtanh_sel( Icb1029aaaaed8c698862ea9c5e22132c[flogtanh_SEL-1:0]),
.flogtanh( Id8b704aada09411d5f5153d088c1c613),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I24326227bfacd8f0de4b746ba973242b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id8b704aada09411d5f5153d088c1c613 };
assign I79259217f63b2f6263552c434d0e5c93 = (Icb1029aaaaed8c698862ea9c5e22132c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I24326227bfacd8f0de4b746ba973242b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00019_00003_U (
.flogtanh_sel( Ib93ea7028c172373b53cdafecae32a67[flogtanh_SEL-1:0]),
.flogtanh( If64a200b2dac7049b77e5b6bb03b9cc3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic96744b0858aea49e052758e4efd4d8a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If64a200b2dac7049b77e5b6bb03b9cc3 };
assign Ice6db5ba70d3c7499df6723a2df56bfe = (Ib93ea7028c172373b53cdafecae32a67[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic96744b0858aea49e052758e4efd4d8a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00019_00004_U (
.flogtanh_sel( If9628275b000e418f3903daebfdace92[flogtanh_SEL-1:0]),
.flogtanh( Iee1b48cae01fe51344b8d662ace9c6f1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I98de4ec4bf1dc2402f1417c2d42a1e2f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iee1b48cae01fe51344b8d662ace9c6f1 };
assign I28aa517220bf597cf898660f698ef19d = (If9628275b000e418f3903daebfdace92[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I98de4ec4bf1dc2402f1417c2d42a1e2f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00000_U (
.flogtanh_sel( I830202fb6f08f98c7f71893a881bd555[flogtanh_SEL-1:0]),
.flogtanh( Ic879cd355d61eb021250d62841115a52),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1174526f0aeaaaaa3f10802ea73526f2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic879cd355d61eb021250d62841115a52 };
assign I07048dc5cbe24ff72d24902d572face0 = (I830202fb6f08f98c7f71893a881bd555[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1174526f0aeaaaaa3f10802ea73526f2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00001_U (
.flogtanh_sel( I6f38bc9359562f57c1603355e9ee312b[flogtanh_SEL-1:0]),
.flogtanh( I46e2d889b9ba7eccad5529200852ca17),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia49bff02824813d4823f50058348f4e1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I46e2d889b9ba7eccad5529200852ca17 };
assign Iab3876e5107e3a56b1fafe41e16d9482 = (I6f38bc9359562f57c1603355e9ee312b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia49bff02824813d4823f50058348f4e1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00002_U (
.flogtanh_sel( I4701b732d59c26e3790a63c1936f9a24[flogtanh_SEL-1:0]),
.flogtanh( Ia4e080f13520998be95b64eb883f8e32),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I30b6fe386734293d3541f1705a7e2f18  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia4e080f13520998be95b64eb883f8e32 };
assign I511a55c2f4d6d3727dff5825597f55a9 = (I4701b732d59c26e3790a63c1936f9a24[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I30b6fe386734293d3541f1705a7e2f18;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00003_U (
.flogtanh_sel( Ib5d28d8f73d17ab6df6a1291e50c04ab[flogtanh_SEL-1:0]),
.flogtanh( I2ad2ede07f1ffac643211e88bf8ddbd6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If7541af81460bd2457931a0f435716d8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2ad2ede07f1ffac643211e88bf8ddbd6 };
assign I2493237a24acdcab8b5bda10e804a5cf = (Ib5d28d8f73d17ab6df6a1291e50c04ab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If7541af81460bd2457931a0f435716d8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00004_U (
.flogtanh_sel( I81259f391db792339824ad5dd1a0057b[flogtanh_SEL-1:0]),
.flogtanh( I5bc390dc300be5f8bc85f928cca1cd0b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I47cd82d1a6107cbc86188bf1ff4a55a6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5bc390dc300be5f8bc85f928cca1cd0b };
assign I03829256e357ac17c7ca7cae2f980f41 = (I81259f391db792339824ad5dd1a0057b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I47cd82d1a6107cbc86188bf1ff4a55a6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00005_U (
.flogtanh_sel( I6f09ac63effe67a86798b9b4e1690664[flogtanh_SEL-1:0]),
.flogtanh( I3e7efaed64fd3c276e882ab38109d538),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I41f07d0c85ebaf33ef8dd9b96a438df2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3e7efaed64fd3c276e882ab38109d538 };
assign Iae32c44b88fe7ddb5d4f19cf8fff3ba6 = (I6f09ac63effe67a86798b9b4e1690664[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I41f07d0c85ebaf33ef8dd9b96a438df2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00006_U (
.flogtanh_sel( I370b4b3a0048a93ba374a40e170c75a3[flogtanh_SEL-1:0]),
.flogtanh( Ib4738fe629dbe40eefed821b40ab93c8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I95a440b3890f6d285bde57a8d879c9aa  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib4738fe629dbe40eefed821b40ab93c8 };
assign I3bdc5ba374f85dc61346e4868c41a6bf = (I370b4b3a0048a93ba374a40e170c75a3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I95a440b3890f6d285bde57a8d879c9aa;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00007_U (
.flogtanh_sel( I3f8476d0aa0ea2439b67ea1a4adf36c5[flogtanh_SEL-1:0]),
.flogtanh( I30268ed341753c3ab53b65ad43e94923),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2d3ee951489a62634a7b7332d5fd2450  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I30268ed341753c3ab53b65ad43e94923 };
assign I557ef77ce931535467a07a8d70145f55 = (I3f8476d0aa0ea2439b67ea1a4adf36c5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2d3ee951489a62634a7b7332d5fd2450;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00008_U (
.flogtanh_sel( I35b52dba10a8a5b22b518388fecac82d[flogtanh_SEL-1:0]),
.flogtanh( I2f10be9cbe2a935475077c0218031a5a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9f4acc72fd3769c7c300fc36aac958b3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2f10be9cbe2a935475077c0218031a5a };
assign Ib4695d4389db72c5ac7e31809072c290 = (I35b52dba10a8a5b22b518388fecac82d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9f4acc72fd3769c7c300fc36aac958b3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00009_U (
.flogtanh_sel( Ic7db274ed18e6fdecf30381a31238777[flogtanh_SEL-1:0]),
.flogtanh( I41d598b80334ab12e5f53b2a6c721517),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4de1d4373a309ecd3278d1891ddce050  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I41d598b80334ab12e5f53b2a6c721517 };
assign Ie81315a3a14a5ef879d8e3f405936365 = (Ic7db274ed18e6fdecf30381a31238777[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4de1d4373a309ecd3278d1891ddce050;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00010_U (
.flogtanh_sel( I2c4e538a8db759e9799541d9178ec61e[flogtanh_SEL-1:0]),
.flogtanh( I94b3d895ee69e3ab482ff1aa0798c92a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iea0a307bacf40b16646458e5e8ea6d9a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I94b3d895ee69e3ab482ff1aa0798c92a };
assign Ia7520053a7c4a94437c6a780b03a28a5 = (I2c4e538a8db759e9799541d9178ec61e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iea0a307bacf40b16646458e5e8ea6d9a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00011_U (
.flogtanh_sel( Ief6d4c3f5ef8663e111ef99347b023f5[flogtanh_SEL-1:0]),
.flogtanh( I24a25d4725db6bcb4732fa21bc861736),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id171f9ecb8da0298882ae2416c2132d3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I24a25d4725db6bcb4732fa21bc861736 };
assign Ic308a5413f38b96d244cac3b0bc9462c = (Ief6d4c3f5ef8663e111ef99347b023f5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id171f9ecb8da0298882ae2416c2132d3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00012_U (
.flogtanh_sel( Id95e964e5faecb52c72669b0d28a4bf5[flogtanh_SEL-1:0]),
.flogtanh( I1877b73e028c908de9dc734b93cbf8bb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic10ae3db593c8fb6a2d2a414b131dace  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1877b73e028c908de9dc734b93cbf8bb };
assign I034fb3850485fae2d1358041a1c41888 = (Id95e964e5faecb52c72669b0d28a4bf5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic10ae3db593c8fb6a2d2a414b131dace;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00020_00013_U (
.flogtanh_sel( I0fcef4538102ac6d24aa7090d5405afa[flogtanh_SEL-1:0]),
.flogtanh( Ic99b64430e5dfdabe3634fbddeb41b3c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9dd17bc57b2d75f3e50f2b2243ea6e0b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic99b64430e5dfdabe3634fbddeb41b3c };
assign I0e7079db66c15210046b997f319ece89 = (I0fcef4538102ac6d24aa7090d5405afa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9dd17bc57b2d75f3e50f2b2243ea6e0b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00000_U (
.flogtanh_sel( I055019e38eec6badd1739033d43d7d97[flogtanh_SEL-1:0]),
.flogtanh( I3c0ddec6d702a344930fd04f923bb2f1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I69c326b0728bef980588c914c3118d6f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3c0ddec6d702a344930fd04f923bb2f1 };
assign I9a5388f8aa6e9924a309aa8db4c1983b = (I055019e38eec6badd1739033d43d7d97[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I69c326b0728bef980588c914c3118d6f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00001_U (
.flogtanh_sel( I35c20a6e823da77a870b421eef2e0a95[flogtanh_SEL-1:0]),
.flogtanh( I41829e511abe1ddf9b67f899143db19a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I52e368d1bc43a02ad9418f54b3fe08b8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I41829e511abe1ddf9b67f899143db19a };
assign Ief76663994991118b1899ea4ddf4527d = (I35c20a6e823da77a870b421eef2e0a95[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I52e368d1bc43a02ad9418f54b3fe08b8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00002_U (
.flogtanh_sel( I32cc12cdacef1a4ef64577e0fa977f46[flogtanh_SEL-1:0]),
.flogtanh( I41961139f5b650e4f4ba5c2eadda6702),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I548594daa8f38ff594534dfa4d6238d9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I41961139f5b650e4f4ba5c2eadda6702 };
assign I6fb63ea54e492bdbc6d1145affc683e9 = (I32cc12cdacef1a4ef64577e0fa977f46[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I548594daa8f38ff594534dfa4d6238d9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00003_U (
.flogtanh_sel( I26b3f2360ca4a8caee61b2f3a3a08267[flogtanh_SEL-1:0]),
.flogtanh( I8ef0ac3bf43f16d2edf5a5045b0eb498),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1080d88996caef7f760f64532883ee93  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8ef0ac3bf43f16d2edf5a5045b0eb498 };
assign If83ce1cbe3a73472419520c225b288a6 = (I26b3f2360ca4a8caee61b2f3a3a08267[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1080d88996caef7f760f64532883ee93;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00004_U (
.flogtanh_sel( I5ef9b7dc0c63e9ca6a5fb5f7ffa06041[flogtanh_SEL-1:0]),
.flogtanh( I4084e3c9ba635fc4a8d281015bdeb33a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I49f6d04d31956a1134257027fabdb381  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4084e3c9ba635fc4a8d281015bdeb33a };
assign Id1df78ab32daf524b77c0431c782f2bf = (I5ef9b7dc0c63e9ca6a5fb5f7ffa06041[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I49f6d04d31956a1134257027fabdb381;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00005_U (
.flogtanh_sel( If881473b05090f40a027d7eeee7f7ed9[flogtanh_SEL-1:0]),
.flogtanh( I199a14038a0ff6ac25dab60162f8c6c9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2aacba8f2c989ba723b7f65c7c009c64  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I199a14038a0ff6ac25dab60162f8c6c9 };
assign Iff142b88493149045fc0de355b767c16 = (If881473b05090f40a027d7eeee7f7ed9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2aacba8f2c989ba723b7f65c7c009c64;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00006_U (
.flogtanh_sel( I23bd59ab5b038935301396aaf2acefc1[flogtanh_SEL-1:0]),
.flogtanh( Ic6859263f79d29d5f4896d85367be2bf),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If0cf7facd593ca5190b2e20429c1868a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic6859263f79d29d5f4896d85367be2bf };
assign I28c3818247c7c6de11790f6692882b5a = (I23bd59ab5b038935301396aaf2acefc1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If0cf7facd593ca5190b2e20429c1868a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00007_U (
.flogtanh_sel( I874386d94dacf84e699d159af1a49836[flogtanh_SEL-1:0]),
.flogtanh( If0af3259e321390fffe518318f0f2545),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I40d7acfc8d14404d3669e04dbfd61659  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If0af3259e321390fffe518318f0f2545 };
assign Ib451127b69a0a800332a712af77c6d29 = (I874386d94dacf84e699d159af1a49836[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I40d7acfc8d14404d3669e04dbfd61659;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00008_U (
.flogtanh_sel( I95bfe51a759bf4165168e5e3b99d6b34[flogtanh_SEL-1:0]),
.flogtanh( Icafbf36da24f4db99e0ce4eeca6ca338),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I43e5964e737fd1bf55c876d36d1a573d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icafbf36da24f4db99e0ce4eeca6ca338 };
assign I3d601db540da359ae4d22f960d3d5af8 = (I95bfe51a759bf4165168e5e3b99d6b34[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I43e5964e737fd1bf55c876d36d1a573d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00009_U (
.flogtanh_sel( I4ba5b2f9b7ec0937ecd2c9945cf6de87[flogtanh_SEL-1:0]),
.flogtanh( Ia614303d31afc0ef4f15ec5b43231cd8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I85cc34b35ec9a6e377263bc8307ae9af  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia614303d31afc0ef4f15ec5b43231cd8 };
assign I2c1f2476efe593829ade470fe8ec2526 = (I4ba5b2f9b7ec0937ecd2c9945cf6de87[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I85cc34b35ec9a6e377263bc8307ae9af;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00010_U (
.flogtanh_sel( I0b08fb8db0e8a1de3d416907c87fe700[flogtanh_SEL-1:0]),
.flogtanh( I28ff2f86da2016b00bd0c21cbd1b4530),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0bf108b578bd4decc8b7b8d9db13d4a1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I28ff2f86da2016b00bd0c21cbd1b4530 };
assign I7e685b06df8a8c2ac351fa9f9b76a81d = (I0b08fb8db0e8a1de3d416907c87fe700[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0bf108b578bd4decc8b7b8d9db13d4a1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00011_U (
.flogtanh_sel( Ie030d12e5acf9ef4975a17c83b2481c1[flogtanh_SEL-1:0]),
.flogtanh( I2b8c969c11b4117c96470f4f6ed6963a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idcd92c1ab555e9586c17b939903bc6a1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2b8c969c11b4117c96470f4f6ed6963a };
assign I1338d211b5d2d409bfe0df76d2ca2701 = (Ie030d12e5acf9ef4975a17c83b2481c1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idcd92c1ab555e9586c17b939903bc6a1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00012_U (
.flogtanh_sel( Ia7a0e852d3dfcef950804ea0ebb0c80a[flogtanh_SEL-1:0]),
.flogtanh( Iea563639beb7fcb0291b5dc1410951d1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I45f165607aba91f1026657ea9c265bb7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iea563639beb7fcb0291b5dc1410951d1 };
assign Ia40dad546d9c852e2fa8942c62a1c1f8 = (Ia7a0e852d3dfcef950804ea0ebb0c80a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I45f165607aba91f1026657ea9c265bb7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00021_00013_U (
.flogtanh_sel( Iaa4c38d030eab2b7899399aa0d7886d9[flogtanh_SEL-1:0]),
.flogtanh( Ic1b35046657e23f42199e39343a652a8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If6a9b9c0cff23cab0ac2af86f2eab66a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic1b35046657e23f42199e39343a652a8 };
assign I0b0dd019d8bd24684403a29aed668b6d = (Iaa4c38d030eab2b7899399aa0d7886d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If6a9b9c0cff23cab0ac2af86f2eab66a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00000_U (
.flogtanh_sel( Icce7ff1d652d4d9c2be5ecf679059bbe[flogtanh_SEL-1:0]),
.flogtanh( Ie7b26120ee77b43574c1ca171d7ec15f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5f36159573f16b76a28cca6923881ece  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie7b26120ee77b43574c1ca171d7ec15f };
assign I66a304016a9adfd85a2abb6f8fd39afc = (Icce7ff1d652d4d9c2be5ecf679059bbe[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5f36159573f16b76a28cca6923881ece;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00001_U (
.flogtanh_sel( If816bc5eacaea23443602e575ddf60b8[flogtanh_SEL-1:0]),
.flogtanh( I2ed61ced1577d905da91d97592006ed5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icd396e938ee702fab0f788a7a91b90cf  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2ed61ced1577d905da91d97592006ed5 };
assign I177be24718c59688752097fe2a4085c4 = (If816bc5eacaea23443602e575ddf60b8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icd396e938ee702fab0f788a7a91b90cf;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00002_U (
.flogtanh_sel( I3b224a4ded05446cc5300d430bdd1947[flogtanh_SEL-1:0]),
.flogtanh( I332dc26a52194745d19c4d8468e42864),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6cee7c45f29f8e1affd935a441d8a0a7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I332dc26a52194745d19c4d8468e42864 };
assign I7e66a42eb7cdb820cd1297c39f0625e8 = (I3b224a4ded05446cc5300d430bdd1947[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6cee7c45f29f8e1affd935a441d8a0a7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00003_U (
.flogtanh_sel( Ia5fc5cfb0e52237b407b37a3858fccb5[flogtanh_SEL-1:0]),
.flogtanh( Ibb4fefe05e94e055e86a743c40fb1c5e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7d389f1dba81f9205521753c52490695  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibb4fefe05e94e055e86a743c40fb1c5e };
assign If2021f0735c6c5649ebac0d230fda87c = (Ia5fc5cfb0e52237b407b37a3858fccb5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7d389f1dba81f9205521753c52490695;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00004_U (
.flogtanh_sel( I92f8ba6e7f8e9b30fb5b6973eb8fd03e[flogtanh_SEL-1:0]),
.flogtanh( Ia56a76a20d4f11b0e80cbe31820a6977),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I759d027d500e4bf950a89c0a49e135c3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia56a76a20d4f11b0e80cbe31820a6977 };
assign Ie1bf5d97b8f679095d2442bbf9f95608 = (I92f8ba6e7f8e9b30fb5b6973eb8fd03e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I759d027d500e4bf950a89c0a49e135c3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00005_U (
.flogtanh_sel( Icdfa60d2a024dd934f7e6639c6cb2c28[flogtanh_SEL-1:0]),
.flogtanh( I054ebc7f9e3da325ba0c6e329f2ee770),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I378871e4d07eabcf01ff30c299f8f054  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I054ebc7f9e3da325ba0c6e329f2ee770 };
assign I632469889d6bb1c268b45fb805467ebd = (Icdfa60d2a024dd934f7e6639c6cb2c28[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I378871e4d07eabcf01ff30c299f8f054;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00006_U (
.flogtanh_sel( Ifff70b976513eaa42b6bd4b80c98611e[flogtanh_SEL-1:0]),
.flogtanh( I3361df26cc86ca8be1653d9376d0c8e0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id346411c557c6ac494ab4913a44c6cf0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3361df26cc86ca8be1653d9376d0c8e0 };
assign Ie230ba3c73808e102eee9e5868595e7c = (Ifff70b976513eaa42b6bd4b80c98611e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id346411c557c6ac494ab4913a44c6cf0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00007_U (
.flogtanh_sel( Ica12fa8b631b70a6bbe9f6e92bf73ea0[flogtanh_SEL-1:0]),
.flogtanh( I586fbde80f0130c4a6ead49de11efdd9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2ed644da3d2a47eef5788a3139de04ac  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I586fbde80f0130c4a6ead49de11efdd9 };
assign Ie1e9326e4eee006ec07abb6bb7d269a5 = (Ica12fa8b631b70a6bbe9f6e92bf73ea0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2ed644da3d2a47eef5788a3139de04ac;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00008_U (
.flogtanh_sel( Ie69c255335760f706c644b115887269b[flogtanh_SEL-1:0]),
.flogtanh( Ifa087137c8a6028b13bfa95aba19fc34),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6e90f86b20562e80e2935d1886123672  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifa087137c8a6028b13bfa95aba19fc34 };
assign Ica4ec1647bdb5a3aad6db6b447bd7995 = (Ie69c255335760f706c644b115887269b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6e90f86b20562e80e2935d1886123672;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00009_U (
.flogtanh_sel( Idb06676b41de19bc86eae34c292183d9[flogtanh_SEL-1:0]),
.flogtanh( I51a3a6c79c488c092394375891775be3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5c8c09dcb6623c9dee9772f1409ffc98  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I51a3a6c79c488c092394375891775be3 };
assign Ia17295aec0a40c2b46a595dacfede2d5 = (Idb06676b41de19bc86eae34c292183d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5c8c09dcb6623c9dee9772f1409ffc98;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00010_U (
.flogtanh_sel( Ib21d2306d5ded3406fac754e69a10d20[flogtanh_SEL-1:0]),
.flogtanh( I01a7ebdc760227ee40b85828e28238a9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6bbd4143192116282eab3d7fbcb544e6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I01a7ebdc760227ee40b85828e28238a9 };
assign I4c6d3d6fc2d10066a744fdd9405a7902 = (Ib21d2306d5ded3406fac754e69a10d20[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6bbd4143192116282eab3d7fbcb544e6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00011_U (
.flogtanh_sel( Ib41d1aa2dcf81879976fb8964cbf6f79[flogtanh_SEL-1:0]),
.flogtanh( Ib3f9e4c05e363069775e5de9d240b3dc),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5177a497f9d6aae2f1917987542472f0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib3f9e4c05e363069775e5de9d240b3dc };
assign Ia9c043c5e8873fd13e39cf6bd8136c51 = (Ib41d1aa2dcf81879976fb8964cbf6f79[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5177a497f9d6aae2f1917987542472f0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00012_U (
.flogtanh_sel( I5f8f5e246f008b8d8c75f72828337bab[flogtanh_SEL-1:0]),
.flogtanh( I18664482dcc1371fa4b915af96070539),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7cdb256503fb49f4bc9123c0815ea3dd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I18664482dcc1371fa4b915af96070539 };
assign I2e802c75c6ce34b05943b678ecbfacb1 = (I5f8f5e246f008b8d8c75f72828337bab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7cdb256503fb49f4bc9123c0815ea3dd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00022_00013_U (
.flogtanh_sel( Id6625e78da0e14d2eeb19cc8ac6520e0[flogtanh_SEL-1:0]),
.flogtanh( I6a41c6cf78cb25ad1c47550756449002),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia116be2c3a094f1f5e1d04db21123309  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6a41c6cf78cb25ad1c47550756449002 };
assign Ieb3f28762410fb40a0c8a8556b4b3ca0 = (Id6625e78da0e14d2eeb19cc8ac6520e0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia116be2c3a094f1f5e1d04db21123309;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00000_U (
.flogtanh_sel( I6d9ddc6afa559ac35c042df1a9390ce9[flogtanh_SEL-1:0]),
.flogtanh( Iaf660a97d66e0d7f8e26f65229b7683f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I75175fd0c716e6fbc022cbbd73a9fefd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iaf660a97d66e0d7f8e26f65229b7683f };
assign Ie3e0c0e40c7a67ce7f957e74bd2a895d = (I6d9ddc6afa559ac35c042df1a9390ce9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I75175fd0c716e6fbc022cbbd73a9fefd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00001_U (
.flogtanh_sel( I9334055c7833676469670372d3c5cc31[flogtanh_SEL-1:0]),
.flogtanh( I7ded197ff64af1bce0e0d85705900a42),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I31809c8a10f68b5058f8db1db8d2f714  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7ded197ff64af1bce0e0d85705900a42 };
assign I491f2373b2df19a4c22e1787ef034179 = (I9334055c7833676469670372d3c5cc31[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I31809c8a10f68b5058f8db1db8d2f714;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00002_U (
.flogtanh_sel( I0c97d772c737c6ff85b584bf69ccaf93[flogtanh_SEL-1:0]),
.flogtanh( I7c06179d5424165f8a805754834fd98c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9f4163bac1b52f4282b51e6767085f7f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7c06179d5424165f8a805754834fd98c };
assign Ief96603d41b4f670d2bbfa3d3875c903 = (I0c97d772c737c6ff85b584bf69ccaf93[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9f4163bac1b52f4282b51e6767085f7f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00003_U (
.flogtanh_sel( Ic6ce97ae85d91dd8a79f3f9d0da375a2[flogtanh_SEL-1:0]),
.flogtanh( Id364f2a517a0f3109564a025ffd8eec3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iccc62d273c738111d4ec9adea8c3aec8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id364f2a517a0f3109564a025ffd8eec3 };
assign I7a029c27d92754041eb6d605837238dd = (Ic6ce97ae85d91dd8a79f3f9d0da375a2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iccc62d273c738111d4ec9adea8c3aec8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00004_U (
.flogtanh_sel( I83ff9a2750b298b0f7c9b6ce13f574af[flogtanh_SEL-1:0]),
.flogtanh( Ie3ea12584ed3e255073776620d778f06),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0c15c6d14710a00728d755472f83d8aa  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie3ea12584ed3e255073776620d778f06 };
assign I00dad36628d2fa923120fdaa79bf0045 = (I83ff9a2750b298b0f7c9b6ce13f574af[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0c15c6d14710a00728d755472f83d8aa;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00005_U (
.flogtanh_sel( I85699a2a05c343a6a9e828af6d445e9e[flogtanh_SEL-1:0]),
.flogtanh( I38d885c58b4f7333c679b0b5783418df),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5a1afe8d872b05da9e7eb44dd4bafb9f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I38d885c58b4f7333c679b0b5783418df };
assign I3707f68de059df0af5c652fc0478e543 = (I85699a2a05c343a6a9e828af6d445e9e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5a1afe8d872b05da9e7eb44dd4bafb9f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00006_U (
.flogtanh_sel( I51f6e39b24b2554884e381be79f47ff2[flogtanh_SEL-1:0]),
.flogtanh( I69251440f80eb2e177307aec4cb0111f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If40a1a450ba33087149fb6cdcf1f202e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I69251440f80eb2e177307aec4cb0111f };
assign I94af4b6b9dc11935db54ba872889392d = (I51f6e39b24b2554884e381be79f47ff2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If40a1a450ba33087149fb6cdcf1f202e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00007_U (
.flogtanh_sel( I9f65fd05c6929300860c8cbbde5607f2[flogtanh_SEL-1:0]),
.flogtanh( I0a9bcd4a3b79b003b5df8afa0d6b6782),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7079b578409c284713f6b1045c34b659  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0a9bcd4a3b79b003b5df8afa0d6b6782 };
assign I38e2dbba093928b874d447362d89b291 = (I9f65fd05c6929300860c8cbbde5607f2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7079b578409c284713f6b1045c34b659;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00008_U (
.flogtanh_sel( If09761d8f06051d4287ee29ac9c9fa19[flogtanh_SEL-1:0]),
.flogtanh( I36569656996bf98bce33b2d7a4b79def),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I336b37e04a2d76a541fcb62871e0c9d4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I36569656996bf98bce33b2d7a4b79def };
assign Ia48f0029e9e76386f3dd70aacd9adbfa = (If09761d8f06051d4287ee29ac9c9fa19[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I336b37e04a2d76a541fcb62871e0c9d4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00009_U (
.flogtanh_sel( I33bfbe0bcca6d32c86b9576577e3f265[flogtanh_SEL-1:0]),
.flogtanh( I7e408a50d0511909aeb57d5a00535e80),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I82325e0f7a4aa9849d619e8b8617c9b8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7e408a50d0511909aeb57d5a00535e80 };
assign Ic2b20168744fafbe15037ed7fa83da72 = (I33bfbe0bcca6d32c86b9576577e3f265[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I82325e0f7a4aa9849d619e8b8617c9b8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00010_U (
.flogtanh_sel( If2921210b1c05ecbf00af3a2bcb96ef4[flogtanh_SEL-1:0]),
.flogtanh( Iacc6f48dd92dc515be06a681cc5b56e9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8bf35575b614154bed06e946d5daf9eb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iacc6f48dd92dc515be06a681cc5b56e9 };
assign I62fdc8936121a2707d94cf3bd6e660ac = (If2921210b1c05ecbf00af3a2bcb96ef4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8bf35575b614154bed06e946d5daf9eb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00011_U (
.flogtanh_sel( Ib074e38e280474a782da831a3e0028b4[flogtanh_SEL-1:0]),
.flogtanh( Icafa051878ad3421c31ed2550ea09945),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If13d0317f786afef5e7dbbb9d4cd241a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icafa051878ad3421c31ed2550ea09945 };
assign Ia0932b3fd6a5ae6da2bacd2b86ba3a43 = (Ib074e38e280474a782da831a3e0028b4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If13d0317f786afef5e7dbbb9d4cd241a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00012_U (
.flogtanh_sel( I507449dde0bc0c8f53a10759436ec731[flogtanh_SEL-1:0]),
.flogtanh( If4e4f2776b1467e4f03bf15ff5f43c04),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6caaf723f09fdfc7684e94af6fd94d30  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If4e4f2776b1467e4f03bf15ff5f43c04 };
assign I9fce6091885f1bb97d29fb1f543b1a38 = (I507449dde0bc0c8f53a10759436ec731[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6caaf723f09fdfc7684e94af6fd94d30;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00023_00013_U (
.flogtanh_sel( Id55a3e3f2d75baeba71a345fad695c69[flogtanh_SEL-1:0]),
.flogtanh( I9387cd07e38260005bb3e41807d2d794),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3925ce727ac5b2dfff6a5982d034eb80  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9387cd07e38260005bb3e41807d2d794 };
assign Ib402cdbfaa9900820b85bd625415c547 = (Id55a3e3f2d75baeba71a345fad695c69[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3925ce727ac5b2dfff6a5982d034eb80;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00024_00000_U (
.flogtanh_sel( I20984f43d22671639a7a178ad15aec04[flogtanh_SEL-1:0]),
.flogtanh( I8bede290f421e6a05e49244f0d1d3d9b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3b949d926e8052d319c9262a80951516  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8bede290f421e6a05e49244f0d1d3d9b };
assign I518a2736384c14c02f27bfa3d8ea7aff = (I20984f43d22671639a7a178ad15aec04[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3b949d926e8052d319c9262a80951516;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00024_00001_U (
.flogtanh_sel( I59f88336d6bdd50ded87d353fb5ce3e9[flogtanh_SEL-1:0]),
.flogtanh( I6d8c2489fdeb42411f2e12bfa30752d2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7e8e247667ba53ee311f29a82574c0b7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6d8c2489fdeb42411f2e12bfa30752d2 };
assign I847cf7ff866f8a666872c12d6b67b1b1 = (I59f88336d6bdd50ded87d353fb5ce3e9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7e8e247667ba53ee311f29a82574c0b7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00024_00002_U (
.flogtanh_sel( I488635e3f7ed77ea88199f5bffd4b1d6[flogtanh_SEL-1:0]),
.flogtanh( I082715d1b8943faf11d464087542a83e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If6264b63f2c37286744ad61d579d2cc7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I082715d1b8943faf11d464087542a83e };
assign I9e45e3d7117ce48cdbfc5db8c0ccfcf4 = (I488635e3f7ed77ea88199f5bffd4b1d6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If6264b63f2c37286744ad61d579d2cc7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00024_00003_U (
.flogtanh_sel( Ie6893017d21c050ba10d206854f4a9f4[flogtanh_SEL-1:0]),
.flogtanh( I4de91d9613edc5c4d096b717d9df5de4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I71f47913679ccca9ab806c95c1152182  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4de91d9613edc5c4d096b717d9df5de4 };
assign I380ff8528cdba4026fac3c4eda8b2c52 = (Ie6893017d21c050ba10d206854f4a9f4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I71f47913679ccca9ab806c95c1152182;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00024_00004_U (
.flogtanh_sel( Id3f68b4dc0ab60673208b7d2081f3533[flogtanh_SEL-1:0]),
.flogtanh( Ifb2a91a74b87c75592cb046b9bfd9c8b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7b8e7702e50151938e6bb4bcfe59bcad  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifb2a91a74b87c75592cb046b9bfd9c8b };
assign Iee8f9b0654f6f6797f11cae0947e454e = (Id3f68b4dc0ab60673208b7d2081f3533[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7b8e7702e50151938e6bb4bcfe59bcad;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00024_00005_U (
.flogtanh_sel( I433756b944e061a824a89bda241e879f[flogtanh_SEL-1:0]),
.flogtanh( Ie21cffaecd7fe37601dcaef49a0d6cc3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic7799445f86a0bb5bed7a74ebe2531fd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie21cffaecd7fe37601dcaef49a0d6cc3 };
assign Ie3e54a4700d8d0f6478187e06cb6f85d = (I433756b944e061a824a89bda241e879f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic7799445f86a0bb5bed7a74ebe2531fd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00024_00006_U (
.flogtanh_sel( I2eb60a922aa4f7482dd92b9351d53a2d[flogtanh_SEL-1:0]),
.flogtanh( Ia648c9d395ad2727209229807b4224fb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic09ec6636c2f6157512550bfe533ac03  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia648c9d395ad2727209229807b4224fb };
assign I8c0069e8756bcff203ce21ae3170aa42 = (I2eb60a922aa4f7482dd92b9351d53a2d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic09ec6636c2f6157512550bfe533ac03;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00025_00000_U (
.flogtanh_sel( I0867979e1b159c8ceae548930376f482[flogtanh_SEL-1:0]),
.flogtanh( Ib415da845b88e5a8261beaf88b7ec804),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I93edc232c5754d21318c71402ba15dad  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib415da845b88e5a8261beaf88b7ec804 };
assign I856eada207c5006beb8f83f01d5d74c9 = (I0867979e1b159c8ceae548930376f482[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I93edc232c5754d21318c71402ba15dad;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00025_00001_U (
.flogtanh_sel( I4accfbeae8a5ee0dbeab23ef3a116145[flogtanh_SEL-1:0]),
.flogtanh( I6dffcf934a74385aa716db9d7fa29ed1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8af3fc54adca45e7dbf26e3bd793cd7b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6dffcf934a74385aa716db9d7fa29ed1 };
assign I79a46279070c53678a5af54f661c5821 = (I4accfbeae8a5ee0dbeab23ef3a116145[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8af3fc54adca45e7dbf26e3bd793cd7b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00025_00002_U (
.flogtanh_sel( Ic7570b0b7c5bef5758f68562ae4c90f6[flogtanh_SEL-1:0]),
.flogtanh( I13383df545ed8620a17a4fc2493cd770),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If111e57b5685180f787cc00a5ca98c39  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I13383df545ed8620a17a4fc2493cd770 };
assign Ica807adc510a2e32580ca77c18ea0b45 = (Ic7570b0b7c5bef5758f68562ae4c90f6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If111e57b5685180f787cc00a5ca98c39;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00025_00003_U (
.flogtanh_sel( Iceadadc4456881fdeea85934a9bf4d6c[flogtanh_SEL-1:0]),
.flogtanh( I87ea43bfae8fad4e4c26741fd2de5b41),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I13886c8ae8cffd0b01f2f3ce76fbe755  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I87ea43bfae8fad4e4c26741fd2de5b41 };
assign Ia8094903aed8dd0ce8e9ff459a5287b0 = (Iceadadc4456881fdeea85934a9bf4d6c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I13886c8ae8cffd0b01f2f3ce76fbe755;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00025_00004_U (
.flogtanh_sel( I7b2b617ae67424f54961eebce42de77e[flogtanh_SEL-1:0]),
.flogtanh( I6d2022ba184980b8e5bc5edb4f4b0ff3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id2e58c1480df3e5cadf231bbd03aaf8e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6d2022ba184980b8e5bc5edb4f4b0ff3 };
assign Ie018f3003c5f124bddd13c359257bf35 = (I7b2b617ae67424f54961eebce42de77e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id2e58c1480df3e5cadf231bbd03aaf8e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00025_00005_U (
.flogtanh_sel( I953f0f8af76f89b2d9ab4abf19fb411d[flogtanh_SEL-1:0]),
.flogtanh( I68f98b68c9a3836d0c7dc152a2d441da),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5fbf6c0b386eb14a493c94824ba51dea  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I68f98b68c9a3836d0c7dc152a2d441da };
assign Ice18bceb10fec484ffc96155e14c4974 = (I953f0f8af76f89b2d9ab4abf19fb411d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5fbf6c0b386eb14a493c94824ba51dea;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00025_00006_U (
.flogtanh_sel( I915b4736dcb20f831d02e48f4e79f008[flogtanh_SEL-1:0]),
.flogtanh( I2dc3cec85c37aa943f01df545f952e05),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8a77a7011da9a8d0a14e561b73d7df86  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2dc3cec85c37aa943f01df545f952e05 };
assign Ib484aa64b795f7e36198b800f302164f = (I915b4736dcb20f831d02e48f4e79f008[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8a77a7011da9a8d0a14e561b73d7df86;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00026_00000_U (
.flogtanh_sel( Ib7eec587348ae1ca1f00c0a3ad10ad27[flogtanh_SEL-1:0]),
.flogtanh( Ieed49c262f87c86b30d94e9842525ab0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifa70dba64cfba1806028839643ea900b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ieed49c262f87c86b30d94e9842525ab0 };
assign Icdb143a4ce96029c2441758bf2edd7b0 = (Ib7eec587348ae1ca1f00c0a3ad10ad27[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifa70dba64cfba1806028839643ea900b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00026_00001_U (
.flogtanh_sel( I001a212686304248c8359e5fc01227c0[flogtanh_SEL-1:0]),
.flogtanh( Ib9ab475010c98fc4e06df5c98944387a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If81b9c6cecfb4f03c642cf8ad899833a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib9ab475010c98fc4e06df5c98944387a };
assign I3a76f70ca3bfbcacc6f3342aa71f1912 = (I001a212686304248c8359e5fc01227c0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If81b9c6cecfb4f03c642cf8ad899833a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00026_00002_U (
.flogtanh_sel( Ibb7554e012c0fc1223c29b759c900666[flogtanh_SEL-1:0]),
.flogtanh( If7c8bdd5bae4a1bffd4bd2c8015bb738),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia515c4910fdd7af0fbf81e2094be54e0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If7c8bdd5bae4a1bffd4bd2c8015bb738 };
assign I9470c7ab9634c01bb832c9e4ff5496bf = (Ibb7554e012c0fc1223c29b759c900666[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia515c4910fdd7af0fbf81e2094be54e0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00026_00003_U (
.flogtanh_sel( I9aeb9c42b54a05be6bf9b7b88b6860ba[flogtanh_SEL-1:0]),
.flogtanh( I6463249144cd032e1c5af9e2987254b3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic110a8375139cd038f6fad5631ff6df6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6463249144cd032e1c5af9e2987254b3 };
assign I218ee96418a4f5d734d3d71685bc09c7 = (I9aeb9c42b54a05be6bf9b7b88b6860ba[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic110a8375139cd038f6fad5631ff6df6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00026_00004_U (
.flogtanh_sel( I6a5a5966965b0790b906c6fda71aef80[flogtanh_SEL-1:0]),
.flogtanh( I5f9e468fc1bc199574d719d866d52dfc),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5b1da643c42d2bf15855112416b6ee01  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5f9e468fc1bc199574d719d866d52dfc };
assign I924514226fdb5bac110a2650bcb2e85f = (I6a5a5966965b0790b906c6fda71aef80[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5b1da643c42d2bf15855112416b6ee01;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00026_00005_U (
.flogtanh_sel( Ic943083ca65ace6c42d73f4234739a06[flogtanh_SEL-1:0]),
.flogtanh( Ie69f792c606c3162052840dec732ef99),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iefe55f571684afc7c5257ae145de8594  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie69f792c606c3162052840dec732ef99 };
assign Idc57f37015a48393608e2b026bc7065c = (Ic943083ca65ace6c42d73f4234739a06[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iefe55f571684afc7c5257ae145de8594;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00026_00006_U (
.flogtanh_sel( Id0b321686d4c39621024cf0dd99822dc[flogtanh_SEL-1:0]),
.flogtanh( If874254c3c6813ff0d5184b574cb613d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7195c3cd02b5b61f50217c41cd409cf6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If874254c3c6813ff0d5184b574cb613d };
assign I41af7e4c97fc04154fe6de66b82499f5 = (Id0b321686d4c39621024cf0dd99822dc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7195c3cd02b5b61f50217c41cd409cf6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00027_00000_U (
.flogtanh_sel( I0839dd3787442f1b79b87e02436bfdce[flogtanh_SEL-1:0]),
.flogtanh( I90969c917df8480d379afef834c1a253),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I39f71f309736112e18565c8a18bc594a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I90969c917df8480d379afef834c1a253 };
assign I972bee4216f8e532e8fa4bd25fbb9c57 = (I0839dd3787442f1b79b87e02436bfdce[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I39f71f309736112e18565c8a18bc594a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00027_00001_U (
.flogtanh_sel( I89e6a9fd97d8aa4dd3b832c3be4697b2[flogtanh_SEL-1:0]),
.flogtanh( I07280ae3417855f994980fbb95696fc6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4fb6ab2aea28cb0776f52fc291782a27  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I07280ae3417855f994980fbb95696fc6 };
assign Ib303ea0240e7ab5f000dd10e975b2274 = (I89e6a9fd97d8aa4dd3b832c3be4697b2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4fb6ab2aea28cb0776f52fc291782a27;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00027_00002_U (
.flogtanh_sel( I93d4157f48b132642752220059861e98[flogtanh_SEL-1:0]),
.flogtanh( I852c62fffff0fd7bf06939d75fada3eb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I85d1c9d05f286204503b33dc9417c3f4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I852c62fffff0fd7bf06939d75fada3eb };
assign I5971253546899e9a82f387d5eabcc7b3 = (I93d4157f48b132642752220059861e98[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I85d1c9d05f286204503b33dc9417c3f4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00027_00003_U (
.flogtanh_sel( I8fc4faa2891d7fd3479ac1f788f481dc[flogtanh_SEL-1:0]),
.flogtanh( I9e0a2da5a82f1b509bd502554f4760aa),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8827c931edb38391e37eca5443c0f26a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9e0a2da5a82f1b509bd502554f4760aa };
assign I1fc36e6f738fab96df356979e1e3a612 = (I8fc4faa2891d7fd3479ac1f788f481dc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8827c931edb38391e37eca5443c0f26a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00027_00004_U (
.flogtanh_sel( I440f30e9cb4bc89233b46ea00b4cbeb4[flogtanh_SEL-1:0]),
.flogtanh( I6293c2b405087f14b42b423336f6990c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I495c79f2d8ec79a2f03613e0b64bde0e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6293c2b405087f14b42b423336f6990c };
assign Ie2d8c84d8c9a4c8f637068a2ae39fdde = (I440f30e9cb4bc89233b46ea00b4cbeb4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I495c79f2d8ec79a2f03613e0b64bde0e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00027_00005_U (
.flogtanh_sel( I6568bfd8780c11e0b1b049a01f92abd8[flogtanh_SEL-1:0]),
.flogtanh( I70e8d96970e69bc828a6aea5ade3bdd1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I954c51f604d6b8e7557797dd06aec9b7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I70e8d96970e69bc828a6aea5ade3bdd1 };
assign I114c595caa67a3f777f087a634130a6d = (I6568bfd8780c11e0b1b049a01f92abd8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I954c51f604d6b8e7557797dd06aec9b7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00027_00006_U (
.flogtanh_sel( Ibf7dc4da07f9955d5d4c7e1f63f1ad68[flogtanh_SEL-1:0]),
.flogtanh( I0380003f741eedb994793c2cb7e6c5c3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icd91fad15b5b5844144ac5c34218955f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0380003f741eedb994793c2cb7e6c5c3 };
assign Idad14b6383b9af54eb35e72ff3d10035 = (Ibf7dc4da07f9955d5d4c7e1f63f1ad68[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icd91fad15b5b5844144ac5c34218955f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00000_U (
.flogtanh_sel( I7ec1a328587b72a39c462083efea0ee0[flogtanh_SEL-1:0]),
.flogtanh( Ia884fcfa49cfe0b404bf49b99d7381aa),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4caf7dc4da499ea51928aa11326e0eae  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia884fcfa49cfe0b404bf49b99d7381aa };
assign I46e9c76b19ed1ff21f102efe6ee5c732 = (I7ec1a328587b72a39c462083efea0ee0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4caf7dc4da499ea51928aa11326e0eae;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00001_U (
.flogtanh_sel( Iaf028e7ab4dc77a7649f15d603834b5f[flogtanh_SEL-1:0]),
.flogtanh( Ie4ecd4c122ea5b478f3d7d2d632b8bf4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5461e1657c752f83cca50253e1db6772  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie4ecd4c122ea5b478f3d7d2d632b8bf4 };
assign Ic75b8bbb1b80001ec188a0cd25623420 = (Iaf028e7ab4dc77a7649f15d603834b5f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5461e1657c752f83cca50253e1db6772;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00002_U (
.flogtanh_sel( I58db79a8e9f0cd1ded379897ba2f27ae[flogtanh_SEL-1:0]),
.flogtanh( I82e534ecaabf5af6a9b6a567b862800a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib184e1d3a451b69a5206cf83e0b787f6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I82e534ecaabf5af6a9b6a567b862800a };
assign Idc7df6877bdb7e7d392307d78183d31c = (I58db79a8e9f0cd1ded379897ba2f27ae[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib184e1d3a451b69a5206cf83e0b787f6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00003_U (
.flogtanh_sel( I6d3cb4ccb4e51c7e6603d0abd1a082c4[flogtanh_SEL-1:0]),
.flogtanh( I1c9684b45467216a18a3a0d93b555b60),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If6d01c60d560e37c2676de16f9c10d20  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1c9684b45467216a18a3a0d93b555b60 };
assign Ib8b95ece5da3877b261a06e6d0571921 = (I6d3cb4ccb4e51c7e6603d0abd1a082c4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If6d01c60d560e37c2676de16f9c10d20;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00004_U (
.flogtanh_sel( I79f75f49ea8a29d684af396014b2f3ab[flogtanh_SEL-1:0]),
.flogtanh( Ice212c509101d6d41b52ea0cb85dacc0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic191abac086c847828546b8feea4fb23  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ice212c509101d6d41b52ea0cb85dacc0 };
assign Ic99654bf4833c9132912eeb4c0dc92fa = (I79f75f49ea8a29d684af396014b2f3ab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic191abac086c847828546b8feea4fb23;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00005_U (
.flogtanh_sel( I9c5ecd86bedb189fada40fae9d751a68[flogtanh_SEL-1:0]),
.flogtanh( I37ee7a2fab22cf8e6452fb408b849595),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I08c8ec03b53121517a27ff7fa143e5cb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I37ee7a2fab22cf8e6452fb408b849595 };
assign I2461055ef9b1aa2ffca0f5cac3300e71 = (I9c5ecd86bedb189fada40fae9d751a68[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I08c8ec03b53121517a27ff7fa143e5cb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00006_U (
.flogtanh_sel( Iad5f06e1989ead7d306c70a3b02cb8f4[flogtanh_SEL-1:0]),
.flogtanh( I0ec18ade132eede6849e0607af608726),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I52362ce3dd44269cdce0797f54886036  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0ec18ade132eede6849e0607af608726 };
assign I2bc3ffbe5b42b0833206437d3863278e = (Iad5f06e1989ead7d306c70a3b02cb8f4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I52362ce3dd44269cdce0797f54886036;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00007_U (
.flogtanh_sel( If6d1a410df5a4aea6a01337a6074fbd9[flogtanh_SEL-1:0]),
.flogtanh( I4651eab27cb766a1792f9564bcb2764a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib36da02cb5325af53c1cebe6e20b9468  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4651eab27cb766a1792f9564bcb2764a };
assign Id5e02d4c48fa6c3b0d45a9e66f09448f = (If6d1a410df5a4aea6a01337a6074fbd9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib36da02cb5325af53c1cebe6e20b9468;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00008_U (
.flogtanh_sel( I3bc40a4db14566b5099b14cee5f61135[flogtanh_SEL-1:0]),
.flogtanh( Ibbdbc4e4fc2ee018a0e7a4da29e85b56),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8be5606ad0efbff7ccb552566592ef15  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibbdbc4e4fc2ee018a0e7a4da29e85b56 };
assign I40e99289d5762e77a3766eb8251eef00 = (I3bc40a4db14566b5099b14cee5f61135[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8be5606ad0efbff7ccb552566592ef15;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00009_U (
.flogtanh_sel( I7e683fd8235d7cfbf4ff407a286f07de[flogtanh_SEL-1:0]),
.flogtanh( Ic67b9e090d6815b2a745bdc4983f9c69),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie70af982f7791be92f896afe027c8832  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic67b9e090d6815b2a745bdc4983f9c69 };
assign I20beb3fdbe91936f74a200cd8ec9817b = (I7e683fd8235d7cfbf4ff407a286f07de[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie70af982f7791be92f896afe027c8832;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00010_U (
.flogtanh_sel( I97afcedf05e588b7976d6005191dc916[flogtanh_SEL-1:0]),
.flogtanh( I8327267045af5da02c066a5eab25f13a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I93ed828faec287b2295a3f860d818fbe  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8327267045af5da02c066a5eab25f13a };
assign Id435b68afb53bef4afc7b70a9512e955 = (I97afcedf05e588b7976d6005191dc916[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I93ed828faec287b2295a3f860d818fbe;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00011_U (
.flogtanh_sel( Ib8d8eec0aaa662adf2837c9b705fce7e[flogtanh_SEL-1:0]),
.flogtanh( Id91ef7e27c689cdf5ce50d705017e40e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifea8cb28a2e829628ceae6126c81eb1f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id91ef7e27c689cdf5ce50d705017e40e };
assign I0cf5cb4cd472502b84dbf6fe1af0be78 = (Ib8d8eec0aaa662adf2837c9b705fce7e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifea8cb28a2e829628ceae6126c81eb1f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00028_00012_U (
.flogtanh_sel( Icbd765be950123705955e2c5d7ace84b[flogtanh_SEL-1:0]),
.flogtanh( I60498760f3c03cf92ceeb99c5096fe54),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idd12f95ce2cb0eb33dbbb09a235c3ca0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I60498760f3c03cf92ceeb99c5096fe54 };
assign Iacf6340a29a5592b61ea875304a2de48 = (Icbd765be950123705955e2c5d7ace84b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idd12f95ce2cb0eb33dbbb09a235c3ca0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00000_U (
.flogtanh_sel( I706e8f5617cfae1e6fc83db18c8b5fe3[flogtanh_SEL-1:0]),
.flogtanh( I63169dbc533400e0db5e37a8ebeca1aa),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2cfcf8d0beaa4aceb9182c835352b210  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I63169dbc533400e0db5e37a8ebeca1aa };
assign I5dfc71255cba279420b7545df4d35c40 = (I706e8f5617cfae1e6fc83db18c8b5fe3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2cfcf8d0beaa4aceb9182c835352b210;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00001_U (
.flogtanh_sel( I1dd8f8c7f1b673898096b1f3ae383197[flogtanh_SEL-1:0]),
.flogtanh( I150f11a565ad39c59d8f9e4c94d397e2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7bcc86543042aa717d956b83566442d2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I150f11a565ad39c59d8f9e4c94d397e2 };
assign Ibadcb205c7e9a0f3345cac7eb41b5985 = (I1dd8f8c7f1b673898096b1f3ae383197[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7bcc86543042aa717d956b83566442d2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00002_U (
.flogtanh_sel( I10ca8978cf4659265ed25a27d09acc1c[flogtanh_SEL-1:0]),
.flogtanh( Icadb816a238ba165425e5a30bd0bb8e6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4ae99bdc1aca92e0c7ebec69455db910  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icadb816a238ba165425e5a30bd0bb8e6 };
assign I762b2abb876381eff6de97cef0798405 = (I10ca8978cf4659265ed25a27d09acc1c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4ae99bdc1aca92e0c7ebec69455db910;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00003_U (
.flogtanh_sel( Iec4656b32460def4a608b6b0f6486af9[flogtanh_SEL-1:0]),
.flogtanh( I3b55785b9625ac53f6c00ba5a10a481b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I612ab97c8ff0b0000f5321336aa31481  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3b55785b9625ac53f6c00ba5a10a481b };
assign Ib3e7633767b6e09e4ee54f6feaddd31e = (Iec4656b32460def4a608b6b0f6486af9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I612ab97c8ff0b0000f5321336aa31481;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00004_U (
.flogtanh_sel( I5f4475897d1d58965da1b35fe0ef8c01[flogtanh_SEL-1:0]),
.flogtanh( If7317c81c9b6503386cab33fa812e80e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I837c986c9a0267bcb434c774c307542e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If7317c81c9b6503386cab33fa812e80e };
assign I3f193e9c265c1dfaeada63d59db5b79f = (I5f4475897d1d58965da1b35fe0ef8c01[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I837c986c9a0267bcb434c774c307542e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00005_U (
.flogtanh_sel( Ife61469306df3cf220666b187f1496a9[flogtanh_SEL-1:0]),
.flogtanh( I095672e79ca3a6dd8589b7821f06cdb9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7383d68c9e1c7c663a32233a8385435a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I095672e79ca3a6dd8589b7821f06cdb9 };
assign Ie72268e979cf069b88f6eadde789e5ab = (Ife61469306df3cf220666b187f1496a9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7383d68c9e1c7c663a32233a8385435a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00006_U (
.flogtanh_sel( Ib49319b9dfa4914f92f423ceaf840014[flogtanh_SEL-1:0]),
.flogtanh( Ibf2f43980e835dd7ae7535957e3ec131),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8726f6e59d2146674ad4fae01d7f4135  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibf2f43980e835dd7ae7535957e3ec131 };
assign I5732fdb805258fc13c8ba4aaf56574ca = (Ib49319b9dfa4914f92f423ceaf840014[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8726f6e59d2146674ad4fae01d7f4135;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00007_U (
.flogtanh_sel( I93ff2f879233cac9b9f0dd2f4c082c09[flogtanh_SEL-1:0]),
.flogtanh( Iaa980a50205025e3e1b09c6ce8ee53dd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3a754b15a3a7d47b3a9741f4982a0a32  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iaa980a50205025e3e1b09c6ce8ee53dd };
assign I3afe987d8f2c93cc19534a3221d1939c = (I93ff2f879233cac9b9f0dd2f4c082c09[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3a754b15a3a7d47b3a9741f4982a0a32;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00008_U (
.flogtanh_sel( I44597d694e9c5d29280e503d72a27c8d[flogtanh_SEL-1:0]),
.flogtanh( I829aa657f0dd13c3fb86baeda8a3b4c8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9bd8a06d5fdfe50c340c649a678ba2e2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I829aa657f0dd13c3fb86baeda8a3b4c8 };
assign Ic66af6c3c0268cfb0e9f0776c4f4e961 = (I44597d694e9c5d29280e503d72a27c8d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9bd8a06d5fdfe50c340c649a678ba2e2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00009_U (
.flogtanh_sel( I04a19448c5e75af8021ad02d1a708bb0[flogtanh_SEL-1:0]),
.flogtanh( I1ae4334c32094064c19df0dac77bd03d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I215cb4bca0e3579af6474dbd9462304c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1ae4334c32094064c19df0dac77bd03d };
assign Ia605d14205926b3edc6d1c2f69f70ac0 = (I04a19448c5e75af8021ad02d1a708bb0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I215cb4bca0e3579af6474dbd9462304c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00010_U (
.flogtanh_sel( I71a3093121c2f19dcd1412b468652fa8[flogtanh_SEL-1:0]),
.flogtanh( I78788f7e0845e4353145012efa04a48c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6d73cf92b5ad3ded496cf1363c87d3ad  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I78788f7e0845e4353145012efa04a48c };
assign I0071f2168787bd42ab7f2370aed9d0f5 = (I71a3093121c2f19dcd1412b468652fa8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6d73cf92b5ad3ded496cf1363c87d3ad;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00011_U (
.flogtanh_sel( I3ae09c82029c617034fe6aacbe9e94e6[flogtanh_SEL-1:0]),
.flogtanh( I359f3e3bb2a69349f8564466fa81a054),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I47851422267c2963b3c93e029e81fe1e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I359f3e3bb2a69349f8564466fa81a054 };
assign I4936f823841b0ffe32f801f5134c0211 = (I3ae09c82029c617034fe6aacbe9e94e6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I47851422267c2963b3c93e029e81fe1e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00029_00012_U (
.flogtanh_sel( Ie7af6b3b441f910b000a333afad6c76f[flogtanh_SEL-1:0]),
.flogtanh( I7b630e8ac26638fb858dd3b5d2d56385),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie9cd13f4f83e446d41fa362d0ca005c2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7b630e8ac26638fb858dd3b5d2d56385 };
assign I5975ef8f6cf53cf2132cdd9d707e7912 = (Ie7af6b3b441f910b000a333afad6c76f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie9cd13f4f83e446d41fa362d0ca005c2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00000_U (
.flogtanh_sel( I4d71dfea8407aa5b5cbb991bc4fea963[flogtanh_SEL-1:0]),
.flogtanh( I859bef71501c2f2a994a0cdf8a94b2a7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9990a45631a11aa0b051d237de4cb71f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I859bef71501c2f2a994a0cdf8a94b2a7 };
assign I954ff0f9ee871a31774a3d786128fa13 = (I4d71dfea8407aa5b5cbb991bc4fea963[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9990a45631a11aa0b051d237de4cb71f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00001_U (
.flogtanh_sel( I1a082caecc831a90e74674ba35da4183[flogtanh_SEL-1:0]),
.flogtanh( Ib51b9e41161f4273f6469e8965acd7dd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4be57c0a1c49baa53daba558c939eee0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib51b9e41161f4273f6469e8965acd7dd };
assign I31f6bbfbbbd4c20d0c5c71663da1d4c1 = (I1a082caecc831a90e74674ba35da4183[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4be57c0a1c49baa53daba558c939eee0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00002_U (
.flogtanh_sel( Iec1de44616a2354a56ab1f681059d4c5[flogtanh_SEL-1:0]),
.flogtanh( I78bb23c008613c0f07f6f85172482296),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I16d8c346fd377bc293763e9cb683566e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I78bb23c008613c0f07f6f85172482296 };
assign I1898bc3cc6a8b6f71d65c758d1f08366 = (Iec1de44616a2354a56ab1f681059d4c5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I16d8c346fd377bc293763e9cb683566e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00003_U (
.flogtanh_sel( Ie3c2318e64d0e218c3db557404c4aac8[flogtanh_SEL-1:0]),
.flogtanh( I8b883a5bc22b2cde03f4074357be7c88),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9df0b548fc5a23180b48207dc7fc603e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8b883a5bc22b2cde03f4074357be7c88 };
assign If86532f849bd392dbf599eeb2fae0545 = (Ie3c2318e64d0e218c3db557404c4aac8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9df0b548fc5a23180b48207dc7fc603e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00004_U (
.flogtanh_sel( I9a251d50f41e51b1a5cc2475f267e8a0[flogtanh_SEL-1:0]),
.flogtanh( Ic2727e097ffbce70f07fc9f3d9395b54),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0b3b2dd5a443fab695d0ff59634b6cb6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic2727e097ffbce70f07fc9f3d9395b54 };
assign Ia344734d285ac29b53cf401c08a0f987 = (I9a251d50f41e51b1a5cc2475f267e8a0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0b3b2dd5a443fab695d0ff59634b6cb6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00005_U (
.flogtanh_sel( I9b5767a49f7b9dcb8fdaea924835033c[flogtanh_SEL-1:0]),
.flogtanh( I096397439036b0056c979054528ce1fd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6f66b0df384980fcbf6a92e5a197575e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I096397439036b0056c979054528ce1fd };
assign I502a8e382aa0881dc86f3c13e0566ca3 = (I9b5767a49f7b9dcb8fdaea924835033c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6f66b0df384980fcbf6a92e5a197575e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00006_U (
.flogtanh_sel( I6ca1e6700a19d03621a193c7240bff54[flogtanh_SEL-1:0]),
.flogtanh( Ifcc83d9007aafdf32acf04f062e008c8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2aff93633ddb7f63312e991dab99cfca  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifcc83d9007aafdf32acf04f062e008c8 };
assign Ic462cebbfc39190b22d20013259e39eb = (I6ca1e6700a19d03621a193c7240bff54[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2aff93633ddb7f63312e991dab99cfca;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00007_U (
.flogtanh_sel( I931c597ff12bffce581f653346202f83[flogtanh_SEL-1:0]),
.flogtanh( I53c01c60f4061d970e4491564ddf88ae),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic17e0c2adccfc8b88818591fb7c3958a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I53c01c60f4061d970e4491564ddf88ae };
assign I385d03def4cfb49f54867687ebd710ed = (I931c597ff12bffce581f653346202f83[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic17e0c2adccfc8b88818591fb7c3958a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00008_U (
.flogtanh_sel( Ia3a2c5d59f6340917ca3933c05ba4678[flogtanh_SEL-1:0]),
.flogtanh( I0b4d34aa164c014f9315debd37fa534b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I835b69f77b77fcb0bb1cc9a05a9964c4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0b4d34aa164c014f9315debd37fa534b };
assign If8aa3ec1b5a4a3c122da82467be917da = (Ia3a2c5d59f6340917ca3933c05ba4678[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I835b69f77b77fcb0bb1cc9a05a9964c4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00009_U (
.flogtanh_sel( Ie83d0a8ee5ed214bc7577467748aaa04[flogtanh_SEL-1:0]),
.flogtanh( Iac97aad4ca2c93e387ff0c1340143029),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iac61d3d6b4ebec5460d07a209317dbf6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iac97aad4ca2c93e387ff0c1340143029 };
assign I8daf79a0a2ee1bac7f055af441539fa4 = (Ie83d0a8ee5ed214bc7577467748aaa04[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iac61d3d6b4ebec5460d07a209317dbf6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00010_U (
.flogtanh_sel( Iaac29552e5fc65aaf4f0116f917b707c[flogtanh_SEL-1:0]),
.flogtanh( I8b4c2d8a5f2b796029575ecf3b89e2b9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I762215c24e6cfbb27328534b48f6c013  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8b4c2d8a5f2b796029575ecf3b89e2b9 };
assign I6261e0d339762cb2364421e6b87086cb = (Iaac29552e5fc65aaf4f0116f917b707c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I762215c24e6cfbb27328534b48f6c013;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00011_U (
.flogtanh_sel( Ie2c8eac7204b98139c03b6fbfff9af36[flogtanh_SEL-1:0]),
.flogtanh( I06dd747316fa36a8dbdbb4ddf011230b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I278647e72fba32b7725004a889c40fb0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I06dd747316fa36a8dbdbb4ddf011230b };
assign I0e2f746715b901feb69f6b3c94f3a828 = (Ie2c8eac7204b98139c03b6fbfff9af36[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I278647e72fba32b7725004a889c40fb0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00030_00012_U (
.flogtanh_sel( Ied7fcdaec662cb3c2f89f131986fa102[flogtanh_SEL-1:0]),
.flogtanh( I1594e7dfaedd9e7f5818dc4d639bb663),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib6b14ee93e905e08b910d6011d780bf9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1594e7dfaedd9e7f5818dc4d639bb663 };
assign I7b8da162c08f8aa2ae90522ee1526cf6 = (Ied7fcdaec662cb3c2f89f131986fa102[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib6b14ee93e905e08b910d6011d780bf9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00000_U (
.flogtanh_sel( Ib16a17d6430570b45a304d847ee2b11c[flogtanh_SEL-1:0]),
.flogtanh( Ic8111eb95e6b6ab35bcd8e2cafcd0c1e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6f89d12b0e9b153b01cd8fd0e548a5ab  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic8111eb95e6b6ab35bcd8e2cafcd0c1e };
assign I5e8ecdbb018402b2fbc0049ee44bae8c = (Ib16a17d6430570b45a304d847ee2b11c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6f89d12b0e9b153b01cd8fd0e548a5ab;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00001_U (
.flogtanh_sel( I42169e454756fe4d1c5f17f2eeb2e091[flogtanh_SEL-1:0]),
.flogtanh( I650b4641d233096a77ae15c8254a29b1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I63ba8ed824c286ff8f68ffb6cb10a12c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I650b4641d233096a77ae15c8254a29b1 };
assign I06d859184884c07a14c83d2f06587ad5 = (I42169e454756fe4d1c5f17f2eeb2e091[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I63ba8ed824c286ff8f68ffb6cb10a12c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00002_U (
.flogtanh_sel( I6fde38a3a92e06fa77123e3279813c41[flogtanh_SEL-1:0]),
.flogtanh( Ia905d37c471bdf7258a547be95b85e4f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib54c1747fb4316314527140212c7cc60  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia905d37c471bdf7258a547be95b85e4f };
assign I79e3e49f57d47231c0fe6aaafdbc57f1 = (I6fde38a3a92e06fa77123e3279813c41[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib54c1747fb4316314527140212c7cc60;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00003_U (
.flogtanh_sel( Id8ee16437e8d6d6da6d37440e04097b6[flogtanh_SEL-1:0]),
.flogtanh( Icfc2b5de1aa36d81de3f163880d48a68),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idfaaf824ddb5452930ca1997f057e321  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icfc2b5de1aa36d81de3f163880d48a68 };
assign I12c07042202f66db926861c9ce7c2b25 = (Id8ee16437e8d6d6da6d37440e04097b6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idfaaf824ddb5452930ca1997f057e321;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00004_U (
.flogtanh_sel( Ibf249d8e5acced9b064132575f40e001[flogtanh_SEL-1:0]),
.flogtanh( I3c6893d360627cd954db1c20f3c9d319),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I372410e0c71fce0d0a592bf9f16f822d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3c6893d360627cd954db1c20f3c9d319 };
assign I9d0fdb45b9e86bd409740e538a690320 = (Ibf249d8e5acced9b064132575f40e001[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I372410e0c71fce0d0a592bf9f16f822d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00005_U (
.flogtanh_sel( I580659084e3d17b48de6b1c66154fcf5[flogtanh_SEL-1:0]),
.flogtanh( Ibc971e0b7ade69365d2c23f30ba0c1ea),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie9392382734808bcff4da7e0c7f8e4d3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibc971e0b7ade69365d2c23f30ba0c1ea };
assign Id5fd6f25dc3df22a322434ae3c90dea6 = (I580659084e3d17b48de6b1c66154fcf5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie9392382734808bcff4da7e0c7f8e4d3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00006_U (
.flogtanh_sel( I7a14e45d43ab77b265501902152c8616[flogtanh_SEL-1:0]),
.flogtanh( I562d9a1676d27c7966d2920bb6be3b38),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If703357df55e47b3ab1fbb1126ad5160  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I562d9a1676d27c7966d2920bb6be3b38 };
assign Id812a8ea2a3b4a912d151be582833fcf = (I7a14e45d43ab77b265501902152c8616[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If703357df55e47b3ab1fbb1126ad5160;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00007_U (
.flogtanh_sel( I81ba868784103e0eb05a44d981d4d666[flogtanh_SEL-1:0]),
.flogtanh( I8aa258f382bea1eb300b006c3083bec1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I69e05d54d008abdfb8d0b2d1ddc0fd49  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8aa258f382bea1eb300b006c3083bec1 };
assign Ifd3638d44e1ba2285891fac152dee327 = (I81ba868784103e0eb05a44d981d4d666[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I69e05d54d008abdfb8d0b2d1ddc0fd49;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00008_U (
.flogtanh_sel( Ic6b88783957cbaf253648a30b22f6b1c[flogtanh_SEL-1:0]),
.flogtanh( Iec0e7232ec94c15d7d50866ad5eb85fb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic79dc94346350619e49087d1d399bc39  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iec0e7232ec94c15d7d50866ad5eb85fb };
assign Idd1b6014de2f053554ed09c29bf3e640 = (Ic6b88783957cbaf253648a30b22f6b1c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic79dc94346350619e49087d1d399bc39;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00009_U (
.flogtanh_sel( I4103c218a85a1d08db5c4f4b5686b2e5[flogtanh_SEL-1:0]),
.flogtanh( I0d252b23e06d25aee4afd84b4c5b4ba9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib805b36c4865846137bb8c620ee711bb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0d252b23e06d25aee4afd84b4c5b4ba9 };
assign I0d96336eb4d5071d7e1d350e86513b25 = (I4103c218a85a1d08db5c4f4b5686b2e5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib805b36c4865846137bb8c620ee711bb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00010_U (
.flogtanh_sel( I0e6c0958af503e4a120a49d02a432863[flogtanh_SEL-1:0]),
.flogtanh( I430703cef7ec173f9099c8391132e5c4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8af4ba916324c47b2773e25e81eec395  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I430703cef7ec173f9099c8391132e5c4 };
assign I31e5b2cdc3dc571eafa37510076bcc64 = (I0e6c0958af503e4a120a49d02a432863[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8af4ba916324c47b2773e25e81eec395;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00011_U (
.flogtanh_sel( I8f76b31e8f15c0e5fe24dcb723418111[flogtanh_SEL-1:0]),
.flogtanh( I5788d966ba8393f5d76dcfcb9294b52e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I43bf51dd2065c4699e2efb0d23ca67fc  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5788d966ba8393f5d76dcfcb9294b52e };
assign Ia8849f78971a45ed0daa2489e7d27dd7 = (I8f76b31e8f15c0e5fe24dcb723418111[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I43bf51dd2065c4699e2efb0d23ca67fc;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00031_00012_U (
.flogtanh_sel( Id1457221b58344b60070aa026436df2c[flogtanh_SEL-1:0]),
.flogtanh( Ied561890134d28b451f26da773ea5525),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie42fb8850ec075e738c9265ef746d0a2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ied561890134d28b451f26da773ea5525 };
assign Ie4749f8e9ad2b370f9f9814b5a463c43 = (Id1457221b58344b60070aa026436df2c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie42fb8850ec075e738c9265ef746d0a2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00032_00000_U (
.flogtanh_sel( Icc31966508e03d8869e81d8aeb243705[flogtanh_SEL-1:0]),
.flogtanh( I52e018ad790a1e406777510a0f4b6c29),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I734fecd29be258bbcf174ce05a4ad7c7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I52e018ad790a1e406777510a0f4b6c29 };
assign I3096d11098113da669ee0a94686e600d = (Icc31966508e03d8869e81d8aeb243705[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I734fecd29be258bbcf174ce05a4ad7c7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00032_00001_U (
.flogtanh_sel( I9dcccf542ba434b6e0fde6f012f98f92[flogtanh_SEL-1:0]),
.flogtanh( I25eb66d8589cbb35b32cd25539a24f7f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I90c0a469b49cec5817be9ee089d7f035  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I25eb66d8589cbb35b32cd25539a24f7f };
assign I09a1d04c307fcb8a0e30925d86df3fe9 = (I9dcccf542ba434b6e0fde6f012f98f92[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I90c0a469b49cec5817be9ee089d7f035;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00032_00002_U (
.flogtanh_sel( I51ccbb824a5e1e340eefd173c4491728[flogtanh_SEL-1:0]),
.flogtanh( Icd4716d0d66d95a532544461c4872d11),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I20467038010337e3e125bf2a7e1302d4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icd4716d0d66d95a532544461c4872d11 };
assign Idb0a98cea3ee6cd4308bfc2414a003e1 = (I51ccbb824a5e1e340eefd173c4491728[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I20467038010337e3e125bf2a7e1302d4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00032_00003_U (
.flogtanh_sel( Ib7ae1730dcd8bc708bbfcc6a9f97ac66[flogtanh_SEL-1:0]),
.flogtanh( I266ba4229056534d310d982253b5f9b9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idc01d14ecbd22e73d7ee052989eacff6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I266ba4229056534d310d982253b5f9b9 };
assign Id4788855f9a503e8b506d012aaeea445 = (Ib7ae1730dcd8bc708bbfcc6a9f97ac66[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idc01d14ecbd22e73d7ee052989eacff6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00032_00004_U (
.flogtanh_sel( I4714f5c91203fcfa552f0fcf71b87442[flogtanh_SEL-1:0]),
.flogtanh( I86498c8c820d276ac12764b5df267252),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If3410ef0f48854e7b788d74904d03dad  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I86498c8c820d276ac12764b5df267252 };
assign I5b937934e7aae1f916c2848889f12685 = (I4714f5c91203fcfa552f0fcf71b87442[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If3410ef0f48854e7b788d74904d03dad;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00032_00005_U (
.flogtanh_sel( I3b6d1e84fdd1019249886fa5fe65895b[flogtanh_SEL-1:0]),
.flogtanh( I7bb9ad1a2cd32966746b05b7604a09b6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icba9bcbb58a3fef701c5572510dbba65  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7bb9ad1a2cd32966746b05b7604a09b6 };
assign I9275bb36e58e0f17964e13ee7f027ab7 = (I3b6d1e84fdd1019249886fa5fe65895b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icba9bcbb58a3fef701c5572510dbba65;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00033_00000_U (
.flogtanh_sel( Ia8a7d4207dbabc7970bf36f3fe74f72d[flogtanh_SEL-1:0]),
.flogtanh( Id0998cc2848a6a72ed2701a8e720946e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ice5cb3b187d142f36c9fe4673952b229  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id0998cc2848a6a72ed2701a8e720946e };
assign I02330ade2eed926076cc071e45eed82c = (Ia8a7d4207dbabc7970bf36f3fe74f72d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ice5cb3b187d142f36c9fe4673952b229;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00033_00001_U (
.flogtanh_sel( I84047457b43ef33874f4550c3b773460[flogtanh_SEL-1:0]),
.flogtanh( If1ed051cd94d42e7836f82c10538b302),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id382353b13f6d198e0e9b90c5c3c16b3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If1ed051cd94d42e7836f82c10538b302 };
assign I296bc392d4223cbdd6f77be6523df819 = (I84047457b43ef33874f4550c3b773460[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id382353b13f6d198e0e9b90c5c3c16b3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00033_00002_U (
.flogtanh_sel( I5e51563c3e69beca0b463742e6e5f9ee[flogtanh_SEL-1:0]),
.flogtanh( I780afd116929565d1ff9b3833ba242d5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I83efee0bf505cf1258bb68e419ffccf7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I780afd116929565d1ff9b3833ba242d5 };
assign I31b0f2fe98cfddbc05dbd14be8be394b = (I5e51563c3e69beca0b463742e6e5f9ee[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I83efee0bf505cf1258bb68e419ffccf7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00033_00003_U (
.flogtanh_sel( I6c8d14e31c80811ccab1b6ab09d28089[flogtanh_SEL-1:0]),
.flogtanh( I89ee99e699676bcec20031b6cad0e2ac),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id54f91bbae7215f942f539ca0834bd1f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I89ee99e699676bcec20031b6cad0e2ac };
assign Ia71663e8f563041c27cd21a0c9c27a28 = (I6c8d14e31c80811ccab1b6ab09d28089[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id54f91bbae7215f942f539ca0834bd1f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00033_00004_U (
.flogtanh_sel( I50b3b7490c9b65b6e662cc86b163a2df[flogtanh_SEL-1:0]),
.flogtanh( I862b467403c045e4694fb57d59e10064),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I810c80a4b57d13add447ee8964844ce1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I862b467403c045e4694fb57d59e10064 };
assign Ib46b13498ec14ceaa56719f26f18febb = (I50b3b7490c9b65b6e662cc86b163a2df[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I810c80a4b57d13add447ee8964844ce1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00033_00005_U (
.flogtanh_sel( I8351a2110a3d73ad8803cf17e3317017[flogtanh_SEL-1:0]),
.flogtanh( Ic3b554c66f652f027159dbc0fccc5ba3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icf6d317a1bca3a6f3dfafdc9bdc0b805  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic3b554c66f652f027159dbc0fccc5ba3 };
assign I9bc2d5692474b8368c570d92835191b3 = (I8351a2110a3d73ad8803cf17e3317017[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icf6d317a1bca3a6f3dfafdc9bdc0b805;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00034_00000_U (
.flogtanh_sel( I1e6c696951688d581f21ab2302593335[flogtanh_SEL-1:0]),
.flogtanh( I04635713f6d70142b7ab3ecb5ffe6ac9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I47ca60b0a9bec684ec4e52f28f76c6d7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I04635713f6d70142b7ab3ecb5ffe6ac9 };
assign If8b0b96a659183e3651c691a2848b86b = (I1e6c696951688d581f21ab2302593335[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I47ca60b0a9bec684ec4e52f28f76c6d7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00034_00001_U (
.flogtanh_sel( Ie9840e28133eebdca0be313552195c7b[flogtanh_SEL-1:0]),
.flogtanh( I1917eae0dbcc0a941718c3248c7d4b11),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6ae68bcd4f3d39661626e4b671acf4ea  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1917eae0dbcc0a941718c3248c7d4b11 };
assign I87d958c00fc6209d901147831b0c951c = (Ie9840e28133eebdca0be313552195c7b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6ae68bcd4f3d39661626e4b671acf4ea;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00034_00002_U (
.flogtanh_sel( I82812258a8032e273cab7139266be1b6[flogtanh_SEL-1:0]),
.flogtanh( Ifa60c3079164485f31442d9cf12bd2ad),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaa25b6dc9ec478e1fe096bfb9013752c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifa60c3079164485f31442d9cf12bd2ad };
assign Ie4e4eaf3e5d2f581210af8054df71c6c = (I82812258a8032e273cab7139266be1b6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaa25b6dc9ec478e1fe096bfb9013752c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00034_00003_U (
.flogtanh_sel( I27ab6fd9927518e29ed36d7a7a241498[flogtanh_SEL-1:0]),
.flogtanh( I5616405acf49c3e8608ae4d2b544b0d6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If7f010576686a2eb7aa5b2307c02ad6b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5616405acf49c3e8608ae4d2b544b0d6 };
assign I0b557cf102da41afd26936cbdb64b6e8 = (I27ab6fd9927518e29ed36d7a7a241498[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If7f010576686a2eb7aa5b2307c02ad6b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00034_00004_U (
.flogtanh_sel( I05b0f33a3808ac53b29d8d8309447650[flogtanh_SEL-1:0]),
.flogtanh( Ie6f9ae463fa1add4de23463435a23d25),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie8a683efbffce7c5676fa831573299d7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie6f9ae463fa1add4de23463435a23d25 };
assign I49eb064043f91112c854e31e4eb9b885 = (I05b0f33a3808ac53b29d8d8309447650[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie8a683efbffce7c5676fa831573299d7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00034_00005_U (
.flogtanh_sel( If150ebf242231f0d22c996a71552f6eb[flogtanh_SEL-1:0]),
.flogtanh( Ib16a67d67a4650e53547312e3af60363),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I50a4545b75d92b3c3209d473f8d0647c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib16a67d67a4650e53547312e3af60363 };
assign I1039bc43e88eee527d2ed6adb8c7d1ba = (If150ebf242231f0d22c996a71552f6eb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I50a4545b75d92b3c3209d473f8d0647c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00035_00000_U (
.flogtanh_sel( If2d0a2b58510715e74787cb60719cb5b[flogtanh_SEL-1:0]),
.flogtanh( I8fa4ad645ca2ef21dea8669d2e2afbe2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib0e11d415f14d70a626c6f0dfeed2e37  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8fa4ad645ca2ef21dea8669d2e2afbe2 };
assign I9aab16e89f1b64117caece8ca8af5940 = (If2d0a2b58510715e74787cb60719cb5b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib0e11d415f14d70a626c6f0dfeed2e37;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00035_00001_U (
.flogtanh_sel( Ib6745a6d17034a29501e022bd846bf2f[flogtanh_SEL-1:0]),
.flogtanh( I41ea2e3d798ff8e0a95f04e4773c59b4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3a6167a349b5dce1dfa66859bfd5eee7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I41ea2e3d798ff8e0a95f04e4773c59b4 };
assign I343df614f97cf732e57cf2ad3f95dc9e = (Ib6745a6d17034a29501e022bd846bf2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3a6167a349b5dce1dfa66859bfd5eee7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00035_00002_U (
.flogtanh_sel( Iae09c127dfe86c9f7bdbeff447c777f5[flogtanh_SEL-1:0]),
.flogtanh( Id7f4c6208197cdbf48fecdb2a18b81fc),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I566fd98c8c6ebf6e2d8ebace4b8b358b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id7f4c6208197cdbf48fecdb2a18b81fc };
assign Ie02de90d8eb06b16314946d21299500c = (Iae09c127dfe86c9f7bdbeff447c777f5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I566fd98c8c6ebf6e2d8ebace4b8b358b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00035_00003_U (
.flogtanh_sel( I742128de6b237ed48e3a7ccd3788f0d7[flogtanh_SEL-1:0]),
.flogtanh( I0adb66417482782dd71da1678c1f7412),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib777f0ff44b2847294370d74f741b70b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0adb66417482782dd71da1678c1f7412 };
assign I3353a7916b569f2c0ca122180608dccc = (I742128de6b237ed48e3a7ccd3788f0d7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib777f0ff44b2847294370d74f741b70b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00035_00004_U (
.flogtanh_sel( Id5e8fda13ba8f6d95d694d0f30da75bb[flogtanh_SEL-1:0]),
.flogtanh( I2abe89a1366a1ad862266ad88101baa2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6cd7374654c74b4be21b6a3639ddac0f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2abe89a1366a1ad862266ad88101baa2 };
assign Ibfe760474fcac99f1e5ffa2e008fef99 = (Id5e8fda13ba8f6d95d694d0f30da75bb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6cd7374654c74b4be21b6a3639ddac0f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00035_00005_U (
.flogtanh_sel( I1aa5a04e40f9b1685c77e4d101c3ccf4[flogtanh_SEL-1:0]),
.flogtanh( I8d10f0c6dc026005f7882ca013283099),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I930319dcb4988822341ac101fef3dc52  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8d10f0c6dc026005f7882ca013283099 };
assign I3caf1211dcbcdc746a3e4c7fbbdae4a8 = (I1aa5a04e40f9b1685c77e4d101c3ccf4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I930319dcb4988822341ac101fef3dc52;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00036_00000_U (
.flogtanh_sel( Ife1adea26d13bc299bb2de241ad4a6ea[flogtanh_SEL-1:0]),
.flogtanh( I4ef16908ce9b89771f94068eec1a983e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If556f828f8cb4c1f1721e9d12977ec5a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4ef16908ce9b89771f94068eec1a983e };
assign I2dcc0d17b9fcac35693bf32b5c5540fd = (Ife1adea26d13bc299bb2de241ad4a6ea[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If556f828f8cb4c1f1721e9d12977ec5a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00036_00001_U (
.flogtanh_sel( Ifcf6c761f0f253921710af87ab1d2247[flogtanh_SEL-1:0]),
.flogtanh( I4f6bcd6e0bcd77730248b69d2b93c904),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If7df1cceb63540263742300063a2febb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4f6bcd6e0bcd77730248b69d2b93c904 };
assign Ie6764a631310e312ba5c2c1e601d828f = (Ifcf6c761f0f253921710af87ab1d2247[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If7df1cceb63540263742300063a2febb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00036_00002_U (
.flogtanh_sel( I1478e6a9113c124bdc4361908af6643f[flogtanh_SEL-1:0]),
.flogtanh( Iea1ae39e18f083fb8f855fd9ad3d4f8e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idb605ffe97f2a0cbc2b260464afd1479  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iea1ae39e18f083fb8f855fd9ad3d4f8e };
assign I220f8e45e5fe6e69f02cded87f12e1e5 = (I1478e6a9113c124bdc4361908af6643f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idb605ffe97f2a0cbc2b260464afd1479;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00036_00003_U (
.flogtanh_sel( I0afd42151925883835844cf5deef6156[flogtanh_SEL-1:0]),
.flogtanh( I795ae30dec63ef2952917eb3355148a2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8690851e49869591791e5202e2ef2432  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I795ae30dec63ef2952917eb3355148a2 };
assign I896cd566a3d078b0f697a788efd223f2 = (I0afd42151925883835844cf5deef6156[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8690851e49869591791e5202e2ef2432;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00036_00004_U (
.flogtanh_sel( I2b4ab0aadffb3a1bb86f45ebc8acf085[flogtanh_SEL-1:0]),
.flogtanh( I188813c5474bf304b59dbe07c78bef6f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I60d3d03ea9219db9501568fb71d87df0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I188813c5474bf304b59dbe07c78bef6f };
assign I7caa41076a293edf18c7c4309fdcfc91 = (I2b4ab0aadffb3a1bb86f45ebc8acf085[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I60d3d03ea9219db9501568fb71d87df0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00036_00005_U (
.flogtanh_sel( Iffa867719ba9c31a8756cc5e6bf81147[flogtanh_SEL-1:0]),
.flogtanh( I1760a42d85513ea751e94a8b829b5f1a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib7f80c4193c311c6c553f15f0d9e0e09  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1760a42d85513ea751e94a8b829b5f1a };
assign I928a0e4951208aab170656596f456209 = (Iffa867719ba9c31a8756cc5e6bf81147[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib7f80c4193c311c6c553f15f0d9e0e09;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00036_00006_U (
.flogtanh_sel( Ibb62b6cb003f0d5549c864075f23d19b[flogtanh_SEL-1:0]),
.flogtanh( I8c652055cfcd230426887e171eaf2511),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3dfabb54fefcb9b9896e52446a1edc25  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8c652055cfcd230426887e171eaf2511 };
assign Ia3d129fd297905bee180293c0c39d9ef = (Ibb62b6cb003f0d5549c864075f23d19b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3dfabb54fefcb9b9896e52446a1edc25;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00036_00007_U (
.flogtanh_sel( I3690d101ae99f258cc58b4482cc378c8[flogtanh_SEL-1:0]),
.flogtanh( I9a88a91b0fcc6dd1a7b4ed24e676d9e1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If35ab032940f067a7905284b5f34a795  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9a88a91b0fcc6dd1a7b4ed24e676d9e1 };
assign Id555c88cf7f0904db74d45cc75c8f5d6 = (I3690d101ae99f258cc58b4482cc378c8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If35ab032940f067a7905284b5f34a795;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00037_00000_U (
.flogtanh_sel( Id597e95ce8a168ab67890085a26870d0[flogtanh_SEL-1:0]),
.flogtanh( I89f6566e2295d58668e63b9529d94df8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I11cbc38d0e7e8bb159707d0b6a312049  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I89f6566e2295d58668e63b9529d94df8 };
assign I1ddfd31bbf062aa5c3c71d61e492e3a2 = (Id597e95ce8a168ab67890085a26870d0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I11cbc38d0e7e8bb159707d0b6a312049;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00037_00001_U (
.flogtanh_sel( I98df60eb8f65641f9cccce4023be905c[flogtanh_SEL-1:0]),
.flogtanh( I08295c218fd06a8900974edc9c2924f2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib39a30cd08168accc0c3ca3bda467878  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I08295c218fd06a8900974edc9c2924f2 };
assign Iae9e023628eb6686708b2656f15616cc = (I98df60eb8f65641f9cccce4023be905c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib39a30cd08168accc0c3ca3bda467878;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00037_00002_U (
.flogtanh_sel( Ibcb4fbdee372353b79c460cdeafdfe4e[flogtanh_SEL-1:0]),
.flogtanh( I0a39fdea8b5bfac1862f199152e26ffe),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I44afd98669c6e6bf5054d677de2b919c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0a39fdea8b5bfac1862f199152e26ffe };
assign If4b100d26126e460c41b8c1bc8fbbb96 = (Ibcb4fbdee372353b79c460cdeafdfe4e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I44afd98669c6e6bf5054d677de2b919c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00037_00003_U (
.flogtanh_sel( I74dbf75966d047a4a9e91c1bc793666f[flogtanh_SEL-1:0]),
.flogtanh( Ib36a71ff310882325be0a2745e48f708),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic75ef170613d6b56ad3928b88f1abef5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib36a71ff310882325be0a2745e48f708 };
assign I85a7fede715578be0634d71e9c7951cd = (I74dbf75966d047a4a9e91c1bc793666f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic75ef170613d6b56ad3928b88f1abef5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00037_00004_U (
.flogtanh_sel( I79b8d9f9447c4c1b551ec6c1e8903040[flogtanh_SEL-1:0]),
.flogtanh( I75e4d037cc2ed0b0f75fc1fe9cb21da3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If541dad0db59ce6598cc87b2ecf6d76a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I75e4d037cc2ed0b0f75fc1fe9cb21da3 };
assign I2d7715a3af03d9664729fa6df85034a2 = (I79b8d9f9447c4c1b551ec6c1e8903040[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If541dad0db59ce6598cc87b2ecf6d76a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00037_00005_U (
.flogtanh_sel( Ib34b66548621fabe0753223712b1369f[flogtanh_SEL-1:0]),
.flogtanh( Iee9e9849924642a9579a10655624fa17),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3e9f3d8ae099408fe2ff46ae3aff430e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iee9e9849924642a9579a10655624fa17 };
assign I571ddcb0a10938e4c0816c965214b4a8 = (Ib34b66548621fabe0753223712b1369f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3e9f3d8ae099408fe2ff46ae3aff430e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00037_00006_U (
.flogtanh_sel( Ie5b3eb4c00bedfaecc3215d43ff28362[flogtanh_SEL-1:0]),
.flogtanh( I0a267feb8313c9fa5c663a3fe68284dd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6688f7cccc769490e870707ba9c14991  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0a267feb8313c9fa5c663a3fe68284dd };
assign I8bf8b0cf27a2654a0e7fdf3255945b67 = (Ie5b3eb4c00bedfaecc3215d43ff28362[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6688f7cccc769490e870707ba9c14991;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00037_00007_U (
.flogtanh_sel( Icf3a1b0b6dbcf959b44379024f3c4169[flogtanh_SEL-1:0]),
.flogtanh( I0e0ff3511e65a1dda10ec944c89d09d7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I89d5eb773f6c952c1ed5e5c57fed6fe1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0e0ff3511e65a1dda10ec944c89d09d7 };
assign I63f82f075d53205b5b556c0054f1a0b8 = (Icf3a1b0b6dbcf959b44379024f3c4169[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I89d5eb773f6c952c1ed5e5c57fed6fe1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00038_00000_U (
.flogtanh_sel( I918c2bbe7c71f8c6a07b0bad8811f4e7[flogtanh_SEL-1:0]),
.flogtanh( I4504a0a17633d26163a0afae21ad0f43),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia55fb2a1a8fcd959e3dd99403cd39a97  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4504a0a17633d26163a0afae21ad0f43 };
assign I3c6fb0df5846a19228a4e6cf9f9106ac = (I918c2bbe7c71f8c6a07b0bad8811f4e7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia55fb2a1a8fcd959e3dd99403cd39a97;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00038_00001_U (
.flogtanh_sel( Iedd960a21b1c08b4a5293cff200218b3[flogtanh_SEL-1:0]),
.flogtanh( Ibd7b7f4ba86b6c61a0dd38f71c67ae05),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I51a2b9abfab582408aeea3130d1e8334  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibd7b7f4ba86b6c61a0dd38f71c67ae05 };
assign I7168b0efdd2fae57292379c9d15c62eb = (Iedd960a21b1c08b4a5293cff200218b3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I51a2b9abfab582408aeea3130d1e8334;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00038_00002_U (
.flogtanh_sel( If9722c28747df3a59b0ecf8200907e98[flogtanh_SEL-1:0]),
.flogtanh( Icddd184270ffda26b803956883400ad0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id1bc8bf048edb72a3564f864e8fb8671  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icddd184270ffda26b803956883400ad0 };
assign Ibe502ebbb366f54a8f8fda4e361308e3 = (If9722c28747df3a59b0ecf8200907e98[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id1bc8bf048edb72a3564f864e8fb8671;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00038_00003_U (
.flogtanh_sel( Ib83df72c8b73a333d0699a8bbbec16be[flogtanh_SEL-1:0]),
.flogtanh( Id3da7061c05091ffc520d4480058e8e9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7aa45db0b1c7bd90b21c438b91070a16  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id3da7061c05091ffc520d4480058e8e9 };
assign Ifce70fefde8f5ea4d2c1857236f66d65 = (Ib83df72c8b73a333d0699a8bbbec16be[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7aa45db0b1c7bd90b21c438b91070a16;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00038_00004_U (
.flogtanh_sel( Ide3798a77f709a9f694523338b081f70[flogtanh_SEL-1:0]),
.flogtanh( Ie63d649228270b34d8ed25e7c4b09883),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4673a5950ad69c59f3cf4001a1dc93d2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie63d649228270b34d8ed25e7c4b09883 };
assign Ice2c390d296e09b117d60905343e9098 = (Ide3798a77f709a9f694523338b081f70[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4673a5950ad69c59f3cf4001a1dc93d2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00038_00005_U (
.flogtanh_sel( I0a9722a805604433562f85c62b168b96[flogtanh_SEL-1:0]),
.flogtanh( I8eed3f7b36c046fff1e41dd52a300d29),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iffb8eaecd6bd058181a4532d83f674a5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8eed3f7b36c046fff1e41dd52a300d29 };
assign I4b94402a53d981e953c21ef316c709b7 = (I0a9722a805604433562f85c62b168b96[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iffb8eaecd6bd058181a4532d83f674a5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00038_00006_U (
.flogtanh_sel( If9480ec13cd538ed03a43e56bd6264a6[flogtanh_SEL-1:0]),
.flogtanh( Iefcebe38e0c2d6d570017e165d70d3b1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0a7e192f836bc8f7c0ea6bd7a66adaa7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iefcebe38e0c2d6d570017e165d70d3b1 };
assign I450c0d6ad5d3b1f18bb28e3a432b5442 = (If9480ec13cd538ed03a43e56bd6264a6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0a7e192f836bc8f7c0ea6bd7a66adaa7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00038_00007_U (
.flogtanh_sel( I433ecf86b7704c5552e5fb5cafe0d529[flogtanh_SEL-1:0]),
.flogtanh( Ia153222350357443978d7426663c3eaa),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic38ac13f1b1f78c5e83379cabf407f5a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia153222350357443978d7426663c3eaa };
assign I2587a5800a5a9ffeabc4dca503e3d964 = (I433ecf86b7704c5552e5fb5cafe0d529[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic38ac13f1b1f78c5e83379cabf407f5a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00039_00000_U (
.flogtanh_sel( I8326f0b2d25139609e2c5e466724f224[flogtanh_SEL-1:0]),
.flogtanh( I06f0fd2d9d46a2fdb4221217ee2496d1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie9b7108feaaa1fd3e2dc5eeba3d6c4e5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I06f0fd2d9d46a2fdb4221217ee2496d1 };
assign I1182655739d7ab5bbe4a6546a5ca36fd = (I8326f0b2d25139609e2c5e466724f224[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie9b7108feaaa1fd3e2dc5eeba3d6c4e5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00039_00001_U (
.flogtanh_sel( Ibbe211d9955cdf2810c9003d1fb78074[flogtanh_SEL-1:0]),
.flogtanh( I9533ff0882ed01409795d7269329fd76),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iab83df9535036f6c0108658ebd03620a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9533ff0882ed01409795d7269329fd76 };
assign I8110a5a62607093b21b7cd088b1d9ee0 = (Ibbe211d9955cdf2810c9003d1fb78074[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iab83df9535036f6c0108658ebd03620a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00039_00002_U (
.flogtanh_sel( If15e950b569a92b590127d0ca6f20a16[flogtanh_SEL-1:0]),
.flogtanh( Ia9eb9821e7dc31c23d7e60839949c1ff),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5dac976084afd52f5b0d21306bcbb511  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia9eb9821e7dc31c23d7e60839949c1ff };
assign I8b611f7c12ddd81de403ba74e212857f = (If15e950b569a92b590127d0ca6f20a16[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5dac976084afd52f5b0d21306bcbb511;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00039_00003_U (
.flogtanh_sel( I03e0532841ba39eb1d4ae823c4de2f7d[flogtanh_SEL-1:0]),
.flogtanh( I3663fc86620d6244a850819bd3ebe72c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I018c59ff182308d3ca739dbe309ba91e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3663fc86620d6244a850819bd3ebe72c };
assign I84a62a133dbceb5a32a7c907f371663d = (I03e0532841ba39eb1d4ae823c4de2f7d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I018c59ff182308d3ca739dbe309ba91e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00039_00004_U (
.flogtanh_sel( I1be81a7b73987ee023e396cec87312d1[flogtanh_SEL-1:0]),
.flogtanh( I11293e7cdeddf352011d46abd6c3bb72),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9a117a38c8db8191f34cfe7a403aa135  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I11293e7cdeddf352011d46abd6c3bb72 };
assign Ia2fc8a1bbc3cb0dd7d89a7f05b04909c = (I1be81a7b73987ee023e396cec87312d1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9a117a38c8db8191f34cfe7a403aa135;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00039_00005_U (
.flogtanh_sel( I4ce1a767a78673590c4074f3f03bad8d[flogtanh_SEL-1:0]),
.flogtanh( Ic9339e415d0f756e34bcd930de63ad87),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I60d5a8f56d1f22d535a53bbba3049a56  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic9339e415d0f756e34bcd930de63ad87 };
assign I2a3eb42a4402e873d081f94a14a99c20 = (I4ce1a767a78673590c4074f3f03bad8d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I60d5a8f56d1f22d535a53bbba3049a56;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00039_00006_U (
.flogtanh_sel( I57806bb7da625881e68ae315543f70d6[flogtanh_SEL-1:0]),
.flogtanh( Icf109f65e24d3a23ecad9e7d4cc54dc1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I270d4c8baa595241fcc0060b18749f4f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icf109f65e24d3a23ecad9e7d4cc54dc1 };
assign I58447d6ae49a6be2d043477a06f83df0 = (I57806bb7da625881e68ae315543f70d6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I270d4c8baa595241fcc0060b18749f4f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00039_00007_U (
.flogtanh_sel( I8b0ab476b4790150575abb06bcdce2b3[flogtanh_SEL-1:0]),
.flogtanh( Idf7dd0ff83b2d56693e729a1a375fabb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I765d0dd290e34cee0116f45ce9527117  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idf7dd0ff83b2d56693e729a1a375fabb };
assign I83292bcda4645233d8e8a1dfe8e5f60b = (I8b0ab476b4790150575abb06bcdce2b3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I765d0dd290e34cee0116f45ce9527117;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00040_00000_U (
.flogtanh_sel( I8846a8961b7d557df4fc62dada679c33[flogtanh_SEL-1:0]),
.flogtanh( I312a248019372261c0959cdc9378ec93),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9ef68d76daf35fa29a0c4168baf64516  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I312a248019372261c0959cdc9378ec93 };
assign Ic5e0a84cf1a2ef907b2456559ea26c75 = (I8846a8961b7d557df4fc62dada679c33[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9ef68d76daf35fa29a0c4168baf64516;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00040_00001_U (
.flogtanh_sel( I7909a0f96a92e93f95023cddc742a5eb[flogtanh_SEL-1:0]),
.flogtanh( I8e311b9891dda272762da2c640019e8c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icc9faf407342c704a8f33b49c1ad8063  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8e311b9891dda272762da2c640019e8c };
assign I2cefbf897bb7f6f67ca500727e85c683 = (I7909a0f96a92e93f95023cddc742a5eb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icc9faf407342c704a8f33b49c1ad8063;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00040_00002_U (
.flogtanh_sel( I43ac4857544c0fb79d04e850435ef673[flogtanh_SEL-1:0]),
.flogtanh( I1874dd9f7c0a93310873173561402912),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibdfcf91a62d88e9b8d011a22c8100106  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1874dd9f7c0a93310873173561402912 };
assign If47be2ca4617a426258c51f8d977ba3f = (I43ac4857544c0fb79d04e850435ef673[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibdfcf91a62d88e9b8d011a22c8100106;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00040_00003_U (
.flogtanh_sel( Ia6dfa47c465325c1d9fb9b9c5ce08f01[flogtanh_SEL-1:0]),
.flogtanh( I04adb3964e739a106098a6c4d2f49e94),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6ff243d4d70ead40034f55f7b0c49557  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I04adb3964e739a106098a6c4d2f49e94 };
assign I7c68e0ae30efc4ca4d68b6047119c6c3 = (Ia6dfa47c465325c1d9fb9b9c5ce08f01[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6ff243d4d70ead40034f55f7b0c49557;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00040_00004_U (
.flogtanh_sel( I2e9eda5bea0cc3d88359ce8a7a82f21f[flogtanh_SEL-1:0]),
.flogtanh( I9135b709c3c802a42c7186087b5664cc),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6fe27a172bfa6cd64ae70b8a22f66e4a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9135b709c3c802a42c7186087b5664cc };
assign Iccca1936f4c1c9496205e77b588e9985 = (I2e9eda5bea0cc3d88359ce8a7a82f21f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6fe27a172bfa6cd64ae70b8a22f66e4a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00040_00005_U (
.flogtanh_sel( I53ec2486418e41b2ccfa8fd82777eaf0[flogtanh_SEL-1:0]),
.flogtanh( Ia236dfe34ff4938456d76f787d2db945),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I20b96db33a7f876f9b37e0dd13d39630  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia236dfe34ff4938456d76f787d2db945 };
assign I59d4567d3355fdae5660a1364d1b8d00 = (I53ec2486418e41b2ccfa8fd82777eaf0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I20b96db33a7f876f9b37e0dd13d39630;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00040_00006_U (
.flogtanh_sel( I18387c05cef21970ecbc39c20a87aafb[flogtanh_SEL-1:0]),
.flogtanh( I41c98bae5fbdb31bac0913930573e80c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic1c711155cf28a3491f52352d5fbd05a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I41c98bae5fbdb31bac0913930573e80c };
assign I4600963866dcb9bbea2515c805f885cb = (I18387c05cef21970ecbc39c20a87aafb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic1c711155cf28a3491f52352d5fbd05a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00040_00007_U (
.flogtanh_sel( I2b23eae78cb925008ad59f45e80e165b[flogtanh_SEL-1:0]),
.flogtanh( I226befd72285893998aca87fe34d9aaf),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic99fca70349dfdfdbec515ab163ad20f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I226befd72285893998aca87fe34d9aaf };
assign If26d90629e70c5a871e6f5b14471b8cf = (I2b23eae78cb925008ad59f45e80e165b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic99fca70349dfdfdbec515ab163ad20f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00040_00008_U (
.flogtanh_sel( Ic69eb7677638a90b7a54389d47be46de[flogtanh_SEL-1:0]),
.flogtanh( I20ab7c6174af39aee99492f704b2748c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I71db278548cbf6a478f5f2d7de410dc9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I20ab7c6174af39aee99492f704b2748c };
assign Iedb9bb14951bf67bc8865b0983490c14 = (Ic69eb7677638a90b7a54389d47be46de[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I71db278548cbf6a478f5f2d7de410dc9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00041_00000_U (
.flogtanh_sel( I8cb9a216f4da7c27f678386cb214c59d[flogtanh_SEL-1:0]),
.flogtanh( I0a1c5724ffa14df653142a1f8bcf44a4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I67f75dfd3165ca969119ededc4c25b1d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0a1c5724ffa14df653142a1f8bcf44a4 };
assign I6a3854ed571e8c262aa3ec377c247778 = (I8cb9a216f4da7c27f678386cb214c59d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I67f75dfd3165ca969119ededc4c25b1d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00041_00001_U (
.flogtanh_sel( I48cb720a6323697084ac3bbd8fcadfcb[flogtanh_SEL-1:0]),
.flogtanh( I481973954b81accf069dd80830fba3bc),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia4f05220e30b257689f831feaa0125e9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I481973954b81accf069dd80830fba3bc };
assign I05028975b49ec0c089bd981696f85a8b = (I48cb720a6323697084ac3bbd8fcadfcb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia4f05220e30b257689f831feaa0125e9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00041_00002_U (
.flogtanh_sel( Ib8dc3c1885c92cdcce7fcb58d65d03e7[flogtanh_SEL-1:0]),
.flogtanh( Ia6825c3edc9d2a6832db7a7d684faf98),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieeaf2a662a0f9295b3c3d6454f731098  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia6825c3edc9d2a6832db7a7d684faf98 };
assign Ife732309efcc740cfff5c747aab2e3d6 = (Ib8dc3c1885c92cdcce7fcb58d65d03e7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieeaf2a662a0f9295b3c3d6454f731098;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00041_00003_U (
.flogtanh_sel( Ic3aa51a5c758405fa6e2dbed707555b2[flogtanh_SEL-1:0]),
.flogtanh( I5c964036207f47629302e282d56fef7b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id7e4f0f2bded6e1d39467d074348b324  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5c964036207f47629302e282d56fef7b };
assign Idcef10a0465614cf38e0d6f503b5174a = (Ic3aa51a5c758405fa6e2dbed707555b2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id7e4f0f2bded6e1d39467d074348b324;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00041_00004_U (
.flogtanh_sel( I4d418179c859feb8bc7d750416bb1004[flogtanh_SEL-1:0]),
.flogtanh( I00b74ed4d6730b37c6fbfd42dee42584),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4c556e88e578d8f5d2d529b33a00b9eb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I00b74ed4d6730b37c6fbfd42dee42584 };
assign Ibd4aaf02982068ffbfd1b8b3795d9217 = (I4d418179c859feb8bc7d750416bb1004[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4c556e88e578d8f5d2d529b33a00b9eb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00041_00005_U (
.flogtanh_sel( If207b2adc6f668f85cb76bf54673fe18[flogtanh_SEL-1:0]),
.flogtanh( I0345fc4a507f9e3be3e1d46b71693de1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I25facb36e0360a4ca4ac5803101984c7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0345fc4a507f9e3be3e1d46b71693de1 };
assign I788c64785b992c675fe348a1fa181525 = (If207b2adc6f668f85cb76bf54673fe18[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I25facb36e0360a4ca4ac5803101984c7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00041_00006_U (
.flogtanh_sel( Ib08b8067ea75e210e83526ca4a37217e[flogtanh_SEL-1:0]),
.flogtanh( I9f0735c1cf5d1af7c82a251ef4886f9c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iab18a2d81fc63ba2b35df1cdf08621af  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9f0735c1cf5d1af7c82a251ef4886f9c };
assign Ib235af5b28d56f24372d3f0af816f2c2 = (Ib08b8067ea75e210e83526ca4a37217e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iab18a2d81fc63ba2b35df1cdf08621af;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00041_00007_U (
.flogtanh_sel( I95b30f641cbf7bec1886643c4468017d[flogtanh_SEL-1:0]),
.flogtanh( I861cf5dffb18c84953013dc4026bd08a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icd609cdfdfa1ecb62bba040a015b8de5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I861cf5dffb18c84953013dc4026bd08a };
assign I4c03a6569d1b954d088053e38827e811 = (I95b30f641cbf7bec1886643c4468017d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icd609cdfdfa1ecb62bba040a015b8de5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00041_00008_U (
.flogtanh_sel( I1978531a6f8d1d25ee6d404025ec4753[flogtanh_SEL-1:0]),
.flogtanh( I19722ceada71cc9cc06edde39142ff17),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I00c895c62ee2842ad86d01beab41e900  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I19722ceada71cc9cc06edde39142ff17 };
assign Idda26504e422367082caeafbb29871f9 = (I1978531a6f8d1d25ee6d404025ec4753[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I00c895c62ee2842ad86d01beab41e900;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00042_00000_U (
.flogtanh_sel( I6c9698ba88db16b8d22ccebd58cc541d[flogtanh_SEL-1:0]),
.flogtanh( Id8349128e2c391df008828494da928c6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idd279726169e173c111b7c490a2c4037  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id8349128e2c391df008828494da928c6 };
assign I195c3a82123142d509886ee37dc6fc98 = (I6c9698ba88db16b8d22ccebd58cc541d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idd279726169e173c111b7c490a2c4037;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00042_00001_U (
.flogtanh_sel( I0d8ac5e09b200a55bf5ba6f834cc9174[flogtanh_SEL-1:0]),
.flogtanh( I27209805df490a07f1726875a7b69922),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I125a005c7f9d37d5365496513fef1893  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I27209805df490a07f1726875a7b69922 };
assign I1abb512ca0383c9e7104418e07281841 = (I0d8ac5e09b200a55bf5ba6f834cc9174[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I125a005c7f9d37d5365496513fef1893;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00042_00002_U (
.flogtanh_sel( Ib58b7d3d77a54ff1a180c6fa5f1400e6[flogtanh_SEL-1:0]),
.flogtanh( I7532c1f0624a2d5a94321c89c73e38df),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I62802ceb2a05dc315e7137f31590cc72  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7532c1f0624a2d5a94321c89c73e38df };
assign I00ff1331b1900bb031ee81d2a58c1bd5 = (Ib58b7d3d77a54ff1a180c6fa5f1400e6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I62802ceb2a05dc315e7137f31590cc72;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00042_00003_U (
.flogtanh_sel( Icf6b990098b7ab91800bfcf1e643153c[flogtanh_SEL-1:0]),
.flogtanh( Ife892846e66e2522c06b170811a11ada),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5b0fda1e3b1829738e08b1de1d934a1c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ife892846e66e2522c06b170811a11ada };
assign If65eb5e743a7b1878fb232ef2fe13cb0 = (Icf6b990098b7ab91800bfcf1e643153c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5b0fda1e3b1829738e08b1de1d934a1c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00042_00004_U (
.flogtanh_sel( Ie4308b9ac6fb6de9329ba02b1eeb0e8a[flogtanh_SEL-1:0]),
.flogtanh( Ib905ede2830f7e3c8cf993075f07345c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0f86873fc1d12c964a3757bec70ad780  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib905ede2830f7e3c8cf993075f07345c };
assign I24ae7de3549a84f4f88f561b6017b7a8 = (Ie4308b9ac6fb6de9329ba02b1eeb0e8a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0f86873fc1d12c964a3757bec70ad780;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00042_00005_U (
.flogtanh_sel( I01d4f02a356c51d7e4e1993de0d8eebd[flogtanh_SEL-1:0]),
.flogtanh( Ibf169f844d9e00eca8f3821ddc952ef0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6f41f58cfeab93cd06c32cd2537426dd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibf169f844d9e00eca8f3821ddc952ef0 };
assign I449c77140475475b138d839a74078337 = (I01d4f02a356c51d7e4e1993de0d8eebd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6f41f58cfeab93cd06c32cd2537426dd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00042_00006_U (
.flogtanh_sel( I36c351e3641b01cc43e1dd5de0a649e5[flogtanh_SEL-1:0]),
.flogtanh( I3137f75629e72f78abdac088e18608d5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibf529f3a5b5f9d44d2e072b2cfb0c987  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3137f75629e72f78abdac088e18608d5 };
assign Ia9e102d8679943c079f16c0228f0f0d1 = (I36c351e3641b01cc43e1dd5de0a649e5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibf529f3a5b5f9d44d2e072b2cfb0c987;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00042_00007_U (
.flogtanh_sel( I4fc983e94c5b8f7bafca61fb0d351c08[flogtanh_SEL-1:0]),
.flogtanh( I8fbcabc2f5c30fcf1c5b46de5dfe887d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I189af406b34e849a5700be4ea8d7a22b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8fbcabc2f5c30fcf1c5b46de5dfe887d };
assign Ibf1c9d86665f696d91c554db748ff42b = (I4fc983e94c5b8f7bafca61fb0d351c08[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I189af406b34e849a5700be4ea8d7a22b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00042_00008_U (
.flogtanh_sel( I1fcb82fdf96cda14a55fa6358cb62c1e[flogtanh_SEL-1:0]),
.flogtanh( Ie7acfb624aa6242b558481350c85fda3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2e6d80f71d9e42ef5e32d8e43c9ad77e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie7acfb624aa6242b558481350c85fda3 };
assign Ieb0336a1974a2aec0966f4f59f460802 = (I1fcb82fdf96cda14a55fa6358cb62c1e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2e6d80f71d9e42ef5e32d8e43c9ad77e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00043_00000_U (
.flogtanh_sel( I665e54ea6bdca483149d3b7f3ee42a2b[flogtanh_SEL-1:0]),
.flogtanh( I11e0b915338d5d649c800455b9a7695f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8a8379ec2c6c9c360b2c32c34e63902d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I11e0b915338d5d649c800455b9a7695f };
assign Ic0819ccefe784a6379716b3633ae0196 = (I665e54ea6bdca483149d3b7f3ee42a2b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8a8379ec2c6c9c360b2c32c34e63902d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00043_00001_U (
.flogtanh_sel( I925df2307b5af6d1b166e5435641d3bd[flogtanh_SEL-1:0]),
.flogtanh( Ia9e4e68dcd3d0281decde939eed0c3bd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic89ee3a7462610019feee4023e1ab63e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia9e4e68dcd3d0281decde939eed0c3bd };
assign I0c4bbd1827b1859caabb067e864ce4b3 = (I925df2307b5af6d1b166e5435641d3bd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic89ee3a7462610019feee4023e1ab63e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00043_00002_U (
.flogtanh_sel( I9b14f48aa357d09e460a445da86cdf89[flogtanh_SEL-1:0]),
.flogtanh( Id508f63a381fc565a28fe4e662b33efb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I49b0d9feed7042dc0551398d48b36f7f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id508f63a381fc565a28fe4e662b33efb };
assign I004c98da87996b77b5761d366210f782 = (I9b14f48aa357d09e460a445da86cdf89[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I49b0d9feed7042dc0551398d48b36f7f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00043_00003_U (
.flogtanh_sel( I78e94ecb6c92fa8ee24edaff33b6f82d[flogtanh_SEL-1:0]),
.flogtanh( I33582dc83370e68b0ae7b22b553276b4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icfbd9d5dfe741fd84977d13887a54dee  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I33582dc83370e68b0ae7b22b553276b4 };
assign Ia457938da4efe847cb06f645f2a54a52 = (I78e94ecb6c92fa8ee24edaff33b6f82d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icfbd9d5dfe741fd84977d13887a54dee;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00043_00004_U (
.flogtanh_sel( I5ebeb9ce5adee72a7c9527ea6d3a3028[flogtanh_SEL-1:0]),
.flogtanh( I8aeca996ad6820edcc6fcbaa8a0f15ce),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib2b669872ca023cf13754a529eab5ad5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8aeca996ad6820edcc6fcbaa8a0f15ce };
assign I7e0474089ebc1c34747be1bc17a81d72 = (I5ebeb9ce5adee72a7c9527ea6d3a3028[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib2b669872ca023cf13754a529eab5ad5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00043_00005_U (
.flogtanh_sel( I90d7b28ec09142ca8086836fc0c5ea0d[flogtanh_SEL-1:0]),
.flogtanh( Ica86e8037319b868c8cb89f3cb02b136),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ife9a683c5c06abb98e9a9da56244cadf  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ica86e8037319b868c8cb89f3cb02b136 };
assign Ib0b46b99e61d724ae664d9d1fec1e29f = (I90d7b28ec09142ca8086836fc0c5ea0d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ife9a683c5c06abb98e9a9da56244cadf;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00043_00006_U (
.flogtanh_sel( I27d9985415e6d0b117e5a4c2863aa7f8[flogtanh_SEL-1:0]),
.flogtanh( Ia95013b19d9fc12d19ff9924007113d4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic2a2da3827248989cad50ff9fcc8822e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia95013b19d9fc12d19ff9924007113d4 };
assign I56d1025271f1f7704a40dd7f0df02b0b = (I27d9985415e6d0b117e5a4c2863aa7f8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic2a2da3827248989cad50ff9fcc8822e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00043_00007_U (
.flogtanh_sel( Idf9b563e5d10c2bdbcc07e81d74467eb[flogtanh_SEL-1:0]),
.flogtanh( Ifcf979b713b014f22c1c8ce1d42132c2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifcbb960ba610a378b0472f005bea218a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifcf979b713b014f22c1c8ce1d42132c2 };
assign I72c2256ba47cf03f95143df8f741fd83 = (Idf9b563e5d10c2bdbcc07e81d74467eb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifcbb960ba610a378b0472f005bea218a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00043_00008_U (
.flogtanh_sel( Ie351922194483938302ff6cafc477e4a[flogtanh_SEL-1:0]),
.flogtanh( I973b3306021532f286cf248084398c26),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9527b33b0941a515601b7fb75c0eba34  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I973b3306021532f286cf248084398c26 };
assign I733c3fa4d84e5680792b16a70bb1a51d = (Ie351922194483938302ff6cafc477e4a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9527b33b0941a515601b7fb75c0eba34;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00000_U (
.flogtanh_sel( Ifb2da5faf236ca8636677bc1dc35c4db[flogtanh_SEL-1:0]),
.flogtanh( Iea7940bb396d1a436f56806fc533edee),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia65e331b9f0ec80ee7860b2c4a6c1e55  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iea7940bb396d1a436f56806fc533edee };
assign If367d63311c96726517240de13bd2a4b = (Ifb2da5faf236ca8636677bc1dc35c4db[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia65e331b9f0ec80ee7860b2c4a6c1e55;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00001_U (
.flogtanh_sel( Ie15825d216685ae241b528fa9c158ff3[flogtanh_SEL-1:0]),
.flogtanh( Ied55045b003302c294591a8d2a6a39fd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2cbdbbf07d938e2f4847fdf594a010c8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ied55045b003302c294591a8d2a6a39fd };
assign Icc6d895d943e14f2801c22e79ce190e8 = (Ie15825d216685ae241b528fa9c158ff3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2cbdbbf07d938e2f4847fdf594a010c8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00002_U (
.flogtanh_sel( Id92c2d8bc61245c0c8e40bec2424c3c8[flogtanh_SEL-1:0]),
.flogtanh( Ib64e948413d5dce1d9309fe95c0919ab),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I260ec6308196983b8aeaddcac953709d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib64e948413d5dce1d9309fe95c0919ab };
assign Ieb664ac9be65fba2e25960141f7fb4b6 = (Id92c2d8bc61245c0c8e40bec2424c3c8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I260ec6308196983b8aeaddcac953709d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00003_U (
.flogtanh_sel( Icd9fd8d7114b6e894dbee493b6797df6[flogtanh_SEL-1:0]),
.flogtanh( I682fe6c6c621db5dd867574e8573d8ed),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I456482f0ce8cb6c76d2b19b69cd0f4fc  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I682fe6c6c621db5dd867574e8573d8ed };
assign I66071f20991b414140869a2e3b750471 = (Icd9fd8d7114b6e894dbee493b6797df6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I456482f0ce8cb6c76d2b19b69cd0f4fc;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00004_U (
.flogtanh_sel( I29ff688c085f2b18e7a3af969f18af76[flogtanh_SEL-1:0]),
.flogtanh( I508b57f6ebc45eb70aa7b114096a7d12),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie9d6a3cf41e366e12a6d90a61163fb48  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I508b57f6ebc45eb70aa7b114096a7d12 };
assign Iffeefa89a2ba7d032db5db64cbf05e20 = (I29ff688c085f2b18e7a3af969f18af76[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie9d6a3cf41e366e12a6d90a61163fb48;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00005_U (
.flogtanh_sel( I6d56db9fcfe69dfcd747521a1ff62297[flogtanh_SEL-1:0]),
.flogtanh( I8e82b8914260669ed1d88a690467a7b4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieb526cf88e7ac70a26f05c0f56d37c91  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8e82b8914260669ed1d88a690467a7b4 };
assign I9ab3cea6ee8d8473221da21bae06066b = (I6d56db9fcfe69dfcd747521a1ff62297[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieb526cf88e7ac70a26f05c0f56d37c91;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00006_U (
.flogtanh_sel( I2f17f7c79a0118b39a63894917c6affa[flogtanh_SEL-1:0]),
.flogtanh( I525feb94b558fb4bb8db8eead9f05afa),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If4ccf2222e01f9418f342054b342412f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I525feb94b558fb4bb8db8eead9f05afa };
assign I3403ce6e697b523a9f441d8fd5e2d420 = (I2f17f7c79a0118b39a63894917c6affa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If4ccf2222e01f9418f342054b342412f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00007_U (
.flogtanh_sel( I7350af5d5ee09ad28c459e3674a829ab[flogtanh_SEL-1:0]),
.flogtanh( Ie5e4cf2b42054822a9091f5ef67cd968),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0875d93243187e274b27f729a86dd9fa  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie5e4cf2b42054822a9091f5ef67cd968 };
assign Ia98a70144e466b356d2998948dc4b602 = (I7350af5d5ee09ad28c459e3674a829ab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0875d93243187e274b27f729a86dd9fa;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00008_U (
.flogtanh_sel( I67b6415c5135e3d6a41d56d98d3f8315[flogtanh_SEL-1:0]),
.flogtanh( I0d08d26e31c8b69ed8c089cdcd055a50),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibd4f6d59420fe37742ef3ae1f22c152c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0d08d26e31c8b69ed8c089cdcd055a50 };
assign Ie4ca0836695d951ee09622892ee35928 = (I67b6415c5135e3d6a41d56d98d3f8315[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibd4f6d59420fe37742ef3ae1f22c152c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00009_U (
.flogtanh_sel( I4a6fffd8bb7244599383f2aa3a1c8916[flogtanh_SEL-1:0]),
.flogtanh( I877f44c880a781381bfa8a8f8471d697),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2f726cba2feffeaeeadff790c6909402  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I877f44c880a781381bfa8a8f8471d697 };
assign I485a48b4ff4da08f977425fd10e6d392 = (I4a6fffd8bb7244599383f2aa3a1c8916[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2f726cba2feffeaeeadff790c6909402;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00010_U (
.flogtanh_sel( I7dbcd21016231546b76aab175cac9f74[flogtanh_SEL-1:0]),
.flogtanh( I7fc78273dc765cf1c03b3c1a043b35f8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id8d5b7c74ba1b051e3e4eb87d812e028  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7fc78273dc765cf1c03b3c1a043b35f8 };
assign Ie8c79e6a5378808c0ead5a4b24319ce9 = (I7dbcd21016231546b76aab175cac9f74[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id8d5b7c74ba1b051e3e4eb87d812e028;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00011_U (
.flogtanh_sel( I9aeff3dc44ed0d0f32518590a900dcc9[flogtanh_SEL-1:0]),
.flogtanh( Ie67275a4b3fdc050f0f6e7ac7d1eebfc),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2c853ac0b4a3ac567a4db08ba5e9e26d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie67275a4b3fdc050f0f6e7ac7d1eebfc };
assign I9ca81c841a75a9ac242835956509e0fe = (I9aeff3dc44ed0d0f32518590a900dcc9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2c853ac0b4a3ac567a4db08ba5e9e26d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00012_U (
.flogtanh_sel( I988b7d5d56d22d2c77c5c8c125129a50[flogtanh_SEL-1:0]),
.flogtanh( I41f9acc96650353174155a5f378d5cc5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifa2b0aa146869b9f6238969c5649acc7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I41f9acc96650353174155a5f378d5cc5 };
assign Id50f18f642f3b00ffa34986f78a0eae6 = (I988b7d5d56d22d2c77c5c8c125129a50[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifa2b0aa146869b9f6238969c5649acc7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00013_U (
.flogtanh_sel( Iff35cd97f2a6d37a7861b9cc1a655ef5[flogtanh_SEL-1:0]),
.flogtanh( I0d73c905b2ed777acd71d560928dcf0b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib4322244b363748db4a0543933452669  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0d73c905b2ed777acd71d560928dcf0b };
assign I75838ca09e301b8e1301cbf603a1f8c2 = (Iff35cd97f2a6d37a7861b9cc1a655ef5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib4322244b363748db4a0543933452669;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00014_U (
.flogtanh_sel( Ifb3f2a1bedfe41c73d198046a2a3f177[flogtanh_SEL-1:0]),
.flogtanh( I2b6b1c25caf8b00d19ccc98156a8ca2b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idbd452a90ce7a7c82d5d2d7f57fbd72c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2b6b1c25caf8b00d19ccc98156a8ca2b };
assign Id968b34075e351ab01d65abcb4ed8cca = (Ifb3f2a1bedfe41c73d198046a2a3f177[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idbd452a90ce7a7c82d5d2d7f57fbd72c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00044_00015_U (
.flogtanh_sel( I37ddc6ccbc188a3eb8c33a501de820be[flogtanh_SEL-1:0]),
.flogtanh( I28ea2b207bcd3518a85ff150466a6a08),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I28ceab58b644f619bb359f153087cb9b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I28ea2b207bcd3518a85ff150466a6a08 };
assign I84da4ce7441e132e775167c1cd81dbe5 = (I37ddc6ccbc188a3eb8c33a501de820be[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I28ceab58b644f619bb359f153087cb9b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00000_U (
.flogtanh_sel( Ica608f1136da397e2ab61bd4a5d83201[flogtanh_SEL-1:0]),
.flogtanh( I7d0a1c64b2e85e1bf0bf99423321466b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaf75fbdcad76103a769669bc20d0c5b7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7d0a1c64b2e85e1bf0bf99423321466b };
assign If19dc22d45cc4664c85a043ec4c00617 = (Ica608f1136da397e2ab61bd4a5d83201[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaf75fbdcad76103a769669bc20d0c5b7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00001_U (
.flogtanh_sel( I80636a3df4541bf29780bcb4d0ee48f9[flogtanh_SEL-1:0]),
.flogtanh( I3b9b9b41b54ff194314b572a15daf606),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4a34573ee0f529e4088f1b5969eee325  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3b9b9b41b54ff194314b572a15daf606 };
assign Ibf482db0f5058be72061267c42ebc292 = (I80636a3df4541bf29780bcb4d0ee48f9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4a34573ee0f529e4088f1b5969eee325;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00002_U (
.flogtanh_sel( I9ad99d544187db3cc7090b92c9933a31[flogtanh_SEL-1:0]),
.flogtanh( Ic914f847e623d9c52e2d9ae5076c21c3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0602ea657e22176e268c3f005b327c5f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic914f847e623d9c52e2d9ae5076c21c3 };
assign I6d2dbb953a58b91dafa7f0d34d41bdc3 = (I9ad99d544187db3cc7090b92c9933a31[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0602ea657e22176e268c3f005b327c5f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00003_U (
.flogtanh_sel( Iaa8a2b6fcd469869efcf0b75ca38e68f[flogtanh_SEL-1:0]),
.flogtanh( I46fc20938dd554b23b5af5f7c3e39480),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I48ef1d4bacb30b7602392e7298e88c40  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I46fc20938dd554b23b5af5f7c3e39480 };
assign Ib393146d81d3cf031466543311cee2ad = (Iaa8a2b6fcd469869efcf0b75ca38e68f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I48ef1d4bacb30b7602392e7298e88c40;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00004_U (
.flogtanh_sel( I9a171d2d8eee362a0073ab7b139d3037[flogtanh_SEL-1:0]),
.flogtanh( I1fa8b37b4697ae60cf399285d9524b8d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I36272af5470aa53e7c61cbc896f26290  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1fa8b37b4697ae60cf399285d9524b8d };
assign I42564ec6a794ea803795f0b5b3523a93 = (I9a171d2d8eee362a0073ab7b139d3037[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I36272af5470aa53e7c61cbc896f26290;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00005_U (
.flogtanh_sel( I84cdcba86bc5991feb391003cd7be40b[flogtanh_SEL-1:0]),
.flogtanh( I66c8261df769288836e188ecb32b6dc6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I146bdc684c432e98b5e1c3b274f3272c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I66c8261df769288836e188ecb32b6dc6 };
assign I4a0033a180d7edce81fcfef603532e28 = (I84cdcba86bc5991feb391003cd7be40b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I146bdc684c432e98b5e1c3b274f3272c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00006_U (
.flogtanh_sel( If9e5c3a848acce5daf570458f78f6aad[flogtanh_SEL-1:0]),
.flogtanh( I267714c8a5aa14bae9c74da272a60aa5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I723e72d69796cee0c174c82c2514cd7c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I267714c8a5aa14bae9c74da272a60aa5 };
assign Ic7a21921e2716fba55aad2e351f4498a = (If9e5c3a848acce5daf570458f78f6aad[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I723e72d69796cee0c174c82c2514cd7c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00007_U (
.flogtanh_sel( I73247d4348333f67a491fc607b15af0e[flogtanh_SEL-1:0]),
.flogtanh( I47a34c8d2174c12f96041e82ad835db2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I305b258a587eb0f55a48679ab7ddcf91  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I47a34c8d2174c12f96041e82ad835db2 };
assign I9a3f0b4867087790c78f674b719dbf7b = (I73247d4348333f67a491fc607b15af0e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I305b258a587eb0f55a48679ab7ddcf91;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00008_U (
.flogtanh_sel( I021c745eee4b85a2cd91d9d8d2b18b2c[flogtanh_SEL-1:0]),
.flogtanh( If99ca487495a015063fd8dc54ae596aa),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia8a328c524c386c6008d76d6c920ab03  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If99ca487495a015063fd8dc54ae596aa };
assign I138f008a6206a1067bb0e22ce3d90990 = (I021c745eee4b85a2cd91d9d8d2b18b2c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia8a328c524c386c6008d76d6c920ab03;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00009_U (
.flogtanh_sel( I1381c0a0bd28b1c5542992084635b355[flogtanh_SEL-1:0]),
.flogtanh( I1043f1b92b49a8c304a23c0b5c615def),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5269f5ff21c0c874811b85f6a028c113  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1043f1b92b49a8c304a23c0b5c615def };
assign I48ad9b737892d7c49340ed679f46e034 = (I1381c0a0bd28b1c5542992084635b355[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5269f5ff21c0c874811b85f6a028c113;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00010_U (
.flogtanh_sel( Ie74eeddc21428254a8fc4c3e293b5eb7[flogtanh_SEL-1:0]),
.flogtanh( Icafa102383ef33455236ba268b1b7460),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I93671d398af3e4f197eb71233121de97  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icafa102383ef33455236ba268b1b7460 };
assign I04a9c9765fd468a7e841577f09fc287b = (Ie74eeddc21428254a8fc4c3e293b5eb7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I93671d398af3e4f197eb71233121de97;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00011_U (
.flogtanh_sel( Ib1d0f94258b45de4bfe610086d8990c5[flogtanh_SEL-1:0]),
.flogtanh( I677fca8017154fed3e6cd54362e829db),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia26b08bdae3e484e917194c100e1763d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I677fca8017154fed3e6cd54362e829db };
assign I7b929c228c865112f00bc6b4dcc95b52 = (Ib1d0f94258b45de4bfe610086d8990c5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia26b08bdae3e484e917194c100e1763d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00012_U (
.flogtanh_sel( I138d6d5d60df37870cdbb1d9c51a94af[flogtanh_SEL-1:0]),
.flogtanh( I826fe051a6b09d5cacf712431ce89b7c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9fa2896c4dbd25ed089fce8d5ce372b2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I826fe051a6b09d5cacf712431ce89b7c };
assign I2b54a135e59945901e9c11580a29ee3d = (I138d6d5d60df37870cdbb1d9c51a94af[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9fa2896c4dbd25ed089fce8d5ce372b2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00013_U (
.flogtanh_sel( I706378735e63e15c8d5395446ea41db8[flogtanh_SEL-1:0]),
.flogtanh( I23f781ebfa449cec7975b94179d72259),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1e4586148b049d4493e1cafe947c3983  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I23f781ebfa449cec7975b94179d72259 };
assign I566221060f06e724676ec9bec861d7de = (I706378735e63e15c8d5395446ea41db8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1e4586148b049d4493e1cafe947c3983;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00014_U (
.flogtanh_sel( If8680a7fc4f5532a660006bf4ca6a66e[flogtanh_SEL-1:0]),
.flogtanh( Ia383b5dc3b7ce1bc7987926535639668),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I375aeddea735459513ef97aec26fc8d1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia383b5dc3b7ce1bc7987926535639668 };
assign Icd9a876a0feb16ea62bcad5be2004dac = (If8680a7fc4f5532a660006bf4ca6a66e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I375aeddea735459513ef97aec26fc8d1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00045_00015_U (
.flogtanh_sel( Ic59d1ff3051a95166c3c2d5a2881221b[flogtanh_SEL-1:0]),
.flogtanh( I40ae857caffae41564c2ecb0c7e9777b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I683f128be784d4e752ea5881c1d483a8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I40ae857caffae41564c2ecb0c7e9777b };
assign I8f8273c4cb2a9ace8a09847efd4bdec7 = (Ic59d1ff3051a95166c3c2d5a2881221b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I683f128be784d4e752ea5881c1d483a8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00000_U (
.flogtanh_sel( I54a551af28c505601cdfaf8faaa94afb[flogtanh_SEL-1:0]),
.flogtanh( I569d56a2673a104f3050d851d767af8a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iacd3b2128fa021305b3de888d7612cf8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I569d56a2673a104f3050d851d767af8a };
assign I96ef4b631a7f63e19f67f3920685f0e6 = (I54a551af28c505601cdfaf8faaa94afb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iacd3b2128fa021305b3de888d7612cf8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00001_U (
.flogtanh_sel( I6a3124c03eb83d41c16704133bd1cfde[flogtanh_SEL-1:0]),
.flogtanh( I2022005072d2979dae84b6e4491a3ce2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0976b3262637cf38babc31162e3f6cea  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2022005072d2979dae84b6e4491a3ce2 };
assign I9e2de71442b8f504358e582087a6d19f = (I6a3124c03eb83d41c16704133bd1cfde[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0976b3262637cf38babc31162e3f6cea;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00002_U (
.flogtanh_sel( Ie9ee27b9761af611ab96f0010abd47a3[flogtanh_SEL-1:0]),
.flogtanh( I98524ad028e4d832ebbcd92956dac08c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I484113b853de9a5684592b8318430da2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I98524ad028e4d832ebbcd92956dac08c };
assign I1fb13d7500f5ac3821c424bd3688cf4e = (Ie9ee27b9761af611ab96f0010abd47a3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I484113b853de9a5684592b8318430da2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00003_U (
.flogtanh_sel( I305436919f84066a22ab1417ebabd737[flogtanh_SEL-1:0]),
.flogtanh( I4d24e2ba47093eee6669f537374ecce7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4b4a443a54b030b20a3e86ba0f63c1ee  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4d24e2ba47093eee6669f537374ecce7 };
assign I2aabda12ff89e708d04b4399472b5203 = (I305436919f84066a22ab1417ebabd737[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4b4a443a54b030b20a3e86ba0f63c1ee;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00004_U (
.flogtanh_sel( I78e63717f436493b756efa32d66cdefd[flogtanh_SEL-1:0]),
.flogtanh( I227232e7189020459c16b3413e881b80),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifb32581537c4402e5345932d83e1388f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I227232e7189020459c16b3413e881b80 };
assign I8c733a5d394e6b8d045eede5cc7451f6 = (I78e63717f436493b756efa32d66cdefd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifb32581537c4402e5345932d83e1388f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00005_U (
.flogtanh_sel( Ic965ba971642db19ca773eb68dc0b9bf[flogtanh_SEL-1:0]),
.flogtanh( If4359aebd4cc66c75cf2a44f681ccc72),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib032b0c1073c1a3689b8f70a8a1f94b5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If4359aebd4cc66c75cf2a44f681ccc72 };
assign I4f45dd50d2825ab338b8a2a8264096c0 = (Ic965ba971642db19ca773eb68dc0b9bf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib032b0c1073c1a3689b8f70a8a1f94b5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00006_U (
.flogtanh_sel( I579480a66a5f6331fb46de13090ce888[flogtanh_SEL-1:0]),
.flogtanh( I8d2e10b8c474f1a915825ec78072ad56),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3ac6148b8dfcfb0816a01ff2a77b905d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8d2e10b8c474f1a915825ec78072ad56 };
assign Ib45caf6b563d22144be3e9225a99a1cd = (I579480a66a5f6331fb46de13090ce888[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3ac6148b8dfcfb0816a01ff2a77b905d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00007_U (
.flogtanh_sel( I38d78b447217271a63f30f78b424e2ae[flogtanh_SEL-1:0]),
.flogtanh( Ie5b3748f3c81d9eeec767d546b29cbd8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie090d9460623450a9654f24bda1be1f7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie5b3748f3c81d9eeec767d546b29cbd8 };
assign I9d6730140c690037b5ca58aa30103f5b = (I38d78b447217271a63f30f78b424e2ae[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie090d9460623450a9654f24bda1be1f7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00008_U (
.flogtanh_sel( I4c8d7e5474b19a7c63444d0cb6143728[flogtanh_SEL-1:0]),
.flogtanh( Ib764a6d1978dc61cb4499b15c45cb1b4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I42979deb711e94d6a366a9c125277bc7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib764a6d1978dc61cb4499b15c45cb1b4 };
assign I9df5b63f66c162d517daa69f5d0e6095 = (I4c8d7e5474b19a7c63444d0cb6143728[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I42979deb711e94d6a366a9c125277bc7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00009_U (
.flogtanh_sel( Ia4bc4b7414bf31305ec8f63e7eda61e7[flogtanh_SEL-1:0]),
.flogtanh( I4fbe7db2d4288676183dc69ed56c9c68),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I12b0827207c31ed0661711adddb9b59f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4fbe7db2d4288676183dc69ed56c9c68 };
assign I1b40adfd6fa6c943dfa8d230d9e65514 = (Ia4bc4b7414bf31305ec8f63e7eda61e7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I12b0827207c31ed0661711adddb9b59f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00010_U (
.flogtanh_sel( Ibbebe287d56c7d627f3ffcf706575e77[flogtanh_SEL-1:0]),
.flogtanh( I99f0cc5986099cb57fbebf9e5e262c56),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If605c57ab8c22fa2cbb1e7f815274d80  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I99f0cc5986099cb57fbebf9e5e262c56 };
assign I0eb3df4d4094e09e6c4b3c788baed61f = (Ibbebe287d56c7d627f3ffcf706575e77[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If605c57ab8c22fa2cbb1e7f815274d80;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00011_U (
.flogtanh_sel( I83867e6ee369fff7e39ef5c8d5398fef[flogtanh_SEL-1:0]),
.flogtanh( I4f5bb7e206563a334d7e2dd100b37c35),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I82ed5aaddf52d30eba9c0116ef5e9a8c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4f5bb7e206563a334d7e2dd100b37c35 };
assign Id6f7923a16cc5adc96a730083153ca6d = (I83867e6ee369fff7e39ef5c8d5398fef[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I82ed5aaddf52d30eba9c0116ef5e9a8c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00012_U (
.flogtanh_sel( I1d40df7dbf99674f987bd06db714a702[flogtanh_SEL-1:0]),
.flogtanh( I59ecb14b5f34ebab3da4784709de66a4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I54e9afa2959a5a02f60ea11cfee788af  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I59ecb14b5f34ebab3da4784709de66a4 };
assign Idf8ebc0d747ae143aa61866e33d458c0 = (I1d40df7dbf99674f987bd06db714a702[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I54e9afa2959a5a02f60ea11cfee788af;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00013_U (
.flogtanh_sel( I92f42789cb81760ff2973e3a5fe915c3[flogtanh_SEL-1:0]),
.flogtanh( I54f5a8caf0e1c2df9477b37157d94995),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I31b86d750f70d42455bd426e8d3e494f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I54f5a8caf0e1c2df9477b37157d94995 };
assign Id682e531735437bc24abbf3d3d51e18b = (I92f42789cb81760ff2973e3a5fe915c3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I31b86d750f70d42455bd426e8d3e494f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00014_U (
.flogtanh_sel( Idbd5f2a25ab05808721cf9c403017565[flogtanh_SEL-1:0]),
.flogtanh( I77e1bed2da0ccf1475dcfe908d64f82c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic2923e2c0a77b23dbe0724bf452ea190  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I77e1bed2da0ccf1475dcfe908d64f82c };
assign I05ecce409cca00ea5b0df25de5a50cf2 = (Idbd5f2a25ab05808721cf9c403017565[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic2923e2c0a77b23dbe0724bf452ea190;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00046_00015_U (
.flogtanh_sel( I7ca5f07d6d3c2a045dfd55ae5214dd65[flogtanh_SEL-1:0]),
.flogtanh( I1a450ec193ccde2946f6ca20c0fa894c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie5fbbda327dbf0e90ad68ba42242fe21  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1a450ec193ccde2946f6ca20c0fa894c };
assign I831d214dcb4f8d534b5ddaaeaeeb81ce = (I7ca5f07d6d3c2a045dfd55ae5214dd65[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie5fbbda327dbf0e90ad68ba42242fe21;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00000_U (
.flogtanh_sel( I7f4e1445c68abbadce23944b99d206f9[flogtanh_SEL-1:0]),
.flogtanh( I01fbfc3b5c14733738f93a3487e54f35),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I261e7001e9ca425607de438bef1f7f4d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I01fbfc3b5c14733738f93a3487e54f35 };
assign Ia540866403683bc30504bace19bdda7b = (I7f4e1445c68abbadce23944b99d206f9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I261e7001e9ca425607de438bef1f7f4d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00001_U (
.flogtanh_sel( Id9f28016678e5e2127d9f0aa93e0b534[flogtanh_SEL-1:0]),
.flogtanh( Icff5d12020f78478c77210d9c692dfbe),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I27aac717f95c8b5b7114810c77bb0761  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icff5d12020f78478c77210d9c692dfbe };
assign I05fb1982415bd3fa78dd9a00af7a3d4a = (Id9f28016678e5e2127d9f0aa93e0b534[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I27aac717f95c8b5b7114810c77bb0761;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00002_U (
.flogtanh_sel( I6b939c57a8b7c7c51ab43e1b1df12f6a[flogtanh_SEL-1:0]),
.flogtanh( I6eb28698ab4105a74c6510dbcfefbc3c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id3820975eb9b8205aed04d02e9c21afb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6eb28698ab4105a74c6510dbcfefbc3c };
assign I977864efb0d94149cce7dc4d165f11de = (I6b939c57a8b7c7c51ab43e1b1df12f6a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id3820975eb9b8205aed04d02e9c21afb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00003_U (
.flogtanh_sel( Ic5d0df586d56bf4cb322d4c3ad677385[flogtanh_SEL-1:0]),
.flogtanh( I7cc0f835ad7a18683e1fdb5bcbfb7f2f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifbd4c6cc29fdd08d49bd7fd9f68051b3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7cc0f835ad7a18683e1fdb5bcbfb7f2f };
assign I9362b615a612599239e3b752a9334e8c = (Ic5d0df586d56bf4cb322d4c3ad677385[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifbd4c6cc29fdd08d49bd7fd9f68051b3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00004_U (
.flogtanh_sel( I2e287724873cf6761799eaf464ed6302[flogtanh_SEL-1:0]),
.flogtanh( I9389a0dfe5a82a903c89e1a468f0ad57),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2e9993aa302580a47147469355f65dcf  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9389a0dfe5a82a903c89e1a468f0ad57 };
assign I5d4fb4b5a5ad3dc48beebfa0e0cebbed = (I2e287724873cf6761799eaf464ed6302[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2e9993aa302580a47147469355f65dcf;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00005_U (
.flogtanh_sel( Ia7a10cffe31a53aafa1104b97543280b[flogtanh_SEL-1:0]),
.flogtanh( Idc4ce4afd846e212526d21a5e0cd1c14),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I187d0d6496e96f11c9c2c241213d405e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idc4ce4afd846e212526d21a5e0cd1c14 };
assign Ifb9b29c43f435452cc761218c509f5df = (Ia7a10cffe31a53aafa1104b97543280b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I187d0d6496e96f11c9c2c241213d405e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00006_U (
.flogtanh_sel( Ieeb089c6a18791a2227c8571913d689a[flogtanh_SEL-1:0]),
.flogtanh( I38a0ba1e69b467d4aed306e76ec3bfdb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1fd12d5a4d0a5d8d08117f57f2f4880e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I38a0ba1e69b467d4aed306e76ec3bfdb };
assign If2143db72bf9a02b64eb45b3a4faa39d = (Ieeb089c6a18791a2227c8571913d689a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1fd12d5a4d0a5d8d08117f57f2f4880e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00007_U (
.flogtanh_sel( Ib29b00328971c3cd67209a5ea5b63b0a[flogtanh_SEL-1:0]),
.flogtanh( I66279b0fa707a272f43ee929cb297945),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iba9bee3dd12c2559872c8498e4cd6f2b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I66279b0fa707a272f43ee929cb297945 };
assign Ice780b1695a8e80607a03dee3c426ffe = (Ib29b00328971c3cd67209a5ea5b63b0a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iba9bee3dd12c2559872c8498e4cd6f2b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00008_U (
.flogtanh_sel( I517e0868f2bb9a22c287a1f3eeaad2f3[flogtanh_SEL-1:0]),
.flogtanh( Ib091954846c14743e01fd4e7bafda1b5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8fecfe7601fa0d166db2b2fc9746129e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib091954846c14743e01fd4e7bafda1b5 };
assign I90b0296f5ef87dfaa6110fc2e9d6ed9d = (I517e0868f2bb9a22c287a1f3eeaad2f3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8fecfe7601fa0d166db2b2fc9746129e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00009_U (
.flogtanh_sel( I2bc9f76469e2a3f9846560ad1975cf54[flogtanh_SEL-1:0]),
.flogtanh( I3b8663f2adecb8da2c84dbb37341e25f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic3d6ada81005c125c29d8ff0abe88185  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3b8663f2adecb8da2c84dbb37341e25f };
assign Icd37da8ea84a606529e32b2db4eb7f5f = (I2bc9f76469e2a3f9846560ad1975cf54[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic3d6ada81005c125c29d8ff0abe88185;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00010_U (
.flogtanh_sel( I9f089315e435cd69d2929fdd936a8a77[flogtanh_SEL-1:0]),
.flogtanh( I19bc03089c6c288e1778bd1f197a3ce3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iddb333f6cb7253e92ba9e485a95c59c1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I19bc03089c6c288e1778bd1f197a3ce3 };
assign Ie626a24e3680f7d3995dd0c2ce60cbcc = (I9f089315e435cd69d2929fdd936a8a77[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iddb333f6cb7253e92ba9e485a95c59c1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00011_U (
.flogtanh_sel( I9b54c9fb4179423c731217286e329930[flogtanh_SEL-1:0]),
.flogtanh( I0988382a446b21da209d49d0d00bd6df),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I64f8fb4dc07decbd4e91436847143c23  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0988382a446b21da209d49d0d00bd6df };
assign Iebee55168fb47664095b11c9f6641124 = (I9b54c9fb4179423c731217286e329930[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I64f8fb4dc07decbd4e91436847143c23;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00012_U (
.flogtanh_sel( I82fb41ab743146badfd2e82258afb310[flogtanh_SEL-1:0]),
.flogtanh( I19f5cb50b27b6c5e40012df9397aa288),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I65c608dc3e2923360416cb08cfba6aeb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I19f5cb50b27b6c5e40012df9397aa288 };
assign Ic0954671eb1dc893c3932e456800fadf = (I82fb41ab743146badfd2e82258afb310[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I65c608dc3e2923360416cb08cfba6aeb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00013_U (
.flogtanh_sel( I5619b91de99eead78befdcba1c62411e[flogtanh_SEL-1:0]),
.flogtanh( I706ca74386e5778b30eca35432429bc3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I70bae72ccecf63dd5a367bf40b4ac870  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I706ca74386e5778b30eca35432429bc3 };
assign Ia4131464996aabab8aae1db85f6a50e4 = (I5619b91de99eead78befdcba1c62411e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I70bae72ccecf63dd5a367bf40b4ac870;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00014_U (
.flogtanh_sel( I83dd2047dece99cd841b2e7955819d57[flogtanh_SEL-1:0]),
.flogtanh( If6af0cc7a120b2897c3a69d54a554e86),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I32e73ad10e9df77b20d3eda78deeafac  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If6af0cc7a120b2897c3a69d54a554e86 };
assign I2de1ca2c390bdd3011fff4a359bb5332 = (I83dd2047dece99cd841b2e7955819d57[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I32e73ad10e9df77b20d3eda78deeafac;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00047_00015_U (
.flogtanh_sel( I8c927e66ccbf4d19f07af5ef9fbfe3fb[flogtanh_SEL-1:0]),
.flogtanh( I88ebe846173f486b07d2051a80bd055f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4688025bd745934e70eaa03f3bb7d089  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I88ebe846173f486b07d2051a80bd055f };
assign I6fb55222b69475b7168874423226ec9c = (I8c927e66ccbf4d19f07af5ef9fbfe3fb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4688025bd745934e70eaa03f3bb7d089;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00048_00000_U (
.flogtanh_sel( I0793fa8938acdf65486e5582d01b9e5a[flogtanh_SEL-1:0]),
.flogtanh( I2c577b130db6f4673704c858d454f3ea),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2c6ba69dd7827396366ce8e6513f8d4c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2c577b130db6f4673704c858d454f3ea };
assign I9b09b800a9dcd8ac36f25cb0324e748d = (I0793fa8938acdf65486e5582d01b9e5a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2c6ba69dd7827396366ce8e6513f8d4c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00048_00001_U (
.flogtanh_sel( Ied68d7ba0ee9974eb33767e737760b4d[flogtanh_SEL-1:0]),
.flogtanh( I383f23d4e769bbdc1c8acd9c660a0b3e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iecde1ff7e98a3f2aa847d1e55403f00f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I383f23d4e769bbdc1c8acd9c660a0b3e };
assign I74ac0327175f50f508a5013df298df02 = (Ied68d7ba0ee9974eb33767e737760b4d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iecde1ff7e98a3f2aa847d1e55403f00f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00048_00002_U (
.flogtanh_sel( I95ba37056659b29fd4318a68d85445e8[flogtanh_SEL-1:0]),
.flogtanh( Iea20a6ecf4bbf907d1a102bde797284f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I28ae9c81892f556ffbc3ed65b7ec0fb5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iea20a6ecf4bbf907d1a102bde797284f };
assign Ica26f542586d50c56ce0f3c00f36b388 = (I95ba37056659b29fd4318a68d85445e8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I28ae9c81892f556ffbc3ed65b7ec0fb5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00048_00003_U (
.flogtanh_sel( I08d7051a18f358d08728f1c401c15c47[flogtanh_SEL-1:0]),
.flogtanh( I77d655383c0c22b1af75d9308fab2e4f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1bfb39b04609b92c72d95b724eb3cae0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I77d655383c0c22b1af75d9308fab2e4f };
assign I7c6862830daffc98cb2c1fc121d82c38 = (I08d7051a18f358d08728f1c401c15c47[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1bfb39b04609b92c72d95b724eb3cae0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00048_00004_U (
.flogtanh_sel( I768b6f55827ac49eb6ac2655e9397be1[flogtanh_SEL-1:0]),
.flogtanh( I4a4ebb2f3389d67c4b7671e12fc5cd92),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I73ba173234b8583fa63ea947b5d2f957  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4a4ebb2f3389d67c4b7671e12fc5cd92 };
assign Icf19dd665616a8c96146b3ab9f46c741 = (I768b6f55827ac49eb6ac2655e9397be1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I73ba173234b8583fa63ea947b5d2f957;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00048_00005_U (
.flogtanh_sel( Ic66f737fe60c55d4c10e5d72b307a061[flogtanh_SEL-1:0]),
.flogtanh( Ibc927d678e218397e23147b5c0654fd9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9f0cce614937f873f39006b334729d72  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibc927d678e218397e23147b5c0654fd9 };
assign I97f2813ec39bbf1513faf66b3e38838a = (Ic66f737fe60c55d4c10e5d72b307a061[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9f0cce614937f873f39006b334729d72;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00048_00006_U (
.flogtanh_sel( I5653779f15c6c9b0f3b26927c48d6234[flogtanh_SEL-1:0]),
.flogtanh( Ib0358b6f47edcd54971935de215203f8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I129867553993fbc89983071472910fa4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib0358b6f47edcd54971935de215203f8 };
assign I716ee53e79883f69aa045380a357e913 = (I5653779f15c6c9b0f3b26927c48d6234[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I129867553993fbc89983071472910fa4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00048_00007_U (
.flogtanh_sel( Iac550729fc437fd67151fab57134ec88[flogtanh_SEL-1:0]),
.flogtanh( Iaa6f2bbd8a343ebf878da57badb4572b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2d6c9368bf6cc6e58ea202397528a736  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iaa6f2bbd8a343ebf878da57badb4572b };
assign I25c324feaca84e80f58075597e8c448f = (Iac550729fc437fd67151fab57134ec88[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2d6c9368bf6cc6e58ea202397528a736;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00048_00008_U (
.flogtanh_sel( I853b03c5826eedc3c67a2fae7a640212[flogtanh_SEL-1:0]),
.flogtanh( I823f1a0d2d757d5ca83dc7b5ca08e0f8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I715eedae273662cb8417d53b77f280c2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I823f1a0d2d757d5ca83dc7b5ca08e0f8 };
assign I7fc190647082a3d71614f46f670167bc = (I853b03c5826eedc3c67a2fae7a640212[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I715eedae273662cb8417d53b77f280c2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00049_00000_U (
.flogtanh_sel( If46a6b47c1c52243cc0bc92d1edb594f[flogtanh_SEL-1:0]),
.flogtanh( I1a650234a61a3ff90ea079e29d322069),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iab6f27ce8700543dfb7a8005ae320445  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1a650234a61a3ff90ea079e29d322069 };
assign Iebdf938a28594624f4d4a337356485cb = (If46a6b47c1c52243cc0bc92d1edb594f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iab6f27ce8700543dfb7a8005ae320445;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00049_00001_U (
.flogtanh_sel( I75b36a9b429cd657afc8151b9613aca6[flogtanh_SEL-1:0]),
.flogtanh( I70a7b1083c9593840759854430ee9d62),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaf6ebea4db33923d6db2c721d1dcd0d4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I70a7b1083c9593840759854430ee9d62 };
assign I3fd068d55154441ffd005999ea823fd0 = (I75b36a9b429cd657afc8151b9613aca6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaf6ebea4db33923d6db2c721d1dcd0d4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00049_00002_U (
.flogtanh_sel( Ife682dd9f677da4d27294fb61b141948[flogtanh_SEL-1:0]),
.flogtanh( I99aa55a3e285e62e9a8b50174e84b68c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic17b627fb3201547b05b457648431ad5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I99aa55a3e285e62e9a8b50174e84b68c };
assign Ic5ca74b66763c6e5591c7c2bfeeb0663 = (Ife682dd9f677da4d27294fb61b141948[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic17b627fb3201547b05b457648431ad5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00049_00003_U (
.flogtanh_sel( Ic2b6177a9c586b274b68b25584e6df2c[flogtanh_SEL-1:0]),
.flogtanh( Ief099d2084b84e0e23599d98102a13b7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iee1fb0a6e0aceddc45640b7ea4b4d0cd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ief099d2084b84e0e23599d98102a13b7 };
assign I5ab556386d2973354a5551ba9823e4ba = (Ic2b6177a9c586b274b68b25584e6df2c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iee1fb0a6e0aceddc45640b7ea4b4d0cd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00049_00004_U (
.flogtanh_sel( I0d23011c4381496a19cced7bf7960546[flogtanh_SEL-1:0]),
.flogtanh( I84aa89bab681c2fc7a8c7c6b47200dec),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I851d25c73aa5ee6bb26c0435353af3b8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I84aa89bab681c2fc7a8c7c6b47200dec };
assign I64f65df774d29696425ba460dda09b68 = (I0d23011c4381496a19cced7bf7960546[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I851d25c73aa5ee6bb26c0435353af3b8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00049_00005_U (
.flogtanh_sel( Ic5992d5eaeafd5dded641a7d9801e763[flogtanh_SEL-1:0]),
.flogtanh( I101b9397639b59fd53a88d17425e0c96),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I35e97af89c2791175cc545646eb7ba92  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I101b9397639b59fd53a88d17425e0c96 };
assign I9e09c25be9f877c1e1aaf79bf12c7943 = (Ic5992d5eaeafd5dded641a7d9801e763[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I35e97af89c2791175cc545646eb7ba92;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00049_00006_U (
.flogtanh_sel( Ic9e7fe68b9045c6c9eb86185b5f5872e[flogtanh_SEL-1:0]),
.flogtanh( Ic302f050dba883d8f4bd20b1030ba14d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I99b5120e2171e49d3320913b9e372936  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic302f050dba883d8f4bd20b1030ba14d };
assign I42c1d469ff97913cbf15e3ebee6fdfa8 = (Ic9e7fe68b9045c6c9eb86185b5f5872e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I99b5120e2171e49d3320913b9e372936;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00049_00007_U (
.flogtanh_sel( I51ad746720b5e6e09ab50f0283552f1a[flogtanh_SEL-1:0]),
.flogtanh( I848425f041888d7433b68900f259732a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idb7353d31a0038c904c4e25c78be46a5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I848425f041888d7433b68900f259732a };
assign If9f2a53dbf6e9b9a335a7657b7a2b468 = (I51ad746720b5e6e09ab50f0283552f1a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idb7353d31a0038c904c4e25c78be46a5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00049_00008_U (
.flogtanh_sel( I0c8964888a1315507f5d71959dd24cf0[flogtanh_SEL-1:0]),
.flogtanh( I2b4671193178503f5329954e74a399b3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I17ae1aa33db4ca2948befb43f1bd3d06  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2b4671193178503f5329954e74a399b3 };
assign I495f8be463b15db906474c518e0741e2 = (I0c8964888a1315507f5d71959dd24cf0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I17ae1aa33db4ca2948befb43f1bd3d06;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00050_00000_U (
.flogtanh_sel( Id4d4f814a0bb3418cbf70c306acf048f[flogtanh_SEL-1:0]),
.flogtanh( I97b93c6d963d51a819b1dc9ab3bf28ea),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ida342ed2e96314bb7c0182b3d895b647  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I97b93c6d963d51a819b1dc9ab3bf28ea };
assign I3e265a7dcf29687248b9275df49771fb = (Id4d4f814a0bb3418cbf70c306acf048f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ida342ed2e96314bb7c0182b3d895b647;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00050_00001_U (
.flogtanh_sel( Ic91bd7b4bd148e526ca21d4a5ba87be9[flogtanh_SEL-1:0]),
.flogtanh( I2593b1b30f4c97845a1f77c3f558b263),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If1d8968112c433d9d9bb309cc916fec9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2593b1b30f4c97845a1f77c3f558b263 };
assign Iffd94cf3a8a4681ff3327c90bf89bd8b = (Ic91bd7b4bd148e526ca21d4a5ba87be9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If1d8968112c433d9d9bb309cc916fec9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00050_00002_U (
.flogtanh_sel( I7959dddc32f0f181b3ba39149afe1016[flogtanh_SEL-1:0]),
.flogtanh( I3a4695c79b62f6baa47cdc939c4e2974),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6a927fb5af8b12fcd5d5b1b2b4e1f4b5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3a4695c79b62f6baa47cdc939c4e2974 };
assign Iea71417e738c6ca54c50aa014cc38627 = (I7959dddc32f0f181b3ba39149afe1016[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6a927fb5af8b12fcd5d5b1b2b4e1f4b5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00050_00003_U (
.flogtanh_sel( I087263600b5f38be072a4f1db787aea7[flogtanh_SEL-1:0]),
.flogtanh( Ibc577b2948aec87c0696c860d7efa1d7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic6b949621a3f4c61ac219919731f8f83  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibc577b2948aec87c0696c860d7efa1d7 };
assign Ic8df04756f67e6dd29f3374c5f86d451 = (I087263600b5f38be072a4f1db787aea7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic6b949621a3f4c61ac219919731f8f83;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00050_00004_U (
.flogtanh_sel( I78d17a56de5cbe08191ef23b9731c485[flogtanh_SEL-1:0]),
.flogtanh( I08401e4e9a1766a0034f45933b5bb29a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie8bfce645fef58bf090818dce30d86e4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I08401e4e9a1766a0034f45933b5bb29a };
assign I546122346a22ad64a6ab2b4978cde095 = (I78d17a56de5cbe08191ef23b9731c485[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie8bfce645fef58bf090818dce30d86e4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00050_00005_U (
.flogtanh_sel( I82f713a43596df3b935d6da6f8041dc2[flogtanh_SEL-1:0]),
.flogtanh( I5e5bb0de4fe6682a6beaa86f6cd1ca32),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ide2a4d41e8d2871f7c52249a8cb48ac1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5e5bb0de4fe6682a6beaa86f6cd1ca32 };
assign Icaae0fb0f460f68d690ab00697355a49 = (I82f713a43596df3b935d6da6f8041dc2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ide2a4d41e8d2871f7c52249a8cb48ac1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00050_00006_U (
.flogtanh_sel( I422987396853a6a39dabb6e7ddbf91fb[flogtanh_SEL-1:0]),
.flogtanh( Ia487e80f0010e7cb34aa12471e62a62f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib58e63392e279cbb87c4e5be4e4b0109  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia487e80f0010e7cb34aa12471e62a62f };
assign I42455e7e4d0c63f97702d204d18a446e = (I422987396853a6a39dabb6e7ddbf91fb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib58e63392e279cbb87c4e5be4e4b0109;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00050_00007_U (
.flogtanh_sel( Ibb6556671e104141dd33188ea5fc024d[flogtanh_SEL-1:0]),
.flogtanh( I3bee9305e2f4456aae800bbb174b7843),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic680a004d350df1379eddb3ed06be34e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3bee9305e2f4456aae800bbb174b7843 };
assign Iaec2f15665e83416bc140890f3cdde9a = (Ibb6556671e104141dd33188ea5fc024d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic680a004d350df1379eddb3ed06be34e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00050_00008_U (
.flogtanh_sel( Ie42ce76076a2a5e887e0112086012da6[flogtanh_SEL-1:0]),
.flogtanh( I14f1aa0dbf6f1f0fbf6b5f996e229a04),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8074f2ecf0e4178d0b8d58f4d6680282  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I14f1aa0dbf6f1f0fbf6b5f996e229a04 };
assign I487391402b6aa27bf212724a37ea9c33 = (Ie42ce76076a2a5e887e0112086012da6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8074f2ecf0e4178d0b8d58f4d6680282;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00051_00000_U (
.flogtanh_sel( I4aea430599b9c0702b3bebd5960b5c91[flogtanh_SEL-1:0]),
.flogtanh( If87afc1cf342dca9986f798c38a69dab),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I20b0882e61c68796b057b0a9d237a979  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If87afc1cf342dca9986f798c38a69dab };
assign Ia9f375709014a9d553d46cff2799b59f = (I4aea430599b9c0702b3bebd5960b5c91[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I20b0882e61c68796b057b0a9d237a979;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00051_00001_U (
.flogtanh_sel( Icbe11a3970136e485eee1bc5053e7273[flogtanh_SEL-1:0]),
.flogtanh( Ibb1c020ea255a966e54c00fc7cc745b5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4c1ecb851699ea3c2642c78fa44b04e6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibb1c020ea255a966e54c00fc7cc745b5 };
assign I34d428a56bd0142a9be9f627f1c3c87f = (Icbe11a3970136e485eee1bc5053e7273[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4c1ecb851699ea3c2642c78fa44b04e6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00051_00002_U (
.flogtanh_sel( I0a7f1ea1719c1f5ff104445a4130a5a8[flogtanh_SEL-1:0]),
.flogtanh( Icae8a2980dd7403caf72820ae508885b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I421cb46488584e6314f701cfe34d3e79  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icae8a2980dd7403caf72820ae508885b };
assign I57db98eb439d59a895dabe029c6a3a8b = (I0a7f1ea1719c1f5ff104445a4130a5a8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I421cb46488584e6314f701cfe34d3e79;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00051_00003_U (
.flogtanh_sel( I1802d759f26dd919bc315bfd4156238d[flogtanh_SEL-1:0]),
.flogtanh( Ic8f858d7f7a16b771933741d31679dc1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibed20c973d23c4058efffc1575d66478  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic8f858d7f7a16b771933741d31679dc1 };
assign I9937af6fcf9d834f308bc3683d524981 = (I1802d759f26dd919bc315bfd4156238d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibed20c973d23c4058efffc1575d66478;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00051_00004_U (
.flogtanh_sel( I2148493e253783fad70f4f2807b83008[flogtanh_SEL-1:0]),
.flogtanh( I9dcf19da38f352fe7fa27c22bff08c19),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2f5e17be80bab46917da109cf7ac3532  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9dcf19da38f352fe7fa27c22bff08c19 };
assign I463f4f370e1ecad71de44780eff10df4 = (I2148493e253783fad70f4f2807b83008[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2f5e17be80bab46917da109cf7ac3532;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00051_00005_U (
.flogtanh_sel( I39e7f78d33aa7f50264908d2efe23634[flogtanh_SEL-1:0]),
.flogtanh( I2bc787aa749db4a5f48bd917715a11d5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I43b6cac96c5c2236629f6ee87f13e0be  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2bc787aa749db4a5f48bd917715a11d5 };
assign I53309409a6059c3bd39f037c23ec3458 = (I39e7f78d33aa7f50264908d2efe23634[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I43b6cac96c5c2236629f6ee87f13e0be;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00051_00006_U (
.flogtanh_sel( I844be5874def16af98de935019f35fe8[flogtanh_SEL-1:0]),
.flogtanh( I3d072e173fd12ac9d802a29a0ff4378c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I54a8f8a82aa219427914ca74da599696  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3d072e173fd12ac9d802a29a0ff4378c };
assign I2603e0b8b93f6680e44c9c8883f6512c = (I844be5874def16af98de935019f35fe8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I54a8f8a82aa219427914ca74da599696;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00051_00007_U (
.flogtanh_sel( Iee5172ba70a6e368b4903f9ff1d93471[flogtanh_SEL-1:0]),
.flogtanh( I2115d62275a57ec7273e3631c0a32872),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I23e89a266dd6a09d486b129eea48fae5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2115d62275a57ec7273e3631c0a32872 };
assign Iab354cc9ac1173335c0efeef694f3567 = (Iee5172ba70a6e368b4903f9ff1d93471[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I23e89a266dd6a09d486b129eea48fae5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00051_00008_U (
.flogtanh_sel( I1f34b473283291e0970879465c005e2f[flogtanh_SEL-1:0]),
.flogtanh( I91bc663fcd7f86a066b8b3f93b1dcfc2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8b68b47c8e9b4055b176745aec55b3b2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I91bc663fcd7f86a066b8b3f93b1dcfc2 };
assign I6c19936ca2edeb0e261e880a1055e964 = (I1f34b473283291e0970879465c005e2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8b68b47c8e9b4055b176745aec55b3b2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00000_U (
.flogtanh_sel( Ie1e0b5120737a7f4bf845618ccd22239[flogtanh_SEL-1:0]),
.flogtanh( I988c0d94f97329dd1cff7d913cb449e7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1195ee9289f2afca25519bb6d493e73a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I988c0d94f97329dd1cff7d913cb449e7 };
assign Ifebfa58419ecd22a334ed4b67f5c3581 = (Ie1e0b5120737a7f4bf845618ccd22239[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1195ee9289f2afca25519bb6d493e73a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00001_U (
.flogtanh_sel( I8abec3020ee5358f8768e5595e9992b4[flogtanh_SEL-1:0]),
.flogtanh( If444a37a85774dcc2769ffd74b785e46),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2844ec353c6ac19013e7a64d350f0204  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If444a37a85774dcc2769ffd74b785e46 };
assign I71a28e8525f07dabeabe4b4f45f353d0 = (I8abec3020ee5358f8768e5595e9992b4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2844ec353c6ac19013e7a64d350f0204;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00002_U (
.flogtanh_sel( I6fe683073211a484cb6e3c416b365d9f[flogtanh_SEL-1:0]),
.flogtanh( Idbb89639b8399b57b190efd898643328),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie4848a127b84c06712bd2b40d80b214d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idbb89639b8399b57b190efd898643328 };
assign I514830acdad20c4ff3d078477e939b4b = (I6fe683073211a484cb6e3c416b365d9f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie4848a127b84c06712bd2b40d80b214d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00003_U (
.flogtanh_sel( Id7d764da58ade36853e8a45b5ee19dc3[flogtanh_SEL-1:0]),
.flogtanh( Ib1d70f302858eb7c78fb834071616a9b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id93016d32ebfabc6e464df96ae3aa74c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib1d70f302858eb7c78fb834071616a9b };
assign I036342f6be0f2e2f1f4927099a5c4a78 = (Id7d764da58ade36853e8a45b5ee19dc3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id93016d32ebfabc6e464df96ae3aa74c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00004_U (
.flogtanh_sel( I3cee2fdf353643deac7d6bca20c8fb52[flogtanh_SEL-1:0]),
.flogtanh( I82bd4ea32da7ae3a0d5938fc8a1424c5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0ed0efac703623c9a35ffb79a57683dc  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I82bd4ea32da7ae3a0d5938fc8a1424c5 };
assign Iedb655aa25e5f0e35137ec6c3acdc527 = (I3cee2fdf353643deac7d6bca20c8fb52[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0ed0efac703623c9a35ffb79a57683dc;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00005_U (
.flogtanh_sel( Ie9b8f8f0434fe3783c3d8f68fef30e50[flogtanh_SEL-1:0]),
.flogtanh( I6964f2e681e9cdf63fbc0358cb6edcca),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2f1a1b3caf70a00d30678c22f68f9cfe  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6964f2e681e9cdf63fbc0358cb6edcca };
assign I0c59e8c82a31aacbf5977ff778a7ff49 = (Ie9b8f8f0434fe3783c3d8f68fef30e50[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2f1a1b3caf70a00d30678c22f68f9cfe;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00006_U (
.flogtanh_sel( I68cba8ad7742cbb34d0b1fb16be4a58a[flogtanh_SEL-1:0]),
.flogtanh( I41aeb75239ce0d636288e8ceb0665b34),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8acdcab405f76f4bf751e8860a50e614  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I41aeb75239ce0d636288e8ceb0665b34 };
assign I1b6d20c64b9f23fb6c30f723546aa285 = (I68cba8ad7742cbb34d0b1fb16be4a58a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8acdcab405f76f4bf751e8860a50e614;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00007_U (
.flogtanh_sel( Idcea56657d40e0fdf9a1c2d920938fd6[flogtanh_SEL-1:0]),
.flogtanh( Ie0d3fd5e7c38c10fdcae3f1b217c28f4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I88ede5095d3876c7ca6dac02faa3eede  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie0d3fd5e7c38c10fdcae3f1b217c28f4 };
assign I0d66aa55747362354aa81d96057bc4c2 = (Idcea56657d40e0fdf9a1c2d920938fd6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I88ede5095d3876c7ca6dac02faa3eede;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00008_U (
.flogtanh_sel( Ic549ffab8f0ce161a177faa2ffd1326d[flogtanh_SEL-1:0]),
.flogtanh( Ia8b7d74eaf227e697c3eb58b31eb355f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I68bc064fabdc9564021be1d29f3cbb7a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia8b7d74eaf227e697c3eb58b31eb355f };
assign I1ea33707e40a2e41513fdb3118371437 = (Ic549ffab8f0ce161a177faa2ffd1326d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I68bc064fabdc9564021be1d29f3cbb7a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00009_U (
.flogtanh_sel( I4d463d500f93f74b2724972ec1d62439[flogtanh_SEL-1:0]),
.flogtanh( I79034cd4180d03348de2c101927048a7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idfd56dd8b81f3ec49acfa9131d4b78c4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I79034cd4180d03348de2c101927048a7 };
assign I68c85727adecde0aa8aa66ed08c4b502 = (I4d463d500f93f74b2724972ec1d62439[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idfd56dd8b81f3ec49acfa9131d4b78c4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00010_U (
.flogtanh_sel( Iba2f362e263953331649c726afa9c481[flogtanh_SEL-1:0]),
.flogtanh( Id23895e0696cdd27e3087294fb52a65b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I777937fc3cbdcb60a10ee0c0d1f56dc5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id23895e0696cdd27e3087294fb52a65b };
assign Iebd050e29044153d5881ef80b2db8c28 = (Iba2f362e263953331649c726afa9c481[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I777937fc3cbdcb60a10ee0c0d1f56dc5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00052_00011_U (
.flogtanh_sel( I6a053d931fb030e03d4882856d3bda75[flogtanh_SEL-1:0]),
.flogtanh( I43939a168f9f5e476262ace39c6ae483),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2de42de0be5ebc2ee41fb217953cb823  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I43939a168f9f5e476262ace39c6ae483 };
assign I3c057d64cf4fca0238a874f0ced99c76 = (I6a053d931fb030e03d4882856d3bda75[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2de42de0be5ebc2ee41fb217953cb823;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00000_U (
.flogtanh_sel( I27ede93004e0c240efaa56cc8c570910[flogtanh_SEL-1:0]),
.flogtanh( Ie5167faac3e6510d4b208a1bdc0cd44c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ied21906ec121c7c7da1d0268e93ab0a6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie5167faac3e6510d4b208a1bdc0cd44c };
assign I066cd52173ec5dbce9a3f470d73325af = (I27ede93004e0c240efaa56cc8c570910[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ied21906ec121c7c7da1d0268e93ab0a6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00001_U (
.flogtanh_sel( I61a11c1711ca10eefea3438722b40bff[flogtanh_SEL-1:0]),
.flogtanh( I1cad8b885a541dd049093ce60c3f8a06),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I074d42d6f79dd8786745ad7b0f59b3e5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1cad8b885a541dd049093ce60c3f8a06 };
assign Ic7ad59f6a232a997706d17b4098e0324 = (I61a11c1711ca10eefea3438722b40bff[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I074d42d6f79dd8786745ad7b0f59b3e5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00002_U (
.flogtanh_sel( Ia7924c88692cfddf24fb1eff66eacb7e[flogtanh_SEL-1:0]),
.flogtanh( Icd2d69f12d4744ce7b09fce7f27ab830),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I78cfd6df12d7b773c498ed763953c8a2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icd2d69f12d4744ce7b09fce7f27ab830 };
assign Icf8cfc800f0a2aa5140a7f83f035b0cc = (Ia7924c88692cfddf24fb1eff66eacb7e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I78cfd6df12d7b773c498ed763953c8a2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00003_U (
.flogtanh_sel( Ibcfd01e622f7f5a5156dd9b335b4e5e0[flogtanh_SEL-1:0]),
.flogtanh( Ic9ee0243e36f66f462eb3d4ce93fdde9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3e452666c55d9b30beef77c58690c8fd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic9ee0243e36f66f462eb3d4ce93fdde9 };
assign I6bfbf7ff79ff0a6facc9ba5031239644 = (Ibcfd01e622f7f5a5156dd9b335b4e5e0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3e452666c55d9b30beef77c58690c8fd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00004_U (
.flogtanh_sel( I7f6f418ea51b4298da8758bda3f6a21b[flogtanh_SEL-1:0]),
.flogtanh( I5353c3239ddb4d7fa7094e413b5303b1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5524ea6d4e43842521569ba37425b387  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5353c3239ddb4d7fa7094e413b5303b1 };
assign I78ade92efd265027807c861be44a10af = (I7f6f418ea51b4298da8758bda3f6a21b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5524ea6d4e43842521569ba37425b387;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00005_U (
.flogtanh_sel( I7185da8937449e23abdd0f39a4b3ed7d[flogtanh_SEL-1:0]),
.flogtanh( Idfca1b1d8041e5808799499e8c8dcf5e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8153350f4b99d2a42acc18f730911337  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idfca1b1d8041e5808799499e8c8dcf5e };
assign I2bc5a10c587d89d10021aa5eaafb490a = (I7185da8937449e23abdd0f39a4b3ed7d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8153350f4b99d2a42acc18f730911337;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00006_U (
.flogtanh_sel( Idc3e3ffa31d9b76c7cf9358a5b2e65d7[flogtanh_SEL-1:0]),
.flogtanh( I4710d61c763098027934286c6a9f3714),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I685829af9b536012f05d3a22e0d7651b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4710d61c763098027934286c6a9f3714 };
assign I30080cc6c03bbe933165d266558a822c = (Idc3e3ffa31d9b76c7cf9358a5b2e65d7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I685829af9b536012f05d3a22e0d7651b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00007_U (
.flogtanh_sel( I31fe8c887c4aff7c69336676cd31aaa1[flogtanh_SEL-1:0]),
.flogtanh( If6a04c29b7205c5db5f2ff3cf302c45f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibb607d3707048ec1dd1f126852667fcb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If6a04c29b7205c5db5f2ff3cf302c45f };
assign I7e28234bdf66ab5489d36d15678db797 = (I31fe8c887c4aff7c69336676cd31aaa1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibb607d3707048ec1dd1f126852667fcb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00008_U (
.flogtanh_sel( I59684d5fe6bbb4b54ac097bd25fceef5[flogtanh_SEL-1:0]),
.flogtanh( Ib5d9348a114627a8b1f56aca968d20b1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib948458593df6c9b4bef35c88845492d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib5d9348a114627a8b1f56aca968d20b1 };
assign I74b3c9dd3a8168aacd4369b9ff68fdfd = (I59684d5fe6bbb4b54ac097bd25fceef5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib948458593df6c9b4bef35c88845492d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00009_U (
.flogtanh_sel( I86a7cd69148f9590ce91d0aa270d6c54[flogtanh_SEL-1:0]),
.flogtanh( I4e2b59a03731959106d469ffee7b7d33),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifbebc06fa0ddc76aa8053ee669fda467  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4e2b59a03731959106d469ffee7b7d33 };
assign Ia7046faae1ab05978e4b32bd44049fb9 = (I86a7cd69148f9590ce91d0aa270d6c54[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifbebc06fa0ddc76aa8053ee669fda467;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00010_U (
.flogtanh_sel( Iabce1ccdd968980f622f0e137b159d11[flogtanh_SEL-1:0]),
.flogtanh( Ic6d519691c7543b1bd0707a8c9899088),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I059d9b49b8c6de67643992e5ef74d939  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic6d519691c7543b1bd0707a8c9899088 };
assign I0c5250aaca86185fed5978438c8861b6 = (Iabce1ccdd968980f622f0e137b159d11[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I059d9b49b8c6de67643992e5ef74d939;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00053_00011_U (
.flogtanh_sel( Iff02977d7b4c733cca1794246f630931[flogtanh_SEL-1:0]),
.flogtanh( Icc6bde490bd8df2ce5efe8cfb24cf5f5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I141b6f8e6baa353f2527dc1171c95908  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icc6bde490bd8df2ce5efe8cfb24cf5f5 };
assign Ic78949e07e643f571f23df7e8f15d9fb = (Iff02977d7b4c733cca1794246f630931[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I141b6f8e6baa353f2527dc1171c95908;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00000_U (
.flogtanh_sel( I9026c904e5ead7ff2994c4f781d61466[flogtanh_SEL-1:0]),
.flogtanh( I861bd8df5caf968dc6edd7a05d690033),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I891992837c6e3d393516506efec821e1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I861bd8df5caf968dc6edd7a05d690033 };
assign Ifb8b3586a5b69b20cf03eabf51344ab6 = (I9026c904e5ead7ff2994c4f781d61466[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I891992837c6e3d393516506efec821e1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00001_U (
.flogtanh_sel( I99d7489ba87c629c6dd9702a9bbfd3c8[flogtanh_SEL-1:0]),
.flogtanh( I6f44882493f9eadbdbe1ac46a3d2a43b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9739e5853bd26c50167491b69e92ed6f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6f44882493f9eadbdbe1ac46a3d2a43b };
assign I9ea09f27ce4484f2e7fc3a6b6d6ecb7c = (I99d7489ba87c629c6dd9702a9bbfd3c8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9739e5853bd26c50167491b69e92ed6f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00002_U (
.flogtanh_sel( Ifaf191e0d00ba6da7019c2efcf08e1d9[flogtanh_SEL-1:0]),
.flogtanh( I5a3ec39885fba8d015009d671a1cb544),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I80c41a49bba592ec70c6ca394bb48845  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5a3ec39885fba8d015009d671a1cb544 };
assign If0b9225e759438be175c4128c78605ea = (Ifaf191e0d00ba6da7019c2efcf08e1d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I80c41a49bba592ec70c6ca394bb48845;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00003_U (
.flogtanh_sel( I4c295991fb08c90862a2f3ba6489000a[flogtanh_SEL-1:0]),
.flogtanh( Ic4e6d76148a8170d1af0c95f370367a5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia96cc576fbc424161dcc350151e4476d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic4e6d76148a8170d1af0c95f370367a5 };
assign I33d941ad9d4858fcfb77f0f6cf99d2ec = (I4c295991fb08c90862a2f3ba6489000a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia96cc576fbc424161dcc350151e4476d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00004_U (
.flogtanh_sel( Iee61d179da125934298400256788cbb8[flogtanh_SEL-1:0]),
.flogtanh( I244bd772f9d750b4e1800e0b0ca67d63),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3abbd492752bc871096dac47e3208d01  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I244bd772f9d750b4e1800e0b0ca67d63 };
assign Ia0868eee7e7e0640ce1a4d3ca9c001cb = (Iee61d179da125934298400256788cbb8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3abbd492752bc871096dac47e3208d01;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00005_U (
.flogtanh_sel( If87c84440426fb24070372dc1d4bf315[flogtanh_SEL-1:0]),
.flogtanh( I00c203d60e09f1cccdadb8ebff2de650),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iff5e7ff31a18e5a3947f16c456cb4bf2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I00c203d60e09f1cccdadb8ebff2de650 };
assign Icb3ab2c67a87b2ee158e0021b72fc186 = (If87c84440426fb24070372dc1d4bf315[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iff5e7ff31a18e5a3947f16c456cb4bf2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00006_U (
.flogtanh_sel( Ib9259a807b31c1b7a528d336bfc403ee[flogtanh_SEL-1:0]),
.flogtanh( I20c7780e77b49d31808e59cae58968a9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6f437a921b54934b3a5d13eb2d8e4b5e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I20c7780e77b49d31808e59cae58968a9 };
assign I5b64997d083769666741c794dd92fb7f = (Ib9259a807b31c1b7a528d336bfc403ee[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6f437a921b54934b3a5d13eb2d8e4b5e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00007_U (
.flogtanh_sel( I411c4d909b2a571e685cd703245516d7[flogtanh_SEL-1:0]),
.flogtanh( Ia332fad029505e5975156f8e13910358),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieb8e5fdc6ac722d69775b46b0f081bf7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia332fad029505e5975156f8e13910358 };
assign I0a3323aac825506435068f6746aee974 = (I411c4d909b2a571e685cd703245516d7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieb8e5fdc6ac722d69775b46b0f081bf7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00008_U (
.flogtanh_sel( If8425453cca8fc8623cb85375c4b8a1d[flogtanh_SEL-1:0]),
.flogtanh( I9cc95185621ad5718a905092c03315f8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8b60818e4831ff872dd58accdbe94b30  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9cc95185621ad5718a905092c03315f8 };
assign Ibec442c099da091afcf75a7c970bf8ea = (If8425453cca8fc8623cb85375c4b8a1d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8b60818e4831ff872dd58accdbe94b30;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00009_U (
.flogtanh_sel( I654b497f62df75fa283127b5de29b1ad[flogtanh_SEL-1:0]),
.flogtanh( Iba2a341076f0506aeac3769e71b91f43),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9e1401baae9fab762f3ac1382b4658ed  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iba2a341076f0506aeac3769e71b91f43 };
assign If3a79ede332c39a8d2a276de833242f6 = (I654b497f62df75fa283127b5de29b1ad[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9e1401baae9fab762f3ac1382b4658ed;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00010_U (
.flogtanh_sel( I2768519342f7b8a1ee40c1d5ac502b66[flogtanh_SEL-1:0]),
.flogtanh( Ic9e82f153d0e690d5ea47ee159523b72),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I19e98430858ce2db7853b31e4a8409f0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic9e82f153d0e690d5ea47ee159523b72 };
assign I49ccb3e14fe61618806e791ecb4f4eae = (I2768519342f7b8a1ee40c1d5ac502b66[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I19e98430858ce2db7853b31e4a8409f0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00054_00011_U (
.flogtanh_sel( I8e354c1c5ba44fe5430887248ce0c43b[flogtanh_SEL-1:0]),
.flogtanh( Ia265b95249953a7867c611d475d01169),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I58ed96e69f7ce8d98d44b992f52fe7ca  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia265b95249953a7867c611d475d01169 };
assign I461ebbf3a02ae63e2eb27531b1370f24 = (I8e354c1c5ba44fe5430887248ce0c43b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I58ed96e69f7ce8d98d44b992f52fe7ca;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00000_U (
.flogtanh_sel( I8970d8a8aea29913e8696c14c153d16e[flogtanh_SEL-1:0]),
.flogtanh( I5ef2899606d7f08aa6d0028f9f113e38),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie2b3c1982842e9b4f2befd0fce03a1cf  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5ef2899606d7f08aa6d0028f9f113e38 };
assign Ice66c108aa66981051df71e226cb0e4d = (I8970d8a8aea29913e8696c14c153d16e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie2b3c1982842e9b4f2befd0fce03a1cf;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00001_U (
.flogtanh_sel( I3555c6e2fd480a6be11549bf95a9b0b1[flogtanh_SEL-1:0]),
.flogtanh( Idf3a6723fec1ef62c1e37a419590122c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1a66d7f556b0f90b7f7c1321d1998cc3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idf3a6723fec1ef62c1e37a419590122c };
assign I645ff0d8c0a87ba7f792fc83f342b958 = (I3555c6e2fd480a6be11549bf95a9b0b1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1a66d7f556b0f90b7f7c1321d1998cc3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00002_U (
.flogtanh_sel( I8d5600a352e8ba4756f917f912fda6dd[flogtanh_SEL-1:0]),
.flogtanh( I0bde2fc197586c74374ffb402956baf5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I87ace9b2a7e2e5ced87a85ad45c0b0c9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0bde2fc197586c74374ffb402956baf5 };
assign Ica94017f26e96fb22a47add326ee126e = (I8d5600a352e8ba4756f917f912fda6dd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I87ace9b2a7e2e5ced87a85ad45c0b0c9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00003_U (
.flogtanh_sel( I7e99d73c95e7ae5c3fe07a3c60ef52eb[flogtanh_SEL-1:0]),
.flogtanh( I9182b3349816b6ddaffde1cbec78339e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia51a22a9b78f5e3e8b6e86b919ceb13d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9182b3349816b6ddaffde1cbec78339e };
assign Id32e7ad5b1aa825732d9b26d0fa02ca1 = (I7e99d73c95e7ae5c3fe07a3c60ef52eb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia51a22a9b78f5e3e8b6e86b919ceb13d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00004_U (
.flogtanh_sel( I831633aebe5c6a52b98d630205376f3a[flogtanh_SEL-1:0]),
.flogtanh( I5bf9702e2afd6c791b28c76c84aeb886),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibb6b016405d27b6863c2d182e9465a5e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5bf9702e2afd6c791b28c76c84aeb886 };
assign I51b5e641856239367cf43f9b5679b268 = (I831633aebe5c6a52b98d630205376f3a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibb6b016405d27b6863c2d182e9465a5e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00005_U (
.flogtanh_sel( I82e35482de74223be0d2558334ac2dfb[flogtanh_SEL-1:0]),
.flogtanh( Ifbd7b868d9cb7e04bf2189922bcb9c92),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2bd977c2b670677802c6486507b0672f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifbd7b868d9cb7e04bf2189922bcb9c92 };
assign I2d1a5645b126761fc7fb70d24e37189a = (I82e35482de74223be0d2558334ac2dfb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2bd977c2b670677802c6486507b0672f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00006_U (
.flogtanh_sel( Iae2a6f9649ef1bb193e4f0ab5ecbc3e3[flogtanh_SEL-1:0]),
.flogtanh( Ib78e7602e521bc064d5cd9efe10ec6b1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie9cd522fdd4e6e94287e7a8ce329c31e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib78e7602e521bc064d5cd9efe10ec6b1 };
assign I49f5f87662fbb540d72c94bfd1acd060 = (Iae2a6f9649ef1bb193e4f0ab5ecbc3e3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie9cd522fdd4e6e94287e7a8ce329c31e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00007_U (
.flogtanh_sel( Ie8eca65d791ad2f6e8f4ed244f22ae3d[flogtanh_SEL-1:0]),
.flogtanh( I0497115b3dd67c6538039969368e03ae),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1330526fdd2ffaa0137d4735167961b5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0497115b3dd67c6538039969368e03ae };
assign I30253dc91301ca27b5732312c01145e0 = (Ie8eca65d791ad2f6e8f4ed244f22ae3d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1330526fdd2ffaa0137d4735167961b5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00008_U (
.flogtanh_sel( Ic24146b01094df9b9ccd455a791f239d[flogtanh_SEL-1:0]),
.flogtanh( Ieba8e28ee660b8e2d78909d61ced3233),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib9939f977a24ec96a60403bc4e8d4ef3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ieba8e28ee660b8e2d78909d61ced3233 };
assign I143f5e324716a94d24ada126886bf895 = (Ic24146b01094df9b9ccd455a791f239d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib9939f977a24ec96a60403bc4e8d4ef3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00009_U (
.flogtanh_sel( I1c9031fd54ff9417d44c9fb17dc1fc63[flogtanh_SEL-1:0]),
.flogtanh( I12e6fe32f6159ce6bb8be6411af2b7bb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6d268ba2240ef4c0ac98f5e771964820  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I12e6fe32f6159ce6bb8be6411af2b7bb };
assign If64aa8c220b9ab6652e081da7e404e80 = (I1c9031fd54ff9417d44c9fb17dc1fc63[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6d268ba2240ef4c0ac98f5e771964820;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00010_U (
.flogtanh_sel( Idefa20487bc5ba6daff03e6b327d76c6[flogtanh_SEL-1:0]),
.flogtanh( I03392e42f99b06cb65b38122c1e4dc81),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If6639d10ed80985c8e322a85cfe65887  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I03392e42f99b06cb65b38122c1e4dc81 };
assign I1092325b801600fa7ec85fa640167da9 = (Idefa20487bc5ba6daff03e6b327d76c6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If6639d10ed80985c8e322a85cfe65887;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00055_00011_U (
.flogtanh_sel( I6f984fd9ea27b40ab3afeac8afd29ade[flogtanh_SEL-1:0]),
.flogtanh( I32270eb6cf0594020ee19abb2edfe93d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5d4d3b9363d24d988468d1782347a41c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I32270eb6cf0594020ee19abb2edfe93d };
assign Ib028686da9c849e827cf249a744b7db3 = (I6f984fd9ea27b40ab3afeac8afd29ade[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5d4d3b9363d24d988468d1782347a41c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00056_00000_U (
.flogtanh_sel( I0be92debced4961df5f461fe81e80bf1[flogtanh_SEL-1:0]),
.flogtanh( Ib135d3d7d338f5ff3a1f504aec754bbd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6461781f905b7694ad26c54d6f8cb062  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib135d3d7d338f5ff3a1f504aec754bbd };
assign I5f3ff7fa8686f7a380302d71b88cfb4b = (I0be92debced4961df5f461fe81e80bf1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6461781f905b7694ad26c54d6f8cb062;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00057_00000_U (
.flogtanh_sel( Ia7bdaba4c6601b7146498aea6c9a3e07[flogtanh_SEL-1:0]),
.flogtanh( Id9cbc2e4b0f437840f028c7273d49416),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I731ddcd050cee04fdfd5724c7236e9fb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id9cbc2e4b0f437840f028c7273d49416 };
assign Ic01904f7c518990eff2dc1de127676c4 = (Ia7bdaba4c6601b7146498aea6c9a3e07[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I731ddcd050cee04fdfd5724c7236e9fb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00058_00000_U (
.flogtanh_sel( Id450c0a1cabe087be051fbf4158e6016[flogtanh_SEL-1:0]),
.flogtanh( I98b5a84c247422b51abf63a705fbb5f7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0306fc584747e83ab0f2be50b228a1ad  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I98b5a84c247422b51abf63a705fbb5f7 };
assign I43f2ddd9780f86af489f8deae51168ec = (Id450c0a1cabe087be051fbf4158e6016[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0306fc584747e83ab0f2be50b228a1ad;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00059_00000_U (
.flogtanh_sel( I656d0d69f6e243746b87ad67764dbc3d[flogtanh_SEL-1:0]),
.flogtanh( I0ae39e89061b4f8c5c0e56eba2f48889),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7b2920a709b708955c261faa5ffda88c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0ae39e89061b4f8c5c0e56eba2f48889 };
assign I0a013fff6c792363bd7feb03d9691db8 = (I656d0d69f6e243746b87ad67764dbc3d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7b2920a709b708955c261faa5ffda88c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00060_00000_U (
.flogtanh_sel( Iab9d870dc1ad159bbaecb20a9b72f005[flogtanh_SEL-1:0]),
.flogtanh( If612cf94a3cefcfb844d6e975ba4aada),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iae6e4e88f9136c6c09f4fe0c9825e2e0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If612cf94a3cefcfb844d6e975ba4aada };
assign I7cf8401bf6893eab0b9f33a0f91ddd05 = (Iab9d870dc1ad159bbaecb20a9b72f005[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iae6e4e88f9136c6c09f4fe0c9825e2e0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00061_00000_U (
.flogtanh_sel( Id53b60854f19e095c38f2c255dc57f29[flogtanh_SEL-1:0]),
.flogtanh( I3dab04eb1045e1b3b6bb47e0f4c390ad),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic729485a48ee429c62eab4aef90b03b8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3dab04eb1045e1b3b6bb47e0f4c390ad };
assign Ic7ccbeaf4ab94d0660eb7a0533723e24 = (Id53b60854f19e095c38f2c255dc57f29[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic729485a48ee429c62eab4aef90b03b8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00062_00000_U (
.flogtanh_sel( If9ba44a2e4a8f0b61692fc69ebeb82bd[flogtanh_SEL-1:0]),
.flogtanh( I447db5cb14c9588418037bbb793a6274),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I009290dfe067ac2cc190b53a07374b34  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I447db5cb14c9588418037bbb793a6274 };
assign I08043393cb7f2558c145a698ea6652c9 = (If9ba44a2e4a8f0b61692fc69ebeb82bd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I009290dfe067ac2cc190b53a07374b34;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00063_00000_U (
.flogtanh_sel( Ief95e8620a1c8ddfd6df673a3a223bd8[flogtanh_SEL-1:0]),
.flogtanh( Ic1227b130f19411495bed64035ea317b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I97455c455bbd84f8085f827abe335a75  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic1227b130f19411495bed64035ea317b };
assign I84865c4f872c0845124b78fabf695c2c = (Ief95e8620a1c8ddfd6df673a3a223bd8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I97455c455bbd84f8085f827abe335a75;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00064_00000_U (
.flogtanh_sel( I61519bc0aa02ed461dbb91851d0ae19e[flogtanh_SEL-1:0]),
.flogtanh( I6861b48d33277dd057c6f09ba630d700),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I89efdab57b5f47e1ff25b260a26b7ce0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6861b48d33277dd057c6f09ba630d700 };
assign I57b9dd7a7deea6695dcd03439c9723cf = (I61519bc0aa02ed461dbb91851d0ae19e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I89efdab57b5f47e1ff25b260a26b7ce0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00065_00000_U (
.flogtanh_sel( Ie0c11d584811174a66ca221baf87c36b[flogtanh_SEL-1:0]),
.flogtanh( I022bebca44e2f0b8f9877dd0e709b29f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9f27d55531f208c5e3b038a7e263fc48  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I022bebca44e2f0b8f9877dd0e709b29f };
assign I1cd6b35bcdfd461db69a4c1bdb1d387f = (Ie0c11d584811174a66ca221baf87c36b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9f27d55531f208c5e3b038a7e263fc48;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00066_00000_U (
.flogtanh_sel( If10f4f45ff0fd17541735934ad20f187[flogtanh_SEL-1:0]),
.flogtanh( I8e3d5a48955fe19e24975579d55f4e14),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib61c6917f61d77ed3c4a7cccf800147a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8e3d5a48955fe19e24975579d55f4e14 };
assign I40a1ecabded8add5bffe316f2d8beda9 = (If10f4f45ff0fd17541735934ad20f187[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib61c6917f61d77ed3c4a7cccf800147a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00067_00000_U (
.flogtanh_sel( I445919f07a6fa8654211301a9a6126bd[flogtanh_SEL-1:0]),
.flogtanh( I7ee915ffb1c7b8985788c5e6af532ce3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id6b11b9d84008c2444e2d5bd86e5415d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7ee915ffb1c7b8985788c5e6af532ce3 };
assign I7c52ae4af926267b5e27a530202fcce0 = (I445919f07a6fa8654211301a9a6126bd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id6b11b9d84008c2444e2d5bd86e5415d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00068_00000_U (
.flogtanh_sel( I64102b82893352549abd2e2132b19476[flogtanh_SEL-1:0]),
.flogtanh( Ia897087d82c2deac4697755c31766241),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3ee69feaef543b025d4267eb09c2cde9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia897087d82c2deac4697755c31766241 };
assign I1a5c6c50817db8bde279d5f0b5095d76 = (I64102b82893352549abd2e2132b19476[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3ee69feaef543b025d4267eb09c2cde9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00069_00000_U (
.flogtanh_sel( I1fc1933fe891ac26f35a42a1b242d919[flogtanh_SEL-1:0]),
.flogtanh( I4c23326dc80b54231289f9f18c4db711),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7ebbfe102249fcdd69f0088cd52a1fbb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4c23326dc80b54231289f9f18c4db711 };
assign Idf0c1b85712fcbbbcc12915158ebff62 = (I1fc1933fe891ac26f35a42a1b242d919[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7ebbfe102249fcdd69f0088cd52a1fbb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00070_00000_U (
.flogtanh_sel( I84dfba8bcf8ad3b85f9472fd60d607b5[flogtanh_SEL-1:0]),
.flogtanh( I8326b063a9b9688fb3014667c49ada1b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic50e81e4594d56cfd739f7f9791b1e15  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I8326b063a9b9688fb3014667c49ada1b };
assign I6b32298e8c61e75d0a38bca3084c0528 = (I84dfba8bcf8ad3b85f9472fd60d607b5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic50e81e4594d56cfd739f7f9791b1e15;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00071_00000_U (
.flogtanh_sel( I4302fccefe5ee13161f9ad49f9ddf43c[flogtanh_SEL-1:0]),
.flogtanh( Ic41133a438fcea4a1cad9f5e5ee05a03),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2968c281ccf212e6a4d456ef3e6a820e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic41133a438fcea4a1cad9f5e5ee05a03 };
assign I5b0d72cedc120406402076148e2d30b0 = (I4302fccefe5ee13161f9ad49f9ddf43c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2968c281ccf212e6a4d456ef3e6a820e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00072_00000_U (
.flogtanh_sel( I59d7153724d3b3805af799692fbe245a[flogtanh_SEL-1:0]),
.flogtanh( I1ac5e426032b874b250cb8adad5b345a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idd368451dfa1cd543cc66f44f3def824  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1ac5e426032b874b250cb8adad5b345a };
assign Iaf624549f73b0d13c1a73c850b99f810 = (I59d7153724d3b3805af799692fbe245a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idd368451dfa1cd543cc66f44f3def824;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00073_00000_U (
.flogtanh_sel( Id1650d0e39be078027493f58e9bbcbdd[flogtanh_SEL-1:0]),
.flogtanh( If9aca7e28f987bf6c7f2fb9b6f11962f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib979f9151b0b4c7c6e850780ce01cd5c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If9aca7e28f987bf6c7f2fb9b6f11962f };
assign Iaaf7efeae9f6dc9e8222dc2b10122000 = (Id1650d0e39be078027493f58e9bbcbdd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib979f9151b0b4c7c6e850780ce01cd5c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00074_00000_U (
.flogtanh_sel( If40ad4aca8dbb3bf7dde8c2ff2e5b8f2[flogtanh_SEL-1:0]),
.flogtanh( Id98a58cd8017fd149ea4f5b295f7ec80),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie3b60e864d739cc4d2c015bc0e4d85ed  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id98a58cd8017fd149ea4f5b295f7ec80 };
assign Iea1cd2321d2ac9b891b344e2ba2363d3 = (If40ad4aca8dbb3bf7dde8c2ff2e5b8f2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie3b60e864d739cc4d2c015bc0e4d85ed;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00075_00000_U (
.flogtanh_sel( Ie49f173549396caeab1d13da36e37c65[flogtanh_SEL-1:0]),
.flogtanh( Ib9e45e75ce8cdd3b548eaf3e41a091ce),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id80fb022cc3ea4d663506b98ead354a4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib9e45e75ce8cdd3b548eaf3e41a091ce };
assign Ia544fa24b953fe91800978895e3e610e = (Ie49f173549396caeab1d13da36e37c65[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id80fb022cc3ea4d663506b98ead354a4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00076_00000_U (
.flogtanh_sel( I3002a0e0cdf8e79bc7186a876410d106[flogtanh_SEL-1:0]),
.flogtanh( I9fcedcbd532cefe1e66ec94b22457cf4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I25fc15d8cb0faffee2dd7aadf733ac0e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9fcedcbd532cefe1e66ec94b22457cf4 };
assign I7fa710c37f5f96c3cdc35612a702a71c = (I3002a0e0cdf8e79bc7186a876410d106[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I25fc15d8cb0faffee2dd7aadf733ac0e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00077_00000_U (
.flogtanh_sel( I2b50fa03f584d10e9af3be085a02a12c[flogtanh_SEL-1:0]),
.flogtanh( Ic627802cf228a709638c14adf83091f8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I343f01a96adfc2286191f40a13d92ebf  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic627802cf228a709638c14adf83091f8 };
assign I98fd105696fca11c1075f9bd30013747 = (I2b50fa03f584d10e9af3be085a02a12c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I343f01a96adfc2286191f40a13d92ebf;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00078_00000_U (
.flogtanh_sel( If473d172a7bff5aeae99245bbb72978d[flogtanh_SEL-1:0]),
.flogtanh( Ib6bd27a683e11d238fcb775bb44dd913),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iab18cb1f98768ce17f46117b9a72090a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib6bd27a683e11d238fcb775bb44dd913 };
assign I61345963ceabdaa0f25f8a463fc9fe5d = (If473d172a7bff5aeae99245bbb72978d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iab18cb1f98768ce17f46117b9a72090a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00079_00000_U (
.flogtanh_sel( Ib89f7b5625995290a64bcfb143d978ca[flogtanh_SEL-1:0]),
.flogtanh( I3affcbe66b25dc7f11f98b4e444937a2),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icd8c66b0c9d66db6764cc3566a14cf06  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3affcbe66b25dc7f11f98b4e444937a2 };
assign I9e8375af6af10f4bac3e87e416d430ee = (Ib89f7b5625995290a64bcfb143d978ca[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icd8c66b0c9d66db6764cc3566a14cf06;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00080_00000_U (
.flogtanh_sel( Iebe0c9b4a87d58a1c55e2ee6b01603c4[flogtanh_SEL-1:0]),
.flogtanh( Ib537657951962c85ad92d43777458588),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I51c808cc77479f221a7c60486b75f6ed  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib537657951962c85ad92d43777458588 };
assign Ida1cd844022bbf1b8431225e66b2b78f = (Iebe0c9b4a87d58a1c55e2ee6b01603c4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I51c808cc77479f221a7c60486b75f6ed;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00081_00000_U (
.flogtanh_sel( I104411bb641d2445c7e1385a809bb682[flogtanh_SEL-1:0]),
.flogtanh( Id0af2b1d8b0aa3ba9764ea6a22fafc8c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I18a65513ce78aa9c77275103956df746  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id0af2b1d8b0aa3ba9764ea6a22fafc8c };
assign I30e9ab592e97dbc5fb6ab58d2ffbf8d4 = (I104411bb641d2445c7e1385a809bb682[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I18a65513ce78aa9c77275103956df746;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00082_00000_U (
.flogtanh_sel( I47dd28b4ae4f7151aff5bb271e35b716[flogtanh_SEL-1:0]),
.flogtanh( I3f934c17beeba9f2d2ca58b3677fe1f3),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I004491418434bb0a6a307d305df7dab0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3f934c17beeba9f2d2ca58b3677fe1f3 };
assign I2ec2a6de2be39b1bc259b0be72e35a0f = (I47dd28b4ae4f7151aff5bb271e35b716[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I004491418434bb0a6a307d305df7dab0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00083_00000_U (
.flogtanh_sel( I3a27d5573b748df459b90a5a347f9d09[flogtanh_SEL-1:0]),
.flogtanh( Ie3e094ae62dc2a694777f4792c78c886),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia74f2ce0e44e31217be3962f40588238  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie3e094ae62dc2a694777f4792c78c886 };
assign Ic32e349efae2ca419e095ee5e15a501d = (I3a27d5573b748df459b90a5a347f9d09[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia74f2ce0e44e31217be3962f40588238;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00084_00000_U (
.flogtanh_sel( I2dbef85d2b2b95af39c3a98c4e143253[flogtanh_SEL-1:0]),
.flogtanh( Idea1d2f5e910ebadc99d356dee8646bd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic92636db4722431041a6b48e99b5924d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idea1d2f5e910ebadc99d356dee8646bd };
assign I1befb935ee9cb871c9a7476c1fc0da3f = (I2dbef85d2b2b95af39c3a98c4e143253[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic92636db4722431041a6b48e99b5924d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00085_00000_U (
.flogtanh_sel( I510d39830ae7b0a857ac11baa7c144d3[flogtanh_SEL-1:0]),
.flogtanh( I7cf160bea55d67417a4ee9ce9b252871),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib525e226298f02a92a49a6fe5fcf6527  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7cf160bea55d67417a4ee9ce9b252871 };
assign I01c57f697f2af7d2c6ae904319f10725 = (I510d39830ae7b0a857ac11baa7c144d3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib525e226298f02a92a49a6fe5fcf6527;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00086_00000_U (
.flogtanh_sel( I2751a94a66ea4cb44c512df4c509937f[flogtanh_SEL-1:0]),
.flogtanh( I196915263bfb62cc21659f81572438b4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icefd1ea8daf4aaf25abd3b31256dcaa5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I196915263bfb62cc21659f81572438b4 };
assign Id580f8a2748efff9b6b747c497c16e9c = (I2751a94a66ea4cb44c512df4c509937f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icefd1ea8daf4aaf25abd3b31256dcaa5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00087_00000_U (
.flogtanh_sel( Ic9a003bfb70ac2da6c229fcad09246d4[flogtanh_SEL-1:0]),
.flogtanh( I548af5c4ccd2816978de565c0c02f176),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6f9a280cf50379308d67506d6d6a5c61  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I548af5c4ccd2816978de565c0c02f176 };
assign I77b54488bd26318f14b4364035cd1836 = (Ic9a003bfb70ac2da6c229fcad09246d4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6f9a280cf50379308d67506d6d6a5c61;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00088_00000_U (
.flogtanh_sel( I34ed986182a3311a8cb005b3dccc224b[flogtanh_SEL-1:0]),
.flogtanh( Ifb7004286169cd9b229b083aea58a408),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia4e1d880c6b384bd3b315ab453e03326  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifb7004286169cd9b229b083aea58a408 };
assign I786338397f55073dce91e1c8c5f8e298 = (I34ed986182a3311a8cb005b3dccc224b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia4e1d880c6b384bd3b315ab453e03326;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00089_00000_U (
.flogtanh_sel( Ic79281755397f6099ff30c5d07d7e6de[flogtanh_SEL-1:0]),
.flogtanh( Ib04408fcc6f4d26fcdb5599b03b1b534),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icc8d6c731fe2502a4d041cc5aefcc9d8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib04408fcc6f4d26fcdb5599b03b1b534 };
assign I0e5931219d94c8e8e1f4af081404dcab = (Ic79281755397f6099ff30c5d07d7e6de[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icc8d6c731fe2502a4d041cc5aefcc9d8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00090_00000_U (
.flogtanh_sel( I8d6559ccc33cbc663584923a55b928b5[flogtanh_SEL-1:0]),
.flogtanh( Ifda1a58a6f54318a30faa98dc1982e8e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I311ca38028cb07e4d7a8f3914aec47cc  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifda1a58a6f54318a30faa98dc1982e8e };
assign I8d96b419b010f8076311420d7b9c8a18 = (I8d6559ccc33cbc663584923a55b928b5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I311ca38028cb07e4d7a8f3914aec47cc;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00091_00000_U (
.flogtanh_sel( I4f0a4c241844e390318f11899a0f2c5a[flogtanh_SEL-1:0]),
.flogtanh( I799ce64e6df49e2b62dc6beda4500146),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I68dc05646fbd91403f254c5de1bc3c70  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I799ce64e6df49e2b62dc6beda4500146 };
assign Ife13f962c7a8df3845cde104a959f678 = (I4f0a4c241844e390318f11899a0f2c5a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I68dc05646fbd91403f254c5de1bc3c70;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00092_00000_U (
.flogtanh_sel( I45fffa266ce3838f82d755b59216a4d6[flogtanh_SEL-1:0]),
.flogtanh( Ia592b65aa89be2fcd981cf144683a298),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2550505d6e2fe478dd0c789bc3b823cf  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia592b65aa89be2fcd981cf144683a298 };
assign I7f701ff37ad3fc34d2f4efafe5ff5351 = (I45fffa266ce3838f82d755b59216a4d6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2550505d6e2fe478dd0c789bc3b823cf;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00093_00000_U (
.flogtanh_sel( I8f0e65f5db47d5460d4ec2172807a3e1[flogtanh_SEL-1:0]),
.flogtanh( Ib52365bf14aedf524bb23a4a6fe10551),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idc3ffe555b7641f987c8cc2cc2f7cb59  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib52365bf14aedf524bb23a4a6fe10551 };
assign I43c815a8ce0b2df9744a525328969691 = (I8f0e65f5db47d5460d4ec2172807a3e1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idc3ffe555b7641f987c8cc2cc2f7cb59;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00094_00000_U (
.flogtanh_sel( I34127c0d1af2438e13b6f4709ece80ba[flogtanh_SEL-1:0]),
.flogtanh( Ieba74e8bf3d692612c544af3ce6046fd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie9ab765b69fae4069793331ca0e0e5f7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ieba74e8bf3d692612c544af3ce6046fd };
assign I6c4a1ded9bf39091cf302ebe0103e2f0 = (I34127c0d1af2438e13b6f4709ece80ba[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie9ab765b69fae4069793331ca0e0e5f7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00095_00000_U (
.flogtanh_sel( I3a67de0e76bbf29d8c77c21865abda2f[flogtanh_SEL-1:0]),
.flogtanh( I6cc1587e659f3f97d636485b708b1eeb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I371fef521a66e4761eb7b3e950d6ed5c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6cc1587e659f3f97d636485b708b1eeb };
assign Icd4ff8d14af2699db2b5168027894ebb = (I3a67de0e76bbf29d8c77c21865abda2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I371fef521a66e4761eb7b3e950d6ed5c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00096_00000_U (
.flogtanh_sel( Ic64e64aeb754249b868e14311ea19759[flogtanh_SEL-1:0]),
.flogtanh( I84b09aba55d2335f19faa5762aeedb89),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6dc9b65102f0ca4eccc76b6c0321beba  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I84b09aba55d2335f19faa5762aeedb89 };
assign Ia79d52fe2130426c07890fcaa50137db = (Ic64e64aeb754249b868e14311ea19759[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6dc9b65102f0ca4eccc76b6c0321beba;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00097_00000_U (
.flogtanh_sel( Ic4aa0dc9014c8445f8d9a7723d7263f5[flogtanh_SEL-1:0]),
.flogtanh( I3c4b9082ba72cade4d52924eff135135),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If4ac2065f0165f0a22d459e53b74ba91  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3c4b9082ba72cade4d52924eff135135 };
assign I308aaa8ac500b5589aa4af533a9062bf = (Ic4aa0dc9014c8445f8d9a7723d7263f5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If4ac2065f0165f0a22d459e53b74ba91;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00098_00000_U (
.flogtanh_sel( I47b988d017580bdfe8f443904b1f3aac[flogtanh_SEL-1:0]),
.flogtanh( I65f6c14ae4e7139fd858d7637ec3fd46),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9ee4045d22e1e23f26f255e747bc2c25  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I65f6c14ae4e7139fd858d7637ec3fd46 };
assign Iac91f4037e542d9fda30fadafe7e79ac = (I47b988d017580bdfe8f443904b1f3aac[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9ee4045d22e1e23f26f255e747bc2c25;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00099_00000_U (
.flogtanh_sel( Ica9ff13e8c3850be6c70b0b06c1d9fbf[flogtanh_SEL-1:0]),
.flogtanh( I02425810db970e5ef0b791dc4be103a9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia356c2d6982d65670b4c3b276950011a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I02425810db970e5ef0b791dc4be103a9 };
assign I8cd5970682bc84881489c12ff073212c = (Ica9ff13e8c3850be6c70b0b06c1d9fbf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia356c2d6982d65670b4c3b276950011a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00100_00000_U (
.flogtanh_sel( If2efeb489911f295dd7722cb22ea521d[flogtanh_SEL-1:0]),
.flogtanh( Id0bc7b00dec58136a8016979d8a9faad),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I711a3fd75980a579031be60aa25e1da4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id0bc7b00dec58136a8016979d8a9faad };
assign I1ee27be7e1a38aff0039b21c45f406d1 = (If2efeb489911f295dd7722cb22ea521d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I711a3fd75980a579031be60aa25e1da4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00101_00000_U (
.flogtanh_sel( Iaa16dffcc01e41e6ff17e92bdefe3df5[flogtanh_SEL-1:0]),
.flogtanh( I7c61892052c3c32343ed172d4ae354cc),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I75a05a0c3ecaf5a582e01297b8dde431  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7c61892052c3c32343ed172d4ae354cc };
assign Idf90f01353ad1057e11fd060442f4e53 = (Iaa16dffcc01e41e6ff17e92bdefe3df5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I75a05a0c3ecaf5a582e01297b8dde431;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00102_00000_U (
.flogtanh_sel( Ie8857b9841fbd795a4192976ef7ecc25[flogtanh_SEL-1:0]),
.flogtanh( I7cd312338aa5a86e1b05cc28ab7a2b23),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib50109a1e4490b3bdaefc5bf87674df2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7cd312338aa5a86e1b05cc28ab7a2b23 };
assign Id45f4e0f142b6c3925f24a37dcf7c0ae = (Ie8857b9841fbd795a4192976ef7ecc25[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib50109a1e4490b3bdaefc5bf87674df2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00103_00000_U (
.flogtanh_sel( If12aef69eea28052aa3bdb6ac31af205[flogtanh_SEL-1:0]),
.flogtanh( I88d4372b4f7bfddd2af726c2df391287),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5717425e31d5707f3f1c7010cc261651  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I88d4372b4f7bfddd2af726c2df391287 };
assign I52a9bcfbd2d3a763671f19cfeaf7bb8b = (If12aef69eea28052aa3bdb6ac31af205[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5717425e31d5707f3f1c7010cc261651;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00104_00000_U (
.flogtanh_sel( I0b3c6162ae2b9221738a18a29489887f[flogtanh_SEL-1:0]),
.flogtanh( Ic8978ad86275ac6f4a0cf80ebefc5b27),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie8244d4913aa3720080a883429b5f2e3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic8978ad86275ac6f4a0cf80ebefc5b27 };
assign Ia3cc6acf2cae41e560e09993007ffd2b = (I0b3c6162ae2b9221738a18a29489887f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie8244d4913aa3720080a883429b5f2e3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00105_00000_U (
.flogtanh_sel( I08211bba29e87faf4079152bcc973e7d[flogtanh_SEL-1:0]),
.flogtanh( I99745124c45f37d3882064590394a0aa),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I32bcd4d63f2064e8b6058defcddf1523  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I99745124c45f37d3882064590394a0aa };
assign Iba0d2f08788f2208a648ae7b5414195d = (I08211bba29e87faf4079152bcc973e7d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I32bcd4d63f2064e8b6058defcddf1523;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00106_00000_U (
.flogtanh_sel( Ibff3da265f1c3f21548f5b019e1a9dc1[flogtanh_SEL-1:0]),
.flogtanh( I33fe34f9be3c51b4b93f89c3f862e332),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3d765cb8f72daad8ad6fd19b230ef2e1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I33fe34f9be3c51b4b93f89c3f862e332 };
assign I9f7df6ad60284c812aeb522974578e0b = (Ibff3da265f1c3f21548f5b019e1a9dc1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3d765cb8f72daad8ad6fd19b230ef2e1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00107_00000_U (
.flogtanh_sel( Ie9fa1762d7844b0d781afdfb0771cea9[flogtanh_SEL-1:0]),
.flogtanh( Iecda9a183e74f78b9fd5ce34e80d712e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6c50eab3042fbe8d0a9c1f13b891ca3b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iecda9a183e74f78b9fd5ce34e80d712e };
assign Iab1fb7006598181bd8749ed90c519b13 = (Ie9fa1762d7844b0d781afdfb0771cea9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6c50eab3042fbe8d0a9c1f13b891ca3b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00108_00000_U (
.flogtanh_sel( Ia677d504b9f7fc2698c0345f236428ba[flogtanh_SEL-1:0]),
.flogtanh( I5293b996bbf152abf110df1205ad4856),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7a87da6d33b578f6bc60ca0c4ee59cf5  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5293b996bbf152abf110df1205ad4856 };
assign Ieef3b299ec35075c71ef9fb10525bfc4 = (Ia677d504b9f7fc2698c0345f236428ba[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7a87da6d33b578f6bc60ca0c4ee59cf5;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00109_00000_U (
.flogtanh_sel( Idebce29121c0481df83d755b60ff632c[flogtanh_SEL-1:0]),
.flogtanh( Ia99c08ee345bdc1489ce82a62481ef3b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6ba6d7a611d9e209c8888454e1a9650e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia99c08ee345bdc1489ce82a62481ef3b };
assign I58a7c08adf48d0737c5803e2a818c045 = (Idebce29121c0481df83d755b60ff632c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6ba6d7a611d9e209c8888454e1a9650e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00110_00000_U (
.flogtanh_sel( Iad2c780a6386674d50cca54d8c4ebd86[flogtanh_SEL-1:0]),
.flogtanh( Iaa314530e04145eb73672ebb150858af),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7b6878abc6b5d1bc713bb9128c238d9d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iaa314530e04145eb73672ebb150858af };
assign I30a1c8fcd9a510a6ed559f07dd809b90 = (Iad2c780a6386674d50cca54d8c4ebd86[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7b6878abc6b5d1bc713bb9128c238d9d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00111_00000_U (
.flogtanh_sel( If1d7944e7c4828ddb91ffea28609cbc7[flogtanh_SEL-1:0]),
.flogtanh( I05f7363bfcc34691280079e82f6f5449),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3debbdfea21b3d4d975aff74df6a89a4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I05f7363bfcc34691280079e82f6f5449 };
assign Ic4f5e9d49419e1c57cfa387761ab643d = (If1d7944e7c4828ddb91ffea28609cbc7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3debbdfea21b3d4d975aff74df6a89a4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00112_00000_U (
.flogtanh_sel( I843a68ceb0adab829091f31d0de56eb6[flogtanh_SEL-1:0]),
.flogtanh( Ica5ce135e77ed1d7cbc8277344ffeaeb),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie21e2ff26b0c30eea53233d9142ec128  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ica5ce135e77ed1d7cbc8277344ffeaeb };
assign Id3dd71ea0bf0f2996fbe42b8c3318762 = (I843a68ceb0adab829091f31d0de56eb6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie21e2ff26b0c30eea53233d9142ec128;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00113_00000_U (
.flogtanh_sel( I59701b9eb54dda2744a79cebe7d73f3b[flogtanh_SEL-1:0]),
.flogtanh( Iac98c702c4d9d78460fc7c212bce7841),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9134717dde036edd9737f695d9c791ae  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iac98c702c4d9d78460fc7c212bce7841 };
assign Ib834b91bf81067e8efa9d470023e8b9d = (I59701b9eb54dda2744a79cebe7d73f3b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9134717dde036edd9737f695d9c791ae;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00114_00000_U (
.flogtanh_sel( If63cf5e8f47e4e51176401f0d954ea23[flogtanh_SEL-1:0]),
.flogtanh( I1fe269380ba03e78a8e41c17aa4bd757),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic492036079044fd3af487ee7c84e68d0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1fe269380ba03e78a8e41c17aa4bd757 };
assign Ic6ead78ed741442f17a15a157cd6ef9c = (If63cf5e8f47e4e51176401f0d954ea23[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic492036079044fd3af487ee7c84e68d0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00115_00000_U (
.flogtanh_sel( Id09454844b525697de3e3727d89551e4[flogtanh_SEL-1:0]),
.flogtanh( Ib19549130ee3307413b69c50042f7302),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib6e42f1caafaddc1c964b5b04862f5c1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib19549130ee3307413b69c50042f7302 };
assign I4e257dbd6f196a02dc0f5a2e5f6047d7 = (Id09454844b525697de3e3727d89551e4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib6e42f1caafaddc1c964b5b04862f5c1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00116_00000_U (
.flogtanh_sel( I6d1b2ce4368945b56eee7814638471cc[flogtanh_SEL-1:0]),
.flogtanh( Iad6acaf97d307fdbe0f20bf010acb468),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I54e99c231380749e3d48384c78fbf0e8  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iad6acaf97d307fdbe0f20bf010acb468 };
assign I3dbfbd34d1fdfd4f422d900154123b6b = (I6d1b2ce4368945b56eee7814638471cc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I54e99c231380749e3d48384c78fbf0e8;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00117_00000_U (
.flogtanh_sel( I6079945faa57335b1c902ccf7f960a70[flogtanh_SEL-1:0]),
.flogtanh( I67c9882f9e19df5a7b9bd0d900bb2f75),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4acf64c7b000236974dc1762d0d7223e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I67c9882f9e19df5a7b9bd0d900bb2f75 };
assign I529b763dace1924613d184c6c70c2708 = (I6079945faa57335b1c902ccf7f960a70[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4acf64c7b000236974dc1762d0d7223e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00118_00000_U (
.flogtanh_sel( Ie7752906ac55cf51f3e96e8c0046f1aa[flogtanh_SEL-1:0]),
.flogtanh( I3099768bc986a11350656e472fc21ac1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib5f05c310200a5759e4dd169a9b3ca8c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3099768bc986a11350656e472fc21ac1 };
assign I7a600aeb6cf8c3311c10afa4d82767a1 = (Ie7752906ac55cf51f3e96e8c0046f1aa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib5f05c310200a5759e4dd169a9b3ca8c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00119_00000_U (
.flogtanh_sel( I2d7d4135a94f5df949283c043228791f[flogtanh_SEL-1:0]),
.flogtanh( Ifba5972f9d38199dbc675432a29934e4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibeef99739eace0ce4d691cd2b4075571  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifba5972f9d38199dbc675432a29934e4 };
assign I8c7aab31f8cb705ea13a41a5bd349303 = (I2d7d4135a94f5df949283c043228791f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibeef99739eace0ce4d691cd2b4075571;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00120_00000_U (
.flogtanh_sel( I99c75e3d26c5d01f6ae9abcd05407d8c[flogtanh_SEL-1:0]),
.flogtanh( I0934fb292b19451a050fb3374a7bd1a7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iea5ee3bf75ed967ef2dfc8ed8d9bbc2f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0934fb292b19451a050fb3374a7bd1a7 };
assign I171149dcaab2c0f0e2a10547ad95084d = (I99c75e3d26c5d01f6ae9abcd05407d8c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iea5ee3bf75ed967ef2dfc8ed8d9bbc2f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00121_00000_U (
.flogtanh_sel( I81e6f97621dbfb2fed6fc236005a2b19[flogtanh_SEL-1:0]),
.flogtanh( I9a3d1741c77fb1bbc1a54383874de82a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib10b3fb9882f1a07acee84ad15ad21f1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9a3d1741c77fb1bbc1a54383874de82a };
assign I23b60ca4da2df0ec40c1df62d058deef = (I81e6f97621dbfb2fed6fc236005a2b19[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib10b3fb9882f1a07acee84ad15ad21f1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00122_00000_U (
.flogtanh_sel( Ieac60532dcfc916a65054e35cf31d6d2[flogtanh_SEL-1:0]),
.flogtanh( If89f2ce813bab91af88f73ddc570d5a1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7a74e6f3e2acbd05e92ff91cc8771f91  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If89f2ce813bab91af88f73ddc570d5a1 };
assign I7978d2d800b4438d0644ae3df6bcac9c = (Ieac60532dcfc916a65054e35cf31d6d2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7a74e6f3e2acbd05e92ff91cc8771f91;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00123_00000_U (
.flogtanh_sel( Ib7eb83ba73e0dc17f69c357b6ca555bf[flogtanh_SEL-1:0]),
.flogtanh( Ibc0dfcffac26f4898d42808534f6588f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8f718fbf0d8b43af7002b67f6e0ef202  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibc0dfcffac26f4898d42808534f6588f };
assign Ibc4eddc0f1768e9ec7e38e951a28ec42 = (Ib7eb83ba73e0dc17f69c357b6ca555bf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8f718fbf0d8b43af7002b67f6e0ef202;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00124_00000_U (
.flogtanh_sel( I5139d8a7a099e3c619c60647c15b7420[flogtanh_SEL-1:0]),
.flogtanh( I3a0a6f3d0141e8ad04d89c4bf306a96f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3bf775756dc497fa91654eb7cf0657e9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3a0a6f3d0141e8ad04d89c4bf306a96f };
assign I1c97fd1d21a31af8b5498a79b1a3e7b6 = (I5139d8a7a099e3c619c60647c15b7420[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3bf775756dc497fa91654eb7cf0657e9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00125_00000_U (
.flogtanh_sel( I6ccd2e11ebd5b2de80b120e20650a602[flogtanh_SEL-1:0]),
.flogtanh( I1c875571dd1be1bb28aa15554964b485),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7c6d4cac0d6ff029d636fa006aa59912  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1c875571dd1be1bb28aa15554964b485 };
assign Ie4f063eeaf7ee3f033e2a01ffaca623e = (I6ccd2e11ebd5b2de80b120e20650a602[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7c6d4cac0d6ff029d636fa006aa59912;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00126_00000_U (
.flogtanh_sel( Ie669cebe5fe39e1a841f8dd3c1f6bc57[flogtanh_SEL-1:0]),
.flogtanh( Ide5d5fdcf86b369b015890030a222a0a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I46249ffce3ba1abfbaaf1447070c1990  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ide5d5fdcf86b369b015890030a222a0a };
assign Ibb3d57d510cad00064a331f61f6400a2 = (Ie669cebe5fe39e1a841f8dd3c1f6bc57[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I46249ffce3ba1abfbaaf1447070c1990;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00127_00000_U (
.flogtanh_sel( If32acb9fc212c4af34099acf6df2bc5a[flogtanh_SEL-1:0]),
.flogtanh( I7cf6e8d40e7bd7685a7260638523690c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I13b24152d7160e4e4c0b8de8ca43ce6a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7cf6e8d40e7bd7685a7260638523690c };
assign I9485ae915474a31562ce358666d66245 = (If32acb9fc212c4af34099acf6df2bc5a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I13b24152d7160e4e4c0b8de8ca43ce6a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00128_00000_U (
.flogtanh_sel( I075ce236a181bf925c8ccce91d9bc8cd[flogtanh_SEL-1:0]),
.flogtanh( I52ccac771cc9a1c1797862bc781e1f58),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If1d125c997fc331af17a03fa647c3a1e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I52ccac771cc9a1c1797862bc781e1f58 };
assign Ia54b6f7044a831020e49f1bf48bc063a = (I075ce236a181bf925c8ccce91d9bc8cd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If1d125c997fc331af17a03fa647c3a1e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00129_00000_U (
.flogtanh_sel( I541d4e422b999a0dfca44d275178e1d9[flogtanh_SEL-1:0]),
.flogtanh( I9db2090916f2535b14ed3292e78baa32),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id02c9cea3b4048f89cdb011325b5f874  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9db2090916f2535b14ed3292e78baa32 };
assign Ie71c7babb5d17378d40444b6bbd4e7a6 = (I541d4e422b999a0dfca44d275178e1d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id02c9cea3b4048f89cdb011325b5f874;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00130_00000_U (
.flogtanh_sel( I3e02657f3d9f79338cd083ed024bf96c[flogtanh_SEL-1:0]),
.flogtanh( I5b77a8ce7f495ae61315d1590bfd71b8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaabab9f3f0c05d0d5fba679bbcb14b3d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5b77a8ce7f495ae61315d1590bfd71b8 };
assign Ia0977b79857bdbf058535c30e338c38a = (I3e02657f3d9f79338cd083ed024bf96c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaabab9f3f0c05d0d5fba679bbcb14b3d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00131_00000_U (
.flogtanh_sel( Ia5e5537405ab8edcc7cd43c86837d43d[flogtanh_SEL-1:0]),
.flogtanh( I4e4bb795cf09757c8ad3933c9ce4686f),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2bfaf258762bbc682298a56d3092d369  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4e4bb795cf09757c8ad3933c9ce4686f };
assign I600ea1371a2be66430ac9534583b512b = (Ia5e5537405ab8edcc7cd43c86837d43d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2bfaf258762bbc682298a56d3092d369;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00132_00000_U (
.flogtanh_sel( I07ff388e3b6c7288f0f6c35a345023fe[flogtanh_SEL-1:0]),
.flogtanh( I78c29808e737dab48b5144b232dd02f6),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If15b5be646c24f6e8ab29b0b7646ebe0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I78c29808e737dab48b5144b232dd02f6 };
assign Ife5b9afdbb30c122b84d5378f9cb366d = (I07ff388e3b6c7288f0f6c35a345023fe[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If15b5be646c24f6e8ab29b0b7646ebe0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00133_00000_U (
.flogtanh_sel( I56cb3b3e193ca5068734417fd0ec4e02[flogtanh_SEL-1:0]),
.flogtanh( Ie2ae83a457d79fbddc640d49d626171c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I58a4e50090f1a5028e267e31bf7c2e00  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie2ae83a457d79fbddc640d49d626171c };
assign I27556d599dd1a27ee8f49e819ccbf29a = (I56cb3b3e193ca5068734417fd0ec4e02[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I58a4e50090f1a5028e267e31bf7c2e00;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00134_00000_U (
.flogtanh_sel( I5bbf1765d8f81581d0cf31c0bc755fb3[flogtanh_SEL-1:0]),
.flogtanh( I3711e49a4eec517e47897fb731d75958),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2f87ae03574e521a6911a4dcd3dc4ec3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3711e49a4eec517e47897fb731d75958 };
assign Icce595233ce089eafcca3eae5e71e5f8 = (I5bbf1765d8f81581d0cf31c0bc755fb3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2f87ae03574e521a6911a4dcd3dc4ec3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00135_00000_U (
.flogtanh_sel( Iaa1643095e518846cdede4d5a90dff84[flogtanh_SEL-1:0]),
.flogtanh( Ifda4e727eb6275266f583badb6d4a9ed),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I84e1a5675d75723d7c5fd8ec7a8bd093  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifda4e727eb6275266f583badb6d4a9ed };
assign Icc3cadf40c09be1a8c2847caf0e3e63c = (Iaa1643095e518846cdede4d5a90dff84[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I84e1a5675d75723d7c5fd8ec7a8bd093;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00136_00000_U (
.flogtanh_sel( Iee6e12f4717a3279dd31b874eabae69e[flogtanh_SEL-1:0]),
.flogtanh( I2be66a82c7b58e3c14b5816522b46969),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I905aab3b31d9dd6fecb74ede9f4c56c0  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2be66a82c7b58e3c14b5816522b46969 };
assign Ib43886d923b8c683004713ff25b2f90d = (Iee6e12f4717a3279dd31b874eabae69e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I905aab3b31d9dd6fecb74ede9f4c56c0;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00137_00000_U (
.flogtanh_sel( Ic52a9edbbc5283844d2514ea142ca6e2[flogtanh_SEL-1:0]),
.flogtanh( I826fe7ad9e67061800d5d6543d779864),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I66d3f7876f1fdc9a4d753a3bbd462300  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I826fe7ad9e67061800d5d6543d779864 };
assign I132d9671c582876568c0f7f5335f5227 = (Ic52a9edbbc5283844d2514ea142ca6e2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I66d3f7876f1fdc9a4d753a3bbd462300;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00138_00000_U (
.flogtanh_sel( Ice3e978c8da2a7de5b28542a5589f0a2[flogtanh_SEL-1:0]),
.flogtanh( Ic0c9069041758b53f56a46da81dd2d60),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3cd15e755f29b592bf2c1532e86d8f33  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic0c9069041758b53f56a46da81dd2d60 };
assign I0859c80b42a8c60dade8f05d58ee3701 = (Ice3e978c8da2a7de5b28542a5589f0a2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3cd15e755f29b592bf2c1532e86d8f33;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00139_00000_U (
.flogtanh_sel( I336a425aed221c85ca80b9a97d21d6b1[flogtanh_SEL-1:0]),
.flogtanh( I6f4c5a8de7690fec959861f43c134915),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I14423aefbe6d66dbd2f518ae34f43f61  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6f4c5a8de7690fec959861f43c134915 };
assign Ib3690ec149adde94343d3e617931a287 = (I336a425aed221c85ca80b9a97d21d6b1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I14423aefbe6d66dbd2f518ae34f43f61;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00140_00000_U (
.flogtanh_sel( Ie477c0f3b77bb299ba8b1a410d211ef7[flogtanh_SEL-1:0]),
.flogtanh( I14f1005a8c0fbdc5ca02c032b8891c2b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib1331d92ac9a84842b3e1b81968f241c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I14f1005a8c0fbdc5ca02c032b8891c2b };
assign I41f2bf9ff00f983ad1298c8c83b041cb = (Ie477c0f3b77bb299ba8b1a410d211ef7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib1331d92ac9a84842b3e1b81968f241c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00141_00000_U (
.flogtanh_sel( Ie62920d089ae762603cd33fbf97d92bb[flogtanh_SEL-1:0]),
.flogtanh( Iacd30dfb96f6572ec56eff0a4094ec04),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If5d175d3ad99e5f1a37ca02c5b72b550  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Iacd30dfb96f6572ec56eff0a4094ec04 };
assign Ib5414585cd6976cfce42e42190cc08d7 = (Ie62920d089ae762603cd33fbf97d92bb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If5d175d3ad99e5f1a37ca02c5b72b550;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00142_00000_U (
.flogtanh_sel( I2ca952e4e676537fd5a8fc71ecfa10e9[flogtanh_SEL-1:0]),
.flogtanh( I1c748b8fe4979331bc3fe5aff4b6f9f4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I44e3174343cfa4f55b79f77e80005fbb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1c748b8fe4979331bc3fe5aff4b6f9f4 };
assign I1ca59325ff30db83df5bf0a2cd9706b6 = (I2ca952e4e676537fd5a8fc71ecfa10e9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I44e3174343cfa4f55b79f77e80005fbb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00143_00000_U (
.flogtanh_sel( Iefd31e7ff3c829c88f60bc89d70afcf7[flogtanh_SEL-1:0]),
.flogtanh( I158c7973974f36c2793127964e50d1bd),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7d917703c26558414d5fb997398a8757  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I158c7973974f36c2793127964e50d1bd };
assign Ie2f5b03f3b136e651b8aba92a30d298a = (Iefd31e7ff3c829c88f60bc89d70afcf7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7d917703c26558414d5fb997398a8757;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00144_00000_U (
.flogtanh_sel( Iafa987a413fd8fcacfe872bc0f5bc2d6[flogtanh_SEL-1:0]),
.flogtanh( Id5ea6ba2402275cb925a1848b31ec2e1),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5ff9bb8ef0620b2a968cc99b709723c7  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id5ea6ba2402275cb925a1848b31ec2e1 };
assign I312ce79a8dd2ce3d37c930d42640509b = (Iafa987a413fd8fcacfe872bc0f5bc2d6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5ff9bb8ef0620b2a968cc99b709723c7;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00145_00000_U (
.flogtanh_sel( I305c1ea420d666f258e38c5a65847367[flogtanh_SEL-1:0]),
.flogtanh( I3862f7017bc2bc69844b73f2a79f47f5),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icb83a6adcf84370776ad71a9f5a8735b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3862f7017bc2bc69844b73f2a79f47f5 };
assign I467d5e2554ef25873e0b44e947ee0011 = (I305c1ea420d666f258e38c5a65847367[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icb83a6adcf84370776ad71a9f5a8735b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00146_00000_U (
.flogtanh_sel( I9f040c4088bfab72d74e5332e9710d1a[flogtanh_SEL-1:0]),
.flogtanh( I4ed41fde5449b7112baf000a05484ac4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieaa23d9c0997f273064a57b8071c64c1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4ed41fde5449b7112baf000a05484ac4 };
assign Ice73b514709469fd21cd254bf4ceadd9 = (I9f040c4088bfab72d74e5332e9710d1a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieaa23d9c0997f273064a57b8071c64c1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00147_00000_U (
.flogtanh_sel( Ia2f41f9778324a06daeb185c736516a4[flogtanh_SEL-1:0]),
.flogtanh( I40c4db2872b602bf9d6a4fc4ba5ac34d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I69b89cf26b64d319f7796610e92caec9  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I40c4db2872b602bf9d6a4fc4ba5ac34d };
assign I45ba06a6d6f00c174b1439a6f226a085 = (Ia2f41f9778324a06daeb185c736516a4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I69b89cf26b64d319f7796610e92caec9;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00148_00000_U (
.flogtanh_sel( Id9778ba5fbdbed4d33a092da6b68c414[flogtanh_SEL-1:0]),
.flogtanh( Ibe5ab52bd0f220f7a6aac244c0e3867e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6bf4038fafaa59349f73aa011149067e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibe5ab52bd0f220f7a6aac244c0e3867e };
assign Ic8a272f82736fd599fb3250e970edf9b = (Id9778ba5fbdbed4d33a092da6b68c414[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6bf4038fafaa59349f73aa011149067e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00149_00000_U (
.flogtanh_sel( I27c2c79d0d719c71c8e28218d1174a13[flogtanh_SEL-1:0]),
.flogtanh( I36668064f280c70f9143ee9f39973015),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idbe16e45feac2ab46cd58d32eb0e3113  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I36668064f280c70f9143ee9f39973015 };
assign I5b9710b16effc8bf0695517c6e651836 = (I27c2c79d0d719c71c8e28218d1174a13[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idbe16e45feac2ab46cd58d32eb0e3113;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00150_00000_U (
.flogtanh_sel( I2a9d6a774769b12ae20bc0cee0c36f5c[flogtanh_SEL-1:0]),
.flogtanh( Ief92462253c5a03a42d46ed7087caf9a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I11eb91a1ff576ec2787ec76b0787977c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ief92462253c5a03a42d46ed7087caf9a };
assign I038b42a83025f5eaebf45799d1ebe7b0 = (I2a9d6a774769b12ae20bc0cee0c36f5c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I11eb91a1ff576ec2787ec76b0787977c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00151_00000_U (
.flogtanh_sel( I2c567b75f1399c069b95284f4c36b6d1[flogtanh_SEL-1:0]),
.flogtanh( Idf196345491ff3290796ba7827d31c17),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie45dede493b6ce54a123db34cfedcefe  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Idf196345491ff3290796ba7827d31c17 };
assign I73ddd7cf9272ceab5a663e2244e72d7e = (I2c567b75f1399c069b95284f4c36b6d1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie45dede493b6ce54a123db34cfedcefe;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00152_00000_U (
.flogtanh_sel( If3d3eb609abfd6e315eec803d2e94490[flogtanh_SEL-1:0]),
.flogtanh( I2230f0e48899877bc2bcb3538be81bfa),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I69df2773462a5c7a2802176217eeee01  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I2230f0e48899877bc2bcb3538be81bfa };
assign I16507fab8f9076bfeb419896fa7cdc1d = (If3d3eb609abfd6e315eec803d2e94490[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I69df2773462a5c7a2802176217eeee01;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00153_00000_U (
.flogtanh_sel( I9c58aea7ce986b1d28f5808b347c015d[flogtanh_SEL-1:0]),
.flogtanh( Ibc0ec83d6b8e6be89ddc88ef83f0b03d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id8a3ef0da815bdd206d02be6d7b82c89  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibc0ec83d6b8e6be89ddc88ef83f0b03d };
assign I3dd1f28cf199299aba54e47a429c9b11 = (I9c58aea7ce986b1d28f5808b347c015d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id8a3ef0da815bdd206d02be6d7b82c89;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00154_00000_U (
.flogtanh_sel( Id139c7a783196941100003b6cb0cd1e7[flogtanh_SEL-1:0]),
.flogtanh( Ifc59c1b26ec09b3a7fe5a2b90511c93b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9f74767b10d0981465160f7f9c915826  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifc59c1b26ec09b3a7fe5a2b90511c93b };
assign I49d9203dc6f8c17f17383e8f7e01f005 = (Id139c7a783196941100003b6cb0cd1e7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9f74767b10d0981465160f7f9c915826;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00155_00000_U (
.flogtanh_sel( I524d7614b01460778da3ce98f6aaa3d9[flogtanh_SEL-1:0]),
.flogtanh( I9c6fc8e09cd63551f40accc98d784a44),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6340b82b10836e90efc17d3d8ce27aa4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9c6fc8e09cd63551f40accc98d784a44 };
assign Ibeec86c75d950ee00dd63a2930f08a24 = (I524d7614b01460778da3ce98f6aaa3d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6340b82b10836e90efc17d3d8ce27aa4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00156_00000_U (
.flogtanh_sel( I8acda65f116d5c91cbe2662ac282aa31[flogtanh_SEL-1:0]),
.flogtanh( I26692a6aab1d81d71219a436bee5e10b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ief2d5177fa9a28016b5da2def9de4050  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I26692a6aab1d81d71219a436bee5e10b };
assign I47b2438c3680b2d816168df37d7c491c = (I8acda65f116d5c91cbe2662ac282aa31[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ief2d5177fa9a28016b5da2def9de4050;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00157_00000_U (
.flogtanh_sel( If67dbe22f8d22b3430215fb0deae8204[flogtanh_SEL-1:0]),
.flogtanh( Ieb50592e17305d0f74cbf216be947862),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I49214ecffd1e025db688d04119248a84  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ieb50592e17305d0f74cbf216be947862 };
assign I5983bf2c6c90b872ee6cf58b5e520311 = (If67dbe22f8d22b3430215fb0deae8204[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I49214ecffd1e025db688d04119248a84;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00158_00000_U (
.flogtanh_sel( I9a35cd7512787263abedd6d9913cf507[flogtanh_SEL-1:0]),
.flogtanh( I0071f023f1be4400541c13bc68278417),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icb84682ddc30efd01dcfe2d96a84ba9d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0071f023f1be4400541c13bc68278417 };
assign I6745cacecb7ee86cf3c7ad7eeee6048f = (I9a35cd7512787263abedd6d9913cf507[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icb84682ddc30efd01dcfe2d96a84ba9d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00159_00000_U (
.flogtanh_sel( If9cca23469c5e6001650f1f8b1360ae8[flogtanh_SEL-1:0]),
.flogtanh( Ib2f1635b38ca6090e5ff633cbfa13273),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7f99c71ccc1918b7ee0ca2e9ed84ea17  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib2f1635b38ca6090e5ff633cbfa13273 };
assign Ib9672d20643d856ff31905ab14c0ac87 = (If9cca23469c5e6001650f1f8b1360ae8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7f99c71ccc1918b7ee0ca2e9ed84ea17;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00160_00000_U (
.flogtanh_sel( Icc2606ae8f9a3b425225ae7339112b9d[flogtanh_SEL-1:0]),
.flogtanh( Id2c0bc90fd26e82fe91b5aef7bdd3a29),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifbc9e59e2ea7b320ad2ec483bd58c1c4  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id2c0bc90fd26e82fe91b5aef7bdd3a29 };
assign Ib9dfea1f34a120eda30d5bd919365a6a = (Icc2606ae8f9a3b425225ae7339112b9d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifbc9e59e2ea7b320ad2ec483bd58c1c4;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00161_00000_U (
.flogtanh_sel( I34aa1802d24e074ae54563898929abfa[flogtanh_SEL-1:0]),
.flogtanh( If4a723ce836f5327b85e234ebd195bd9),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I98a7d5627114777569c3ad29fbdf33ce  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If4a723ce836f5327b85e234ebd195bd9 };
assign Ia7bf82c9e5ca4467b5e50beeaeb975e9 = (I34aa1802d24e074ae54563898929abfa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I98a7d5627114777569c3ad29fbdf33ce;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00162_00000_U (
.flogtanh_sel( Icb85b3464dc40e8504c53c377e889c45[flogtanh_SEL-1:0]),
.flogtanh( If63dd5997e033817126a9ebaf38c1955),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic3cf4882216f4f3c63524154ca5bf020  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, If63dd5997e033817126a9ebaf38c1955 };
assign I327c9acb8934729b4ea5486787afa2e8 = (Icb85b3464dc40e8504c53c377e889c45[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic3cf4882216f4f3c63524154ca5bf020;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00163_00000_U (
.flogtanh_sel( Ie595a7d10b5ac84c0301fb55bebd3680[flogtanh_SEL-1:0]),
.flogtanh( Ie2ee6baf8ec357f6131dff92fb480e42),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaa2e0df90fb601ebaddcf0d4afaeedd2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie2ee6baf8ec357f6131dff92fb480e42 };
assign Ieddef08050c38d07e5d38f5bb7b099c0 = (Ie595a7d10b5ac84c0301fb55bebd3680[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaa2e0df90fb601ebaddcf0d4afaeedd2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00164_00000_U (
.flogtanh_sel( I9c217a672cabc05efbdff218637123ba[flogtanh_SEL-1:0]),
.flogtanh( Ibff4d4fca3681fe10807414ed84e4157),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0f5bf0ab35c2588426d461588a882388  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibff4d4fca3681fe10807414ed84e4157 };
assign I39f9e8430db114991bfb27cc46ef3e39 = (I9c217a672cabc05efbdff218637123ba[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0f5bf0ab35c2588426d461588a882388;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00165_00000_U (
.flogtanh_sel( If20f3780b4af857ffe8083056085517a[flogtanh_SEL-1:0]),
.flogtanh( I4540d74c919f50e9b6e40ef6b8cfd279),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic7fc2a5137184b1908cb1293341fcf26  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4540d74c919f50e9b6e40ef6b8cfd279 };
assign I56aa548618a4a15e9a35e04f5eeb823f = (If20f3780b4af857ffe8083056085517a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic7fc2a5137184b1908cb1293341fcf26;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00166_00000_U (
.flogtanh_sel( Ic2e275bfa8ab3d2002d2aa374ac9bfe2[flogtanh_SEL-1:0]),
.flogtanh( I01637ffca829d72accbb5dcee48817ca),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0e1b866232599fcb497ce38c2c68f32a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I01637ffca829d72accbb5dcee48817ca };
assign I1908897b529ca04df7e7da395be4a8ce = (Ic2e275bfa8ab3d2002d2aa374ac9bfe2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0e1b866232599fcb497ce38c2c68f32a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00167_00000_U (
.flogtanh_sel( Iac5798fd9915b6778700da6a14f6a381[flogtanh_SEL-1:0]),
.flogtanh( I7e8af960e934c7cc3cb163d6f8e7d597),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id526a3d6594056c40bd5c1ee1f109925  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7e8af960e934c7cc3cb163d6f8e7d597 };
assign Ib2bbd59cd6098608ed53ac556036534f = (Iac5798fd9915b6778700da6a14f6a381[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id526a3d6594056c40bd5c1ee1f109925;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00168_00000_U (
.flogtanh_sel( Ide3204bf317fdfb993410d338085b174[flogtanh_SEL-1:0]),
.flogtanh( Ifd80d371c8851b9e16193a3e62ddf79a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia75d451c04e28eb476104090e9f952b2  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifd80d371c8851b9e16193a3e62ddf79a };
assign If004552b2047ab1cf23bb50375460b01 = (Ide3204bf317fdfb993410d338085b174[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia75d451c04e28eb476104090e9f952b2;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00169_00000_U (
.flogtanh_sel( Ic3a95140fc1029efa17a6557bc977719[flogtanh_SEL-1:0]),
.flogtanh( I19d2c4bc969133fa59d22f7f2d8cfd4a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib30ec3e9a870536690a38fe069018f42  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I19d2c4bc969133fa59d22f7f2d8cfd4a };
assign If97092e1e2147de199c94a23831cf6b9 = (Ic3a95140fc1029efa17a6557bc977719[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib30ec3e9a870536690a38fe069018f42;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00170_00000_U (
.flogtanh_sel( I647d3a46bb2c7ed0f1ec08760b3858be[flogtanh_SEL-1:0]),
.flogtanh( I532326ad245909d441134296dae9a5d4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I00edc092e1c7c9738943465938a693bd  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I532326ad245909d441134296dae9a5d4 };
assign Ibf74a4dfaab7f7f538d2b5fac7394b63 = (I647d3a46bb2c7ed0f1ec08760b3858be[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I00edc092e1c7c9738943465938a693bd;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00171_00000_U (
.flogtanh_sel( I4816747af9d9fc8dc85fd831336ec710[flogtanh_SEL-1:0]),
.flogtanh( I6ca7199e28b480ac5816bf5b4cfb1eef),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4dc8aa3d45b1cbb2a926179a5cccdf57  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I6ca7199e28b480ac5816bf5b4cfb1eef };
assign I991a7a7d562eb0a8b4b8d8f008ef2225 = (I4816747af9d9fc8dc85fd831336ec710[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4dc8aa3d45b1cbb2a926179a5cccdf57;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00172_00000_U (
.flogtanh_sel( I1f66c026a5437320bd1f4df2ff71663d[flogtanh_SEL-1:0]),
.flogtanh( I0d5b26d24fbce6b236120b5697d0db6b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4a60dfcad5fab348684831c1c5301d02  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0d5b26d24fbce6b236120b5697d0db6b };
assign I64c3d7be41abaa17d6992f9af8e72789 = (I1f66c026a5437320bd1f4df2ff71663d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4a60dfcad5fab348684831c1c5301d02;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00173_00000_U (
.flogtanh_sel( If347c58c328193f420286ea27a4afa20[flogtanh_SEL-1:0]),
.flogtanh( I618d329f2b0f18617d80aa350b79601c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6d9fce52b1224fa10ee9bd3e5a02b68b  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I618d329f2b0f18617d80aa350b79601c };
assign Icb91e63ebabc7a75a54eb7c731df4fa0 = (If347c58c328193f420286ea27a4afa20[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6d9fce52b1224fa10ee9bd3e5a02b68b;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00174_00000_U (
.flogtanh_sel( I7a126c8304be920f2a920315dc61ba7f[flogtanh_SEL-1:0]),
.flogtanh( I58e3a5e842e14d09de91959839798a67),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifcc8638ec8cc700bfafedd844eabe861  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I58e3a5e842e14d09de91959839798a67 };
assign I673d1d0d0daab99bd940c46cc14ef55a = (I7a126c8304be920f2a920315dc61ba7f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifcc8638ec8cc700bfafedd844eabe861;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00175_00000_U (
.flogtanh_sel( I237327d6a74df1fb05537dc3691ebf11[flogtanh_SEL-1:0]),
.flogtanh( Icdecd5095ef818a0915ff3fcb395db5b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I60914917663174bf0a5f6b1b16a0a1ce  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Icdecd5095ef818a0915ff3fcb395db5b };
assign I62cadbd70b07a6a7a2974c7c392696b3 = (I237327d6a74df1fb05537dc3691ebf11[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I60914917663174bf0a5f6b1b16a0a1ce;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00176_00000_U (
.flogtanh_sel( I64a3e8bb4c87b066806d33a5306a2c53[flogtanh_SEL-1:0]),
.flogtanh( I236f843994d3065b6ee70c41f390a3d0),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4ef6d192effc3fb6d583b0370194cd62  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I236f843994d3065b6ee70c41f390a3d0 };
assign Icd8257d7f53d93db989eb56eaeb7e593 = (I64a3e8bb4c87b066806d33a5306a2c53[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4ef6d192effc3fb6d583b0370194cd62;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00177_00000_U (
.flogtanh_sel( Ibbca6ec39234473fb517447a8beacafc[flogtanh_SEL-1:0]),
.flogtanh( I7a9001d6c1d1aa8af79d9b152e596b70),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9fe9281eeaac31b7c9499f5c3e8bfe9a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7a9001d6c1d1aa8af79d9b152e596b70 };
assign I05931ceae6eff26e5a66a44a54d628ae = (Ibbca6ec39234473fb517447a8beacafc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9fe9281eeaac31b7c9499f5c3e8bfe9a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00178_00000_U (
.flogtanh_sel( I78327356176a16fc996188b83b058cbc[flogtanh_SEL-1:0]),
.flogtanh( I56a43a072d463792d9e676c4907b3e76),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I80bc60c27d0ebfc778d59b578732f07e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I56a43a072d463792d9e676c4907b3e76 };
assign I306fec0aa68a0396053a6e0fa1cda38f = (I78327356176a16fc996188b83b058cbc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I80bc60c27d0ebfc778d59b578732f07e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00179_00000_U (
.flogtanh_sel( Ifec496c87a7a2474855067305ac8cba3[flogtanh_SEL-1:0]),
.flogtanh( I336a86e85d3a8a42c4b6458ccb92ae05),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id371abee85a8611bc9f15cb475c76169  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I336a86e85d3a8a42c4b6458ccb92ae05 };
assign Idee8c8144207d676d1f2f9064bbdff45 = (Ifec496c87a7a2474855067305ac8cba3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id371abee85a8611bc9f15cb475c76169;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00180_00000_U (
.flogtanh_sel( I41584165a62caaa37ddebbf79bb8b617[flogtanh_SEL-1:0]),
.flogtanh( Id97f66b78f1e3b6bf0b962b85ca1cde7),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ida40585da3f7140c84ef2d0088d42977  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id97f66b78f1e3b6bf0b962b85ca1cde7 };
assign I5855124d566af739caa6511f8598f2c5 = (I41584165a62caaa37ddebbf79bb8b617[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ida40585da3f7140c84ef2d0088d42977;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00181_00000_U (
.flogtanh_sel( Idf0916d6b025aad6eccb98ada5ba3aca[flogtanh_SEL-1:0]),
.flogtanh( I52c7f0a8f9b4533052b5acd1b5bd5e17),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib175445b5c07a6fd6e4ea0dc6e6952fe  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I52c7f0a8f9b4533052b5acd1b5bd5e17 };
assign I50729db4a8e04f18979707df14cb2419 = (Idf0916d6b025aad6eccb98ada5ba3aca[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib175445b5c07a6fd6e4ea0dc6e6952fe;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00182_00000_U (
.flogtanh_sel( I00ef133d5a53f8f99f35b50327e5272b[flogtanh_SEL-1:0]),
.flogtanh( I3b1db672b1a94502b90451260062a274),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idb001650555c8e77733c2cae7b6f099f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I3b1db672b1a94502b90451260062a274 };
assign Ia3cb3ea64576a3e7332e1fb55953aa3e = (I00ef133d5a53f8f99f35b50327e5272b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idb001650555c8e77733c2cae7b6f099f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00183_00000_U (
.flogtanh_sel( I6f0e302d38d75982d0761e306ce9f146[flogtanh_SEL-1:0]),
.flogtanh( I1a83f91eb1262911ae8d99e305294bf8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icfa6a05bc48790590b66ff78773cc9a6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I1a83f91eb1262911ae8d99e305294bf8 };
assign I3cb1f233951d49f985b0deac6e052bfd = (I6f0e302d38d75982d0761e306ce9f146[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icfa6a05bc48790590b66ff78773cc9a6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00184_00000_U (
.flogtanh_sel( I127eed5de00e10a020717e796de76c7d[flogtanh_SEL-1:0]),
.flogtanh( Id01bfbd86b6321a843e239ca97cec514),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib953adc95f33e5f0f97545b7ac0e6a82  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Id01bfbd86b6321a843e239ca97cec514 };
assign I7015def91103398e54f446ce3e43af01 = (I127eed5de00e10a020717e796de76c7d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib953adc95f33e5f0f97545b7ac0e6a82;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00185_00000_U (
.flogtanh_sel( If9aad73aefb1b225f35e8c813b85fe87[flogtanh_SEL-1:0]),
.flogtanh( I26b769b58e1c21b68dd95c9f38c0362b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3e379d83cf4dae9968eaadd4da9e2b4c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I26b769b58e1c21b68dd95c9f38c0362b };
assign I04874bd1bf257f205b5189c8c20e5a12 = (If9aad73aefb1b225f35e8c813b85fe87[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3e379d83cf4dae9968eaadd4da9e2b4c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00186_00000_U (
.flogtanh_sel( I00a89ac37676521a081a21b1ec1a0798[flogtanh_SEL-1:0]),
.flogtanh( Ic86f9988281398adfe43152beb722c1b),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I51508292b5316d23e45d217d48eb623d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic86f9988281398adfe43152beb722c1b };
assign I937e3a8ede2305ea7c1750283224a870 = (I00a89ac37676521a081a21b1ec1a0798[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I51508292b5316d23e45d217d48eb623d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00187_00000_U (
.flogtanh_sel( I06f3a34f2b1770ef82ddc2a732b3d4fb[flogtanh_SEL-1:0]),
.flogtanh( I9d8ac6c29c2f5df7c2d124dface59e35),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I36d727f90d4a830f79443b4941c9df9c  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9d8ac6c29c2f5df7c2d124dface59e35 };
assign Ia7206430a739a11af4d860096eedd6c3 = (I06f3a34f2b1770ef82ddc2a732b3d4fb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I36d727f90d4a830f79443b4941c9df9c;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00188_00000_U (
.flogtanh_sel( I4744d64a746f16004e3bedaaa41465f1[flogtanh_SEL-1:0]),
.flogtanh( I56b46c426895409b40c3be9b79365a8a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I519b932add092db1a149df22a471d04e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I56b46c426895409b40c3be9b79365a8a };
assign Ibf4c2c00f8e012e9498361bfd3c5b06e = (I4744d64a746f16004e3bedaaa41465f1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I519b932add092db1a149df22a471d04e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00189_00000_U (
.flogtanh_sel( Ifae0cc6cc1c65d24bbe84c4ba938e2ea[flogtanh_SEL-1:0]),
.flogtanh( Ic63de8464f79ae05f27f05c935dbf495),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I44395e9b406cd0ae7b3672e8ff86af4d  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ic63de8464f79ae05f27f05c935dbf495 };
assign I899e5f03cd1d52d11f898959559aaeea = (Ifae0cc6cc1c65d24bbe84c4ba938e2ea[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I44395e9b406cd0ae7b3672e8ff86af4d;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00190_00000_U (
.flogtanh_sel( I1223c21129382d41e4f38ef4bbe60c2f[flogtanh_SEL-1:0]),
.flogtanh( I4d21ee443e5921532d5bf1db7ef93f82),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I08955fcfabffed0ad0c5e398e7872be1  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I4d21ee443e5921532d5bf1db7ef93f82 };
assign I59c80c7ec26f43308b1a646c47160568 = (I1223c21129382d41e4f38ef4bbe60c2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I08955fcfabffed0ad0c5e398e7872be1;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00191_00000_U (
.flogtanh_sel( I14e36e16df00adcd7dc1973d3852d2d9[flogtanh_SEL-1:0]),
.flogtanh( Ieb5fa20abbdb29a7f75021b7afafea31),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I99252b9918c30f2ba5611abc79e08fbb  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ieb5fa20abbdb29a7f75021b7afafea31 };
assign I8a954a331d36266465a0813d2e8b319b = (I14e36e16df00adcd7dc1973d3852d2d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I99252b9918c30f2ba5611abc79e08fbb;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00192_00000_U (
.flogtanh_sel( I0d05ae27b53fb6939e4c2f862a8d20b2[flogtanh_SEL-1:0]),
.flogtanh( I16a12326344aadf4226bd149424a53a8),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9cb632c1ab546359ef5a787a4bc3aaa6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I16a12326344aadf4226bd149424a53a8 };
assign Ib49e53ca8efd9564ee9572eb3089bb51 = (I0d05ae27b53fb6939e4c2f862a8d20b2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9cb632c1ab546359ef5a787a4bc3aaa6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00193_00000_U (
.flogtanh_sel( I97a6fcc08929c3b7d15e36d7706ed13d[flogtanh_SEL-1:0]),
.flogtanh( I07f36b533b48344c13dbb133739712f4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia4ee264b162c3ab4fec78ddb3a4fc6da  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I07f36b533b48344c13dbb133739712f4 };
assign Icbde2c6230e9cc67ef12031e38bb344f = (I97a6fcc08929c3b7d15e36d7706ed13d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia4ee264b162c3ab4fec78ddb3a4fc6da;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00194_00000_U (
.flogtanh_sel( I1f04e86bf27596718836d0a09adbe120[flogtanh_SEL-1:0]),
.flogtanh( I7a0072bf1e5fb0c4de85c6e4447878a4),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I116d3b804a2077edec9cf686b7cf5737  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I7a0072bf1e5fb0c4de85c6e4447878a4 };
assign I2e22e867f6f84a7807b82f64a147022e = (I1f04e86bf27596718836d0a09adbe120[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I116d3b804a2077edec9cf686b7cf5737;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00195_00000_U (
.flogtanh_sel( Ie40873cfd6d10a61a94a761becf588a8[flogtanh_SEL-1:0]),
.flogtanh( I320bafc5a1775d6933bcb9f2d2c84576),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5f89382f736f2688bc2c3696e0796002  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I320bafc5a1775d6933bcb9f2d2c84576 };
assign Id9704e1d8096cd28577c5c357d30b7a4 = (Ie40873cfd6d10a61a94a761becf588a8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5f89382f736f2688bc2c3696e0796002;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00196_00000_U (
.flogtanh_sel( I61960ed74fee948cc12bd1fd8384559a[flogtanh_SEL-1:0]),
.flogtanh( I5ec61756ff7237146f2d83f17eb5bb3a),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie139e712a1c886d4452735c1cd51af2e  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I5ec61756ff7237146f2d83f17eb5bb3a };
assign I4b8554cab486a4fc1e14884a6495016e = (I61960ed74fee948cc12bd1fd8384559a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie139e712a1c886d4452735c1cd51af2e;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00197_00000_U (
.flogtanh_sel( I8533a3ec4be4c49166184c94761eaebc[flogtanh_SEL-1:0]),
.flogtanh( I382008a17338641e68fa859ac2af1d20),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic3137e053b8e22028a8ccdeb9c573170  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I382008a17338641e68fa859ac2af1d20 };
assign Iaa235d085a5916a3b0814c3ed2a9026f = (I8533a3ec4be4c49166184c94761eaebc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic3137e053b8e22028a8ccdeb9c573170;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00198_00000_U (
.flogtanh_sel( I00be319b5bdb85ffaf3bb0eca0b348b6[flogtanh_SEL-1:0]),
.flogtanh( Ifd375ad8038ea2455c0e3b1463b83b7e),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8e15864be74893cd89bc56c0c2df858a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ifd375ad8038ea2455c0e3b1463b83b7e };
assign I5d86ce0b58c0b281d747116a9069ef33 = (I00be319b5bdb85ffaf3bb0eca0b348b6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8e15864be74893cd89bc56c0c2df858a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00199_00000_U (
.flogtanh_sel( Ie889c916b5af185b52ff5e2e3cc23045[flogtanh_SEL-1:0]),
.flogtanh( I0b75763235278d8eca6ca72fc97fb83c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I015b6b916b0b84ddbfded84bca8f849f  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I0b75763235278d8eca6ca72fc97fb83c };
assign Id20394136fb036435bb4680aac64581f = (Ie889c916b5af185b52ff5e2e3cc23045[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I015b6b916b0b84ddbfded84bca8f849f;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00200_00000_U (
.flogtanh_sel( I89697be6dcb2e7f972db498c1b1dea71[flogtanh_SEL-1:0]),
.flogtanh( I9bc4c3b77a9635bb77ad31527d961952),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7ee0d250f9a3166db6bd3f366059804a  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I9bc4c3b77a9635bb77ad31527d961952 };
assign I8a16afac6e470ca69634d7fe9656387a = (I89697be6dcb2e7f972db498c1b1dea71[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7ee0d250f9a3166db6bd3f366059804a;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00201_00000_U (
.flogtanh_sel( If13dfbfff7cd8e197bb44006a3db73bf[flogtanh_SEL-1:0]),
.flogtanh( Ief93f4a7eaaa1f43ea1788dc4629c093),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6fc4b3ab1858416a94ce844cd92277ce  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ief93f4a7eaaa1f43ea1788dc4629c093 };
assign Ic4e7f690bc050f1d1f84eae7ca193e1c = (If13dfbfff7cd8e197bb44006a3db73bf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6fc4b3ab1858416a94ce844cd92277ce;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00202_00000_U (
.flogtanh_sel( I87ed6c3e172c7a06bf6aefe7bf718d70[flogtanh_SEL-1:0]),
.flogtanh( I34b86fbc3949cb2083931ad8edd2444d),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9035dc3d53fc938d0927370681b669b3  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I34b86fbc3949cb2083931ad8edd2444d };
assign Ia60421aa427236540b4d0d08d52ff507 = (I87ed6c3e172c7a06bf6aefe7bf718d70[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9035dc3d53fc938d0927370681b669b3;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00203_00000_U (
.flogtanh_sel( I0db87adc849839fab3a4c9884d5a4882[flogtanh_SEL-1:0]),
.flogtanh( I560c163fb55aa4b56da25f96e9b8ef6c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I162c001a328c8bbc178403bc97725ed6  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, I560c163fb55aa4b56da25f96e9b8ef6c };
assign Icace650ee3865bd7bbddd2d9435c5561 = (I0db87adc849839fab3a4c9884d5a4882[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I162c001a328c8bbc178403bc97725ed6;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00204_00000_U (
.flogtanh_sel( I535e01a6c35fd7b455e4b79b1d4bb414[flogtanh_SEL-1:0]),
.flogtanh( Ib3c46d34c5bc3d2651147b3e764d9786),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5fac1be3058558fcba4ae7c095138a07  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ib3c46d34c5bc3d2651147b3e764d9786 };
assign I7d27d070b96b7810f667e1d1845342d3 = (I535e01a6c35fd7b455e4b79b1d4bb414[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5fac1be3058558fcba4ae7c095138a07;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00205_00000_U (
.flogtanh_sel( Ia2d1c752cc4b405adb97a815e90a7b96[flogtanh_SEL-1:0]),
.flogtanh( Ie5e2ba4fe22870afc81d6cfc708570be),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0e7ff238062811c5a3d3549bbf3bec52  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ie5e2ba4fe22870afc81d6cfc708570be };
assign Ida7ec09c913caa0e78a2c4cbaae517c8 = (Ia2d1c752cc4b405adb97a815e90a7b96[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0e7ff238062811c5a3d3549bbf3bec52;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00206_00000_U (
.flogtanh_sel( I9ac12eb3878f6fc7dc428fe5e7f35d97[flogtanh_SEL-1:0]),
.flogtanh( Ibf3bde181da4f960537516d6c0b2a72c),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie6509743f0bbe16d5f0aae9039db3d21  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ibf3bde181da4f960537516d6c0b2a72c };
assign Ic5eba898858be1f768841ead792d6d86 = (I9ac12eb3878f6fc7dc428fe5e7f35d97[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie6509743f0bbe16d5f0aae9039db3d21;


Ic3da32f100a43f826b89a492544e7812 flogtanh_00207_00000_U (
.flogtanh_sel( If46fa11dfadb0691eaaa0a40836e08d8[flogtanh_SEL-1:0]),
.flogtanh( Ia93f96aa0718f8755e9ebb8cc5d8f405),
.start_in(start_d3),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2b807f3aaa37eaddf34d61f95d436d48  = { {(MAX_SUM_WDTH_L-flogtanh_WDTH){1'b0}}, Ia93f96aa0718f8755e9ebb8cc5d8f405 };
assign I72197797a307c611fa8952533e63d7bf = (If46fa11dfadb0691eaaa0a40836e08d8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2b807f3aaa37eaddf34d61f95d436d48;





Ic9c2f173881d25f8976d723957809f51 fgallag_00000_00000_U (
.fgallag_sel( I97afe24956b7f87cd431f048202bab67[fgallag_SEL-1:0]),
.fgallag( fgallag_00000_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(start_d5),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00000_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00000_00000 };

assign fgallag_final_00000_00000 = (I97afe24956b7f87cd431f048202bab67[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00000_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00000_00001_U (
.fgallag_sel( I117235e3ac8e68e4c1ab34db1612aba0[fgallag_SEL-1:0]),
.fgallag( fgallag_00000_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00000_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00000_00001 };

assign fgallag_final_00000_00001 = (I117235e3ac8e68e4c1ab34db1612aba0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00000_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00000_00002_U (
.fgallag_sel( Ifd700cc9d18f99b63f1947f3ae631976[fgallag_SEL-1:0]),
.fgallag( fgallag_00000_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00000_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00000_00002 };

assign fgallag_final_00000_00002 = (Ifd700cc9d18f99b63f1947f3ae631976[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00000_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00000_00003_U (
.fgallag_sel( Ifffbe3d1007fb07a20d3b37902b3ec95[fgallag_SEL-1:0]),
.fgallag( fgallag_00000_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00000_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00000_00003 };

assign fgallag_final_00000_00003 = (Ifffbe3d1007fb07a20d3b37902b3ec95[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00000_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00000_00004_U (
.fgallag_sel( If5443777169422ea6e1e3f709b970e05[fgallag_SEL-1:0]),
.fgallag( fgallag_00000_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00000_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00000_00004 };

assign fgallag_final_00000_00004 = (If5443777169422ea6e1e3f709b970e05[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00000_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00000_00005_U (
.fgallag_sel( Ifaf9fc93e4609d818aa46751754c17f1[fgallag_SEL-1:0]),
.fgallag( fgallag_00000_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00000_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00000_00005 };

assign fgallag_final_00000_00005 = (Ifaf9fc93e4609d818aa46751754c17f1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00000_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00000_00006_U (
.fgallag_sel( I419caf964986c655df84d043badc37c9[fgallag_SEL-1:0]),
.fgallag( fgallag_00000_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00000_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00000_00006 };

assign fgallag_final_00000_00006 = (I419caf964986c655df84d043badc37c9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00000_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00000_00007_U (
.fgallag_sel( I3095214ac0e6c1323e75ee4ec85e6821[fgallag_SEL-1:0]),
.fgallag( fgallag_00000_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00000_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00000_00007 };

assign fgallag_final_00000_00007 = (I3095214ac0e6c1323e75ee4ec85e6821[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00000_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00001_00000_U (
.fgallag_sel( Ided9739bf63937933250a6d0c37535f9[fgallag_SEL-1:0]),
.fgallag( fgallag_00001_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00001_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00001_00000 };

assign fgallag_final_00001_00000 = (Ided9739bf63937933250a6d0c37535f9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00001_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00001_00001_U (
.fgallag_sel( Id0f139b9f3848b45554ac8429230eea2[fgallag_SEL-1:0]),
.fgallag( fgallag_00001_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00001_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00001_00001 };

assign fgallag_final_00001_00001 = (Id0f139b9f3848b45554ac8429230eea2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00001_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00001_00002_U (
.fgallag_sel( Id9feed58cf9565255abfd0bf7e3ec068[fgallag_SEL-1:0]),
.fgallag( fgallag_00001_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00001_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00001_00002 };

assign fgallag_final_00001_00002 = (Id9feed58cf9565255abfd0bf7e3ec068[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00001_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00001_00003_U (
.fgallag_sel( I30a3be3b5f6ad1880a917eb35659a1bf[fgallag_SEL-1:0]),
.fgallag( fgallag_00001_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00001_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00001_00003 };

assign fgallag_final_00001_00003 = (I30a3be3b5f6ad1880a917eb35659a1bf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00001_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00001_00004_U (
.fgallag_sel( Ie8148d9aa962a733eb65877b902a187d[fgallag_SEL-1:0]),
.fgallag( fgallag_00001_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00001_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00001_00004 };

assign fgallag_final_00001_00004 = (Ie8148d9aa962a733eb65877b902a187d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00001_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00001_00005_U (
.fgallag_sel( I69e98cf3e679183aef6005bb582b18dc[fgallag_SEL-1:0]),
.fgallag( fgallag_00001_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00001_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00001_00005 };

assign fgallag_final_00001_00005 = (I69e98cf3e679183aef6005bb582b18dc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00001_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00001_00006_U (
.fgallag_sel( I7f42a504fc61c9548acebdd8b1858eaa[fgallag_SEL-1:0]),
.fgallag( fgallag_00001_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00001_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00001_00006 };

assign fgallag_final_00001_00006 = (I7f42a504fc61c9548acebdd8b1858eaa[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00001_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00001_00007_U (
.fgallag_sel( I08b1b4639b5a9ca509b943b977f6d4bb[fgallag_SEL-1:0]),
.fgallag( fgallag_00001_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00001_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00001_00007 };

assign fgallag_final_00001_00007 = (I08b1b4639b5a9ca509b943b977f6d4bb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00001_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00002_00000_U (
.fgallag_sel( I8d7296627d886566783e79c01b9fa423[fgallag_SEL-1:0]),
.fgallag( fgallag_00002_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00002_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00002_00000 };

assign fgallag_final_00002_00000 = (I8d7296627d886566783e79c01b9fa423[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00002_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00002_00001_U (
.fgallag_sel( I4fc4c97229a8b1f631a3b505941159e4[fgallag_SEL-1:0]),
.fgallag( fgallag_00002_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00002_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00002_00001 };

assign fgallag_final_00002_00001 = (I4fc4c97229a8b1f631a3b505941159e4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00002_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00002_00002_U (
.fgallag_sel( Ib9b16bf51891c328dba2699eb9bcef95[fgallag_SEL-1:0]),
.fgallag( fgallag_00002_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00002_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00002_00002 };

assign fgallag_final_00002_00002 = (Ib9b16bf51891c328dba2699eb9bcef95[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00002_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00002_00003_U (
.fgallag_sel( I6c30501ec81fce286817788d614a7824[fgallag_SEL-1:0]),
.fgallag( fgallag_00002_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00002_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00002_00003 };

assign fgallag_final_00002_00003 = (I6c30501ec81fce286817788d614a7824[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00002_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00002_00004_U (
.fgallag_sel( Ia4d4f37baec48121a88808075dd655ef[fgallag_SEL-1:0]),
.fgallag( fgallag_00002_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00002_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00002_00004 };

assign fgallag_final_00002_00004 = (Ia4d4f37baec48121a88808075dd655ef[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00002_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00002_00005_U (
.fgallag_sel( I385495ea2bf6442a95ab7561456254ac[fgallag_SEL-1:0]),
.fgallag( fgallag_00002_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00002_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00002_00005 };

assign fgallag_final_00002_00005 = (I385495ea2bf6442a95ab7561456254ac[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00002_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00002_00006_U (
.fgallag_sel( I5128e03d383c226befa6f7422f3a6f04[fgallag_SEL-1:0]),
.fgallag( fgallag_00002_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00002_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00002_00006 };

assign fgallag_final_00002_00006 = (I5128e03d383c226befa6f7422f3a6f04[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00002_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00002_00007_U (
.fgallag_sel( Ib208908bab4c20713cd17e20139c8db3[fgallag_SEL-1:0]),
.fgallag( fgallag_00002_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00002_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00002_00007 };

assign fgallag_final_00002_00007 = (Ib208908bab4c20713cd17e20139c8db3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00002_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00003_00000_U (
.fgallag_sel( Id939992b99a11c09f4688c10ca1a34d1[fgallag_SEL-1:0]),
.fgallag( fgallag_00003_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00003_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00003_00000 };

assign fgallag_final_00003_00000 = (Id939992b99a11c09f4688c10ca1a34d1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00003_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00003_00001_U (
.fgallag_sel( I823453ccb90d5b2b2d9dfc6e8358224d[fgallag_SEL-1:0]),
.fgallag( fgallag_00003_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00003_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00003_00001 };

assign fgallag_final_00003_00001 = (I823453ccb90d5b2b2d9dfc6e8358224d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00003_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00003_00002_U (
.fgallag_sel( I279c5c00b92eb1b872b5afa168b0306e[fgallag_SEL-1:0]),
.fgallag( fgallag_00003_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00003_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00003_00002 };

assign fgallag_final_00003_00002 = (I279c5c00b92eb1b872b5afa168b0306e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00003_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00003_00003_U (
.fgallag_sel( I66f25b1c3c0eb226295179adcca2c3d2[fgallag_SEL-1:0]),
.fgallag( fgallag_00003_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00003_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00003_00003 };

assign fgallag_final_00003_00003 = (I66f25b1c3c0eb226295179adcca2c3d2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00003_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00003_00004_U (
.fgallag_sel( I3068627e91b667d14cd3e55a9371931a[fgallag_SEL-1:0]),
.fgallag( fgallag_00003_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00003_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00003_00004 };

assign fgallag_final_00003_00004 = (I3068627e91b667d14cd3e55a9371931a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00003_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00003_00005_U (
.fgallag_sel( I44c4e0a2d8a7289f8660b81a9ecfa19b[fgallag_SEL-1:0]),
.fgallag( fgallag_00003_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00003_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00003_00005 };

assign fgallag_final_00003_00005 = (I44c4e0a2d8a7289f8660b81a9ecfa19b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00003_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00003_00006_U (
.fgallag_sel( Ibe868e258dc87f0dd1460ba6b8354671[fgallag_SEL-1:0]),
.fgallag( fgallag_00003_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00003_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00003_00006 };

assign fgallag_final_00003_00006 = (Ibe868e258dc87f0dd1460ba6b8354671[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00003_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00003_00007_U (
.fgallag_sel( Idc3083c3021200345e3edd35a9d4725a[fgallag_SEL-1:0]),
.fgallag( fgallag_00003_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00003_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00003_00007 };

assign fgallag_final_00003_00007 = (Idc3083c3021200345e3edd35a9d4725a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00003_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00004_00000_U (
.fgallag_sel( I320d4f19a5b18c23ff407508d47caa77[fgallag_SEL-1:0]),
.fgallag( fgallag_00004_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00004_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00004_00000 };

assign fgallag_final_00004_00000 = (I320d4f19a5b18c23ff407508d47caa77[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00004_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00004_00001_U (
.fgallag_sel( I16becf3c92615d98d5ec51ee9641cc0a[fgallag_SEL-1:0]),
.fgallag( fgallag_00004_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00004_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00004_00001 };

assign fgallag_final_00004_00001 = (I16becf3c92615d98d5ec51ee9641cc0a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00004_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00004_00002_U (
.fgallag_sel( Ifbfacc3b3a0128119943bcbf80176612[fgallag_SEL-1:0]),
.fgallag( fgallag_00004_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00004_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00004_00002 };

assign fgallag_final_00004_00002 = (Ifbfacc3b3a0128119943bcbf80176612[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00004_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00004_00003_U (
.fgallag_sel( I6b4f670c9e8e25984e8891f2440322ab[fgallag_SEL-1:0]),
.fgallag( fgallag_00004_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00004_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00004_00003 };

assign fgallag_final_00004_00003 = (I6b4f670c9e8e25984e8891f2440322ab[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00004_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00004_00004_U (
.fgallag_sel( I19bf0990a30c72421f231772b8627e8e[fgallag_SEL-1:0]),
.fgallag( fgallag_00004_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00004_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00004_00004 };

assign fgallag_final_00004_00004 = (I19bf0990a30c72421f231772b8627e8e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00004_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00004_00005_U (
.fgallag_sel( I3ec3eb096ebe3ee8a47e1cba6487b997[fgallag_SEL-1:0]),
.fgallag( fgallag_00004_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00004_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00004_00005 };

assign fgallag_final_00004_00005 = (I3ec3eb096ebe3ee8a47e1cba6487b997[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00004_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00004_00006_U (
.fgallag_sel( I7379ef16405c461ac44b66c4315df831[fgallag_SEL-1:0]),
.fgallag( fgallag_00004_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00004_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00004_00006 };

assign fgallag_final_00004_00006 = (I7379ef16405c461ac44b66c4315df831[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00004_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00004_00007_U (
.fgallag_sel( I79db45b23d21d533a1f9a6e8f94d403d[fgallag_SEL-1:0]),
.fgallag( fgallag_00004_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00004_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00004_00007 };

assign fgallag_final_00004_00007 = (I79db45b23d21d533a1f9a6e8f94d403d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00004_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00004_00008_U (
.fgallag_sel( I0979534730cc2b53547d413dbb6b75f4[fgallag_SEL-1:0]),
.fgallag( fgallag_00004_00008 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00004_00008 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00004_00008 };

assign fgallag_final_00004_00008 = (I0979534730cc2b53547d413dbb6b75f4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00004_00008 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00004_00009_U (
.fgallag_sel( I5aa2f9c0667d1a6e871efbd4d2bad3a8[fgallag_SEL-1:0]),
.fgallag( fgallag_00004_00009 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00004_00009 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00004_00009 };

assign fgallag_final_00004_00009 = (I5aa2f9c0667d1a6e871efbd4d2bad3a8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00004_00009 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00005_00000_U (
.fgallag_sel( Iadb28dc990ccf2dd3099544de16b8f16[fgallag_SEL-1:0]),
.fgallag( fgallag_00005_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00005_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00005_00000 };

assign fgallag_final_00005_00000 = (Iadb28dc990ccf2dd3099544de16b8f16[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00005_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00005_00001_U (
.fgallag_sel( I1f71aebf698788d6ada66891e9ea756f[fgallag_SEL-1:0]),
.fgallag( fgallag_00005_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00005_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00005_00001 };

assign fgallag_final_00005_00001 = (I1f71aebf698788d6ada66891e9ea756f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00005_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00005_00002_U (
.fgallag_sel( Ib234e9cf7e7616a1ebc6ab99df2a7ccb[fgallag_SEL-1:0]),
.fgallag( fgallag_00005_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00005_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00005_00002 };

assign fgallag_final_00005_00002 = (Ib234e9cf7e7616a1ebc6ab99df2a7ccb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00005_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00005_00003_U (
.fgallag_sel( I297d1edcc583ea4d69da780150f0620c[fgallag_SEL-1:0]),
.fgallag( fgallag_00005_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00005_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00005_00003 };

assign fgallag_final_00005_00003 = (I297d1edcc583ea4d69da780150f0620c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00005_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00005_00004_U (
.fgallag_sel( Ib0a717cbb4fe38a3fc85520ca0826fd9[fgallag_SEL-1:0]),
.fgallag( fgallag_00005_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00005_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00005_00004 };

assign fgallag_final_00005_00004 = (Ib0a717cbb4fe38a3fc85520ca0826fd9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00005_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00005_00005_U (
.fgallag_sel( I037ecd5945b1f1280b4469d73fe1c7ff[fgallag_SEL-1:0]),
.fgallag( fgallag_00005_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00005_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00005_00005 };

assign fgallag_final_00005_00005 = (I037ecd5945b1f1280b4469d73fe1c7ff[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00005_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00005_00006_U (
.fgallag_sel( I367ff6b11b884e02a3065fc7fe811e15[fgallag_SEL-1:0]),
.fgallag( fgallag_00005_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00005_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00005_00006 };

assign fgallag_final_00005_00006 = (I367ff6b11b884e02a3065fc7fe811e15[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00005_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00005_00007_U (
.fgallag_sel( I6fab19692b512166fe9c74b5e987788d[fgallag_SEL-1:0]),
.fgallag( fgallag_00005_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00005_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00005_00007 };

assign fgallag_final_00005_00007 = (I6fab19692b512166fe9c74b5e987788d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00005_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00005_00008_U (
.fgallag_sel( I04dd73af505f618ccdb209b3cf97ceec[fgallag_SEL-1:0]),
.fgallag( fgallag_00005_00008 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00005_00008 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00005_00008 };

assign fgallag_final_00005_00008 = (I04dd73af505f618ccdb209b3cf97ceec[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00005_00008 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00005_00009_U (
.fgallag_sel( If8c559905d4120488d431719c4e8ce24[fgallag_SEL-1:0]),
.fgallag( fgallag_00005_00009 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00005_00009 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00005_00009 };

assign fgallag_final_00005_00009 = (If8c559905d4120488d431719c4e8ce24[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00005_00009 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00006_00000_U (
.fgallag_sel( I20ed4f6f14e20ce3f0e106d1b7782fcd[fgallag_SEL-1:0]),
.fgallag( fgallag_00006_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00006_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00006_00000 };

assign fgallag_final_00006_00000 = (I20ed4f6f14e20ce3f0e106d1b7782fcd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00006_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00006_00001_U (
.fgallag_sel( Ib10626ffa126188c5bf1fc8399107b26[fgallag_SEL-1:0]),
.fgallag( fgallag_00006_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00006_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00006_00001 };

assign fgallag_final_00006_00001 = (Ib10626ffa126188c5bf1fc8399107b26[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00006_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00006_00002_U (
.fgallag_sel( I29007c52357ac7afbda39d72a5bb60af[fgallag_SEL-1:0]),
.fgallag( fgallag_00006_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00006_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00006_00002 };

assign fgallag_final_00006_00002 = (I29007c52357ac7afbda39d72a5bb60af[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00006_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00006_00003_U (
.fgallag_sel( I66d367c046611f145e607a90911cf499[fgallag_SEL-1:0]),
.fgallag( fgallag_00006_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00006_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00006_00003 };

assign fgallag_final_00006_00003 = (I66d367c046611f145e607a90911cf499[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00006_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00006_00004_U (
.fgallag_sel( I9c4c2556f6170a8df61d909855a846ed[fgallag_SEL-1:0]),
.fgallag( fgallag_00006_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00006_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00006_00004 };

assign fgallag_final_00006_00004 = (I9c4c2556f6170a8df61d909855a846ed[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00006_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00006_00005_U (
.fgallag_sel( I6fadc3e8d995bb4317bf7b4377c3c2c5[fgallag_SEL-1:0]),
.fgallag( fgallag_00006_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00006_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00006_00005 };

assign fgallag_final_00006_00005 = (I6fadc3e8d995bb4317bf7b4377c3c2c5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00006_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00006_00006_U (
.fgallag_sel( I99b20e911c189e0616f02376ab736e91[fgallag_SEL-1:0]),
.fgallag( fgallag_00006_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00006_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00006_00006 };

assign fgallag_final_00006_00006 = (I99b20e911c189e0616f02376ab736e91[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00006_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00006_00007_U (
.fgallag_sel( I5793c12f5dbdd8245dbb202d550ca960[fgallag_SEL-1:0]),
.fgallag( fgallag_00006_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00006_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00006_00007 };

assign fgallag_final_00006_00007 = (I5793c12f5dbdd8245dbb202d550ca960[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00006_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00006_00008_U (
.fgallag_sel( Id0660e9637cad1ce1a73d37188060154[fgallag_SEL-1:0]),
.fgallag( fgallag_00006_00008 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00006_00008 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00006_00008 };

assign fgallag_final_00006_00008 = (Id0660e9637cad1ce1a73d37188060154[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00006_00008 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00006_00009_U (
.fgallag_sel( If5a7af7ca023e1393526e888f4220a44[fgallag_SEL-1:0]),
.fgallag( fgallag_00006_00009 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00006_00009 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00006_00009 };

assign fgallag_final_00006_00009 = (If5a7af7ca023e1393526e888f4220a44[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00006_00009 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00007_00000_U (
.fgallag_sel( Id043eb50634e803e53adc1168379a5d0[fgallag_SEL-1:0]),
.fgallag( fgallag_00007_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00007_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00007_00000 };

assign fgallag_final_00007_00000 = (Id043eb50634e803e53adc1168379a5d0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00007_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00007_00001_U (
.fgallag_sel( I1f866dd0b129267550aea1a267d9c91e[fgallag_SEL-1:0]),
.fgallag( fgallag_00007_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00007_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00007_00001 };

assign fgallag_final_00007_00001 = (I1f866dd0b129267550aea1a267d9c91e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00007_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00007_00002_U (
.fgallag_sel( I8c4da05c08210fe33139c3d3e5d75d58[fgallag_SEL-1:0]),
.fgallag( fgallag_00007_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00007_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00007_00002 };

assign fgallag_final_00007_00002 = (I8c4da05c08210fe33139c3d3e5d75d58[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00007_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00007_00003_U (
.fgallag_sel( Ib41f7b823681fdd084b6d8436a407aa8[fgallag_SEL-1:0]),
.fgallag( fgallag_00007_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00007_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00007_00003 };

assign fgallag_final_00007_00003 = (Ib41f7b823681fdd084b6d8436a407aa8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00007_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00007_00004_U (
.fgallag_sel( Ic5b50a785b7acac7e3be4095aa92e50a[fgallag_SEL-1:0]),
.fgallag( fgallag_00007_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00007_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00007_00004 };

assign fgallag_final_00007_00004 = (Ic5b50a785b7acac7e3be4095aa92e50a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00007_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00007_00005_U (
.fgallag_sel( I3ffbe03796b66d00d47fd918be60ab89[fgallag_SEL-1:0]),
.fgallag( fgallag_00007_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00007_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00007_00005 };

assign fgallag_final_00007_00005 = (I3ffbe03796b66d00d47fd918be60ab89[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00007_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00007_00006_U (
.fgallag_sel( Ifc92a916da938ef6164db250be635f88[fgallag_SEL-1:0]),
.fgallag( fgallag_00007_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00007_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00007_00006 };

assign fgallag_final_00007_00006 = (Ifc92a916da938ef6164db250be635f88[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00007_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00007_00007_U (
.fgallag_sel( I8ccd42508ce7d5bd897c2cf0c54caeb3[fgallag_SEL-1:0]),
.fgallag( fgallag_00007_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00007_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00007_00007 };

assign fgallag_final_00007_00007 = (I8ccd42508ce7d5bd897c2cf0c54caeb3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00007_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00007_00008_U (
.fgallag_sel( I4920e7e82749cc036b58a7cd0a03e327[fgallag_SEL-1:0]),
.fgallag( fgallag_00007_00008 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00007_00008 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00007_00008 };

assign fgallag_final_00007_00008 = (I4920e7e82749cc036b58a7cd0a03e327[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00007_00008 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00007_00009_U (
.fgallag_sel( Ie1040b2aa91f272e4449c4b5f9f8f575[fgallag_SEL-1:0]),
.fgallag( fgallag_00007_00009 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00007_00009 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00007_00009 };

assign fgallag_final_00007_00009 = (Ie1040b2aa91f272e4449c4b5f9f8f575[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00007_00009 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00008_00000_U (
.fgallag_sel( I65968fb0f63d52ad96cd8fa270126a1b[fgallag_SEL-1:0]),
.fgallag( fgallag_00008_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00008_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00008_00000 };

assign fgallag_final_00008_00000 = (I65968fb0f63d52ad96cd8fa270126a1b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00008_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00008_00001_U (
.fgallag_sel( I839ac8ee59f51d4c3de92ba5cb26e788[fgallag_SEL-1:0]),
.fgallag( fgallag_00008_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00008_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00008_00001 };

assign fgallag_final_00008_00001 = (I839ac8ee59f51d4c3de92ba5cb26e788[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00008_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00008_00002_U (
.fgallag_sel( I33cd95f1919318a0f3df5df7310d64c6[fgallag_SEL-1:0]),
.fgallag( fgallag_00008_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00008_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00008_00002 };

assign fgallag_final_00008_00002 = (I33cd95f1919318a0f3df5df7310d64c6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00008_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00008_00003_U (
.fgallag_sel( I4933e8d16fba26cd797b25a9ac2a2de8[fgallag_SEL-1:0]),
.fgallag( fgallag_00008_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00008_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00008_00003 };

assign fgallag_final_00008_00003 = (I4933e8d16fba26cd797b25a9ac2a2de8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00008_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00008_00004_U (
.fgallag_sel( I218f7578eb748e31d0002052f30c5842[fgallag_SEL-1:0]),
.fgallag( fgallag_00008_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00008_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00008_00004 };

assign fgallag_final_00008_00004 = (I218f7578eb748e31d0002052f30c5842[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00008_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00008_00005_U (
.fgallag_sel( I2a808d1c42ad758ae3baaaee8129dfb2[fgallag_SEL-1:0]),
.fgallag( fgallag_00008_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00008_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00008_00005 };

assign fgallag_final_00008_00005 = (I2a808d1c42ad758ae3baaaee8129dfb2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00008_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00008_00006_U (
.fgallag_sel( I4e851fd3c114af87f5e8c68c02594e3a[fgallag_SEL-1:0]),
.fgallag( fgallag_00008_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00008_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00008_00006 };

assign fgallag_final_00008_00006 = (I4e851fd3c114af87f5e8c68c02594e3a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00008_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00008_00007_U (
.fgallag_sel( I0da40f88adc46e90f616acdcdb8e0e2c[fgallag_SEL-1:0]),
.fgallag( fgallag_00008_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00008_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00008_00007 };

assign fgallag_final_00008_00007 = (I0da40f88adc46e90f616acdcdb8e0e2c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00008_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00009_00000_U (
.fgallag_sel( I0dee7767e472a5fd71250ae6c57cc8b5[fgallag_SEL-1:0]),
.fgallag( fgallag_00009_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00009_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00009_00000 };

assign fgallag_final_00009_00000 = (I0dee7767e472a5fd71250ae6c57cc8b5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00009_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00009_00001_U (
.fgallag_sel( I9f40be7552b3dd625e5bce0befc5a548[fgallag_SEL-1:0]),
.fgallag( fgallag_00009_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00009_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00009_00001 };

assign fgallag_final_00009_00001 = (I9f40be7552b3dd625e5bce0befc5a548[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00009_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00009_00002_U (
.fgallag_sel( I8fdf98ffd757c8845ed6ffa4ddd1a16b[fgallag_SEL-1:0]),
.fgallag( fgallag_00009_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00009_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00009_00002 };

assign fgallag_final_00009_00002 = (I8fdf98ffd757c8845ed6ffa4ddd1a16b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00009_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00009_00003_U (
.fgallag_sel( I8103b777314a4fa471e0898fde9cde08[fgallag_SEL-1:0]),
.fgallag( fgallag_00009_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00009_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00009_00003 };

assign fgallag_final_00009_00003 = (I8103b777314a4fa471e0898fde9cde08[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00009_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00009_00004_U (
.fgallag_sel( If6c3ee8e0d7dea58043d5be0f4630873[fgallag_SEL-1:0]),
.fgallag( fgallag_00009_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00009_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00009_00004 };

assign fgallag_final_00009_00004 = (If6c3ee8e0d7dea58043d5be0f4630873[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00009_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00009_00005_U (
.fgallag_sel( I711a5171f591f472cdbfc9a0f5e1aa17[fgallag_SEL-1:0]),
.fgallag( fgallag_00009_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00009_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00009_00005 };

assign fgallag_final_00009_00005 = (I711a5171f591f472cdbfc9a0f5e1aa17[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00009_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00009_00006_U (
.fgallag_sel( Ic30bc38184dfbbd694af52640692709d[fgallag_SEL-1:0]),
.fgallag( fgallag_00009_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00009_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00009_00006 };

assign fgallag_final_00009_00006 = (Ic30bc38184dfbbd694af52640692709d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00009_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00009_00007_U (
.fgallag_sel( I422f6fd1d273a3834d04b04ab8e2812d[fgallag_SEL-1:0]),
.fgallag( fgallag_00009_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00009_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00009_00007 };

assign fgallag_final_00009_00007 = (I422f6fd1d273a3834d04b04ab8e2812d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00009_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00010_00000_U (
.fgallag_sel( Ia0fdc60b90ad18b6585ec1ad4e89e80b[fgallag_SEL-1:0]),
.fgallag( fgallag_00010_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00010_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00010_00000 };

assign fgallag_final_00010_00000 = (Ia0fdc60b90ad18b6585ec1ad4e89e80b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00010_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00010_00001_U (
.fgallag_sel( I7809fe7a30d041a7e569ffe890242df8[fgallag_SEL-1:0]),
.fgallag( fgallag_00010_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00010_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00010_00001 };

assign fgallag_final_00010_00001 = (I7809fe7a30d041a7e569ffe890242df8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00010_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00010_00002_U (
.fgallag_sel( I672b14ec1b3c4797545f266727505a85[fgallag_SEL-1:0]),
.fgallag( fgallag_00010_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00010_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00010_00002 };

assign fgallag_final_00010_00002 = (I672b14ec1b3c4797545f266727505a85[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00010_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00010_00003_U (
.fgallag_sel( If9620d20ebaae6245a2c386d9bf5fdb1[fgallag_SEL-1:0]),
.fgallag( fgallag_00010_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00010_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00010_00003 };

assign fgallag_final_00010_00003 = (If9620d20ebaae6245a2c386d9bf5fdb1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00010_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00010_00004_U (
.fgallag_sel( Ic74e22bffd88f32eefe499cde0fafa8a[fgallag_SEL-1:0]),
.fgallag( fgallag_00010_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00010_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00010_00004 };

assign fgallag_final_00010_00004 = (Ic74e22bffd88f32eefe499cde0fafa8a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00010_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00010_00005_U (
.fgallag_sel( I76d38ce67387bd76ab45c9cba7d18b31[fgallag_SEL-1:0]),
.fgallag( fgallag_00010_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00010_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00010_00005 };

assign fgallag_final_00010_00005 = (I76d38ce67387bd76ab45c9cba7d18b31[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00010_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00010_00006_U (
.fgallag_sel( I44413c6f6f6493f8a86abf6eb32604f6[fgallag_SEL-1:0]),
.fgallag( fgallag_00010_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00010_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00010_00006 };

assign fgallag_final_00010_00006 = (I44413c6f6f6493f8a86abf6eb32604f6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00010_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00010_00007_U (
.fgallag_sel( I67f632fca617fe06565ddcaaee8fa8b8[fgallag_SEL-1:0]),
.fgallag( fgallag_00010_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00010_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00010_00007 };

assign fgallag_final_00010_00007 = (I67f632fca617fe06565ddcaaee8fa8b8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00010_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00011_00000_U (
.fgallag_sel( I3fd38a71ce6aa3db1d7a5a9f8a991e12[fgallag_SEL-1:0]),
.fgallag( fgallag_00011_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00011_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00011_00000 };

assign fgallag_final_00011_00000 = (I3fd38a71ce6aa3db1d7a5a9f8a991e12[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00011_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00011_00001_U (
.fgallag_sel( I63e5718bf7d8771ef90b91be73d73264[fgallag_SEL-1:0]),
.fgallag( fgallag_00011_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00011_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00011_00001 };

assign fgallag_final_00011_00001 = (I63e5718bf7d8771ef90b91be73d73264[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00011_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00011_00002_U (
.fgallag_sel( Ie385e1aeb2b0dcf6d2454be3d7708b27[fgallag_SEL-1:0]),
.fgallag( fgallag_00011_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00011_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00011_00002 };

assign fgallag_final_00011_00002 = (Ie385e1aeb2b0dcf6d2454be3d7708b27[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00011_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00011_00003_U (
.fgallag_sel( Ib2d1b7e105b25b492b45da72536d7578[fgallag_SEL-1:0]),
.fgallag( fgallag_00011_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00011_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00011_00003 };

assign fgallag_final_00011_00003 = (Ib2d1b7e105b25b492b45da72536d7578[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00011_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00011_00004_U (
.fgallag_sel( I588abf5ef4c583f0fec422736a0ce6a0[fgallag_SEL-1:0]),
.fgallag( fgallag_00011_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00011_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00011_00004 };

assign fgallag_final_00011_00004 = (I588abf5ef4c583f0fec422736a0ce6a0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00011_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00011_00005_U (
.fgallag_sel( I58bb95c56c7be17c263a2161210d7d8d[fgallag_SEL-1:0]),
.fgallag( fgallag_00011_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00011_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00011_00005 };

assign fgallag_final_00011_00005 = (I58bb95c56c7be17c263a2161210d7d8d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00011_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00011_00006_U (
.fgallag_sel( Ifaf0e1f21b3bd7393c475b5126540a72[fgallag_SEL-1:0]),
.fgallag( fgallag_00011_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00011_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00011_00006 };

assign fgallag_final_00011_00006 = (Ifaf0e1f21b3bd7393c475b5126540a72[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00011_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00011_00007_U (
.fgallag_sel( I7027db9e0450724a6d417d708f1043f2[fgallag_SEL-1:0]),
.fgallag( fgallag_00011_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00011_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00011_00007 };

assign fgallag_final_00011_00007 = (I7027db9e0450724a6d417d708f1043f2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00011_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00012_00000_U (
.fgallag_sel( Iebcb7206d8860b5094459c5d10b4efed[fgallag_SEL-1:0]),
.fgallag( fgallag_00012_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00012_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00012_00000 };

assign fgallag_final_00012_00000 = (Iebcb7206d8860b5094459c5d10b4efed[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00012_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00012_00001_U (
.fgallag_sel( I6bbf2b47a7dc50e66a3d8d258d6e31fb[fgallag_SEL-1:0]),
.fgallag( fgallag_00012_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00012_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00012_00001 };

assign fgallag_final_00012_00001 = (I6bbf2b47a7dc50e66a3d8d258d6e31fb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00012_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00012_00002_U (
.fgallag_sel( I8459abaa907f5afcd11884b1ec8c06c5[fgallag_SEL-1:0]),
.fgallag( fgallag_00012_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00012_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00012_00002 };

assign fgallag_final_00012_00002 = (I8459abaa907f5afcd11884b1ec8c06c5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00012_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00012_00003_U (
.fgallag_sel( Ia16ae2f6ef5000d47b6b84ed058252aa[fgallag_SEL-1:0]),
.fgallag( fgallag_00012_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00012_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00012_00003 };

assign fgallag_final_00012_00003 = (Ia16ae2f6ef5000d47b6b84ed058252aa[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00012_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00012_00004_U (
.fgallag_sel( Ica32690dbc9ea110fefdce92260b125c[fgallag_SEL-1:0]),
.fgallag( fgallag_00012_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00012_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00012_00004 };

assign fgallag_final_00012_00004 = (Ica32690dbc9ea110fefdce92260b125c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00012_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00012_00005_U (
.fgallag_sel( Ic431d9383cce30b1889c92e2be4cb9d0[fgallag_SEL-1:0]),
.fgallag( fgallag_00012_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00012_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00012_00005 };

assign fgallag_final_00012_00005 = (Ic431d9383cce30b1889c92e2be4cb9d0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00012_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00012_00006_U (
.fgallag_sel( Ib9cca4c0e58373c26d5fd9f51f793898[fgallag_SEL-1:0]),
.fgallag( fgallag_00012_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00012_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00012_00006 };

assign fgallag_final_00012_00006 = (Ib9cca4c0e58373c26d5fd9f51f793898[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00012_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00012_00007_U (
.fgallag_sel( I99bf0bc8ac20832b3724b2753f6ca449[fgallag_SEL-1:0]),
.fgallag( fgallag_00012_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00012_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00012_00007 };

assign fgallag_final_00012_00007 = (I99bf0bc8ac20832b3724b2753f6ca449[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00012_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00012_00008_U (
.fgallag_sel( Ie701008f3c60c51ed72c5f964a8fc36e[fgallag_SEL-1:0]),
.fgallag( fgallag_00012_00008 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00012_00008 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00012_00008 };

assign fgallag_final_00012_00008 = (Ie701008f3c60c51ed72c5f964a8fc36e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00012_00008 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00012_00009_U (
.fgallag_sel( I3e2d78f8307a1787f8b2eccba94c7557[fgallag_SEL-1:0]),
.fgallag( fgallag_00012_00009 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00012_00009 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00012_00009 };

assign fgallag_final_00012_00009 = (I3e2d78f8307a1787f8b2eccba94c7557[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00012_00009 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00013_00000_U (
.fgallag_sel( Ic1b4444ab0df9745d29bf893d9b83168[fgallag_SEL-1:0]),
.fgallag( fgallag_00013_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00013_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00013_00000 };

assign fgallag_final_00013_00000 = (Ic1b4444ab0df9745d29bf893d9b83168[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00013_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00013_00001_U (
.fgallag_sel( I5f52dbf600656a8f5dc6b6b8a45ccebe[fgallag_SEL-1:0]),
.fgallag( fgallag_00013_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00013_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00013_00001 };

assign fgallag_final_00013_00001 = (I5f52dbf600656a8f5dc6b6b8a45ccebe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00013_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00013_00002_U (
.fgallag_sel( I7f307af79f45ad4b9511e3961c917078[fgallag_SEL-1:0]),
.fgallag( fgallag_00013_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00013_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00013_00002 };

assign fgallag_final_00013_00002 = (I7f307af79f45ad4b9511e3961c917078[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00013_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00013_00003_U (
.fgallag_sel( Ie17a5be2a16d2efb98c976d7ee882535[fgallag_SEL-1:0]),
.fgallag( fgallag_00013_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00013_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00013_00003 };

assign fgallag_final_00013_00003 = (Ie17a5be2a16d2efb98c976d7ee882535[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00013_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00013_00004_U (
.fgallag_sel( I5f19d2adff2f34a4bebe03f929a09c49[fgallag_SEL-1:0]),
.fgallag( fgallag_00013_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00013_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00013_00004 };

assign fgallag_final_00013_00004 = (I5f19d2adff2f34a4bebe03f929a09c49[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00013_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00013_00005_U (
.fgallag_sel( I3cd69aeed9e869a2096d6dced5c209a0[fgallag_SEL-1:0]),
.fgallag( fgallag_00013_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00013_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00013_00005 };

assign fgallag_final_00013_00005 = (I3cd69aeed9e869a2096d6dced5c209a0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00013_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00013_00006_U (
.fgallag_sel( I359b6a22c9568a13b81670c741281393[fgallag_SEL-1:0]),
.fgallag( fgallag_00013_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00013_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00013_00006 };

assign fgallag_final_00013_00006 = (I359b6a22c9568a13b81670c741281393[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00013_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00013_00007_U (
.fgallag_sel( I24ba99614df383c38bbac50ae8b4487e[fgallag_SEL-1:0]),
.fgallag( fgallag_00013_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00013_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00013_00007 };

assign fgallag_final_00013_00007 = (I24ba99614df383c38bbac50ae8b4487e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00013_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00013_00008_U (
.fgallag_sel( I7498bee46de6b1c946ce95fdcc89f6e5[fgallag_SEL-1:0]),
.fgallag( fgallag_00013_00008 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00013_00008 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00013_00008 };

assign fgallag_final_00013_00008 = (I7498bee46de6b1c946ce95fdcc89f6e5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00013_00008 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00013_00009_U (
.fgallag_sel( I0f644f42cabf871b71e5a82871bc7b5d[fgallag_SEL-1:0]),
.fgallag( fgallag_00013_00009 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00013_00009 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00013_00009 };

assign fgallag_final_00013_00009 = (I0f644f42cabf871b71e5a82871bc7b5d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00013_00009 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00014_00000_U (
.fgallag_sel( I71f9e059726a6cac8bdf0efcc0eadd2b[fgallag_SEL-1:0]),
.fgallag( fgallag_00014_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00014_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00014_00000 };

assign fgallag_final_00014_00000 = (I71f9e059726a6cac8bdf0efcc0eadd2b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00014_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00014_00001_U (
.fgallag_sel( I0c9b2c1da30bfab514bbb556ae7bd4c4[fgallag_SEL-1:0]),
.fgallag( fgallag_00014_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00014_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00014_00001 };

assign fgallag_final_00014_00001 = (I0c9b2c1da30bfab514bbb556ae7bd4c4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00014_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00014_00002_U (
.fgallag_sel( I7918b2e37e96aee94fbccca7e0f75fc4[fgallag_SEL-1:0]),
.fgallag( fgallag_00014_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00014_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00014_00002 };

assign fgallag_final_00014_00002 = (I7918b2e37e96aee94fbccca7e0f75fc4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00014_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00014_00003_U (
.fgallag_sel( I76eebd77eb77e0abcbc727d2c511370a[fgallag_SEL-1:0]),
.fgallag( fgallag_00014_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00014_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00014_00003 };

assign fgallag_final_00014_00003 = (I76eebd77eb77e0abcbc727d2c511370a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00014_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00014_00004_U (
.fgallag_sel( Ibb2288e62110bae5b2d3fe901974e5c7[fgallag_SEL-1:0]),
.fgallag( fgallag_00014_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00014_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00014_00004 };

assign fgallag_final_00014_00004 = (Ibb2288e62110bae5b2d3fe901974e5c7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00014_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00014_00005_U (
.fgallag_sel( I080f931dfef9d8adfb1dc1ee073eb64c[fgallag_SEL-1:0]),
.fgallag( fgallag_00014_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00014_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00014_00005 };

assign fgallag_final_00014_00005 = (I080f931dfef9d8adfb1dc1ee073eb64c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00014_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00014_00006_U (
.fgallag_sel( Ide1106431e3565158bd81ccd6b18f3a1[fgallag_SEL-1:0]),
.fgallag( fgallag_00014_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00014_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00014_00006 };

assign fgallag_final_00014_00006 = (Ide1106431e3565158bd81ccd6b18f3a1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00014_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00014_00007_U (
.fgallag_sel( I63df19931e8d28666cccd79922cbd418[fgallag_SEL-1:0]),
.fgallag( fgallag_00014_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00014_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00014_00007 };

assign fgallag_final_00014_00007 = (I63df19931e8d28666cccd79922cbd418[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00014_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00014_00008_U (
.fgallag_sel( I9a7e4a59447048de90446f877eb06627[fgallag_SEL-1:0]),
.fgallag( fgallag_00014_00008 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00014_00008 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00014_00008 };

assign fgallag_final_00014_00008 = (I9a7e4a59447048de90446f877eb06627[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00014_00008 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00014_00009_U (
.fgallag_sel( I0917e92ed84363ca92fd2074acd74eba[fgallag_SEL-1:0]),
.fgallag( fgallag_00014_00009 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00014_00009 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00014_00009 };

assign fgallag_final_00014_00009 = (I0917e92ed84363ca92fd2074acd74eba[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00014_00009 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00015_00000_U (
.fgallag_sel( Ie3eefdf7b5561a90a6ddd9e6aa432509[fgallag_SEL-1:0]),
.fgallag( fgallag_00015_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00015_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00015_00000 };

assign fgallag_final_00015_00000 = (Ie3eefdf7b5561a90a6ddd9e6aa432509[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00015_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00015_00001_U (
.fgallag_sel( I56eeb10d11e886cff629457a640a1c76[fgallag_SEL-1:0]),
.fgallag( fgallag_00015_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00015_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00015_00001 };

assign fgallag_final_00015_00001 = (I56eeb10d11e886cff629457a640a1c76[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00015_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00015_00002_U (
.fgallag_sel( I7a9eea89c4e76d856df44b6bdc332840[fgallag_SEL-1:0]),
.fgallag( fgallag_00015_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00015_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00015_00002 };

assign fgallag_final_00015_00002 = (I7a9eea89c4e76d856df44b6bdc332840[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00015_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00015_00003_U (
.fgallag_sel( If8d8f4333e893788fcb9ec54256e5b7a[fgallag_SEL-1:0]),
.fgallag( fgallag_00015_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00015_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00015_00003 };

assign fgallag_final_00015_00003 = (If8d8f4333e893788fcb9ec54256e5b7a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00015_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00015_00004_U (
.fgallag_sel( Ie4af0e7e04778d85f5dee73da33376a8[fgallag_SEL-1:0]),
.fgallag( fgallag_00015_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00015_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00015_00004 };

assign fgallag_final_00015_00004 = (Ie4af0e7e04778d85f5dee73da33376a8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00015_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00015_00005_U (
.fgallag_sel( I019a4e997adf54f5f5ca651f80b7901b[fgallag_SEL-1:0]),
.fgallag( fgallag_00015_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00015_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00015_00005 };

assign fgallag_final_00015_00005 = (I019a4e997adf54f5f5ca651f80b7901b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00015_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00015_00006_U (
.fgallag_sel( I10294667f09abbfd4e2f757c414072fc[fgallag_SEL-1:0]),
.fgallag( fgallag_00015_00006 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00015_00006 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00015_00006 };

assign fgallag_final_00015_00006 = (I10294667f09abbfd4e2f757c414072fc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00015_00006 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00015_00007_U (
.fgallag_sel( Id4e8ab8f15b36bd27d1e4ebc5cbe1495[fgallag_SEL-1:0]),
.fgallag( fgallag_00015_00007 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00015_00007 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00015_00007 };

assign fgallag_final_00015_00007 = (Id4e8ab8f15b36bd27d1e4ebc5cbe1495[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00015_00007 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00015_00008_U (
.fgallag_sel( I6c93588ca9e7c623d75314da39e89a91[fgallag_SEL-1:0]),
.fgallag( fgallag_00015_00008 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00015_00008 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00015_00008 };

assign fgallag_final_00015_00008 = (I6c93588ca9e7c623d75314da39e89a91[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00015_00008 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00015_00009_U (
.fgallag_sel( I1020412efc78d12a9ebcbaeb83e5dcea[fgallag_SEL-1:0]),
.fgallag( fgallag_00015_00009 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00015_00009 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00015_00009 };

assign fgallag_final_00015_00009 = (I1020412efc78d12a9ebcbaeb83e5dcea[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00015_00009 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00016_00000_U (
.fgallag_sel( Id0b574f35a83dcfd4481a10043cd1884[fgallag_SEL-1:0]),
.fgallag( fgallag_00016_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00016_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00016_00000 };

assign fgallag_final_00016_00000 = (Id0b574f35a83dcfd4481a10043cd1884[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00016_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00016_00001_U (
.fgallag_sel( Ifc577e5c2c7288373a8c5e3969ac1589[fgallag_SEL-1:0]),
.fgallag( fgallag_00016_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00016_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00016_00001 };

assign fgallag_final_00016_00001 = (Ifc577e5c2c7288373a8c5e3969ac1589[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00016_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00016_00002_U (
.fgallag_sel( Id18a1a17c1cf6e8a2492aa73b62898f2[fgallag_SEL-1:0]),
.fgallag( fgallag_00016_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00016_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00016_00002 };

assign fgallag_final_00016_00002 = (Id18a1a17c1cf6e8a2492aa73b62898f2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00016_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00016_00003_U (
.fgallag_sel( Id8ce8f636723b9f119bb86c25017e6b3[fgallag_SEL-1:0]),
.fgallag( fgallag_00016_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00016_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00016_00003 };

assign fgallag_final_00016_00003 = (Id8ce8f636723b9f119bb86c25017e6b3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00016_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00017_00000_U (
.fgallag_sel( Ic29a18d8d504a2d5280c1d7771346518[fgallag_SEL-1:0]),
.fgallag( fgallag_00017_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00017_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00017_00000 };

assign fgallag_final_00017_00000 = (Ic29a18d8d504a2d5280c1d7771346518[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00017_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00017_00001_U (
.fgallag_sel( I96a79193aa2956b8f901d5fcc9cf65cf[fgallag_SEL-1:0]),
.fgallag( fgallag_00017_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00017_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00017_00001 };

assign fgallag_final_00017_00001 = (I96a79193aa2956b8f901d5fcc9cf65cf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00017_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00017_00002_U (
.fgallag_sel( I8c97a246c749fbef029f8b1671c772bd[fgallag_SEL-1:0]),
.fgallag( fgallag_00017_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00017_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00017_00002 };

assign fgallag_final_00017_00002 = (I8c97a246c749fbef029f8b1671c772bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00017_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00017_00003_U (
.fgallag_sel( If9ba9d221909ce7499725f6fd7d519f8[fgallag_SEL-1:0]),
.fgallag( fgallag_00017_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00017_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00017_00003 };

assign fgallag_final_00017_00003 = (If9ba9d221909ce7499725f6fd7d519f8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00017_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00018_00000_U (
.fgallag_sel( I53a7878f44253f0f1a82d9d27b1a44c3[fgallag_SEL-1:0]),
.fgallag( fgallag_00018_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00018_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00018_00000 };

assign fgallag_final_00018_00000 = (I53a7878f44253f0f1a82d9d27b1a44c3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00018_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00018_00001_U (
.fgallag_sel( Ie0e928125f9d3d17d123d97e00f1fc34[fgallag_SEL-1:0]),
.fgallag( fgallag_00018_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00018_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00018_00001 };

assign fgallag_final_00018_00001 = (Ie0e928125f9d3d17d123d97e00f1fc34[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00018_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00018_00002_U (
.fgallag_sel( I2bd0f77efeca09eebe82ea234e9fe638[fgallag_SEL-1:0]),
.fgallag( fgallag_00018_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00018_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00018_00002 };

assign fgallag_final_00018_00002 = (I2bd0f77efeca09eebe82ea234e9fe638[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00018_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00018_00003_U (
.fgallag_sel( I94f2e7ef9b3463bd598dc9049f6fb0ef[fgallag_SEL-1:0]),
.fgallag( fgallag_00018_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00018_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00018_00003 };

assign fgallag_final_00018_00003 = (I94f2e7ef9b3463bd598dc9049f6fb0ef[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00018_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00019_00000_U (
.fgallag_sel( I6dc16510af6b61b79b339d0fce77ac24[fgallag_SEL-1:0]),
.fgallag( fgallag_00019_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00019_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00019_00000 };

assign fgallag_final_00019_00000 = (I6dc16510af6b61b79b339d0fce77ac24[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00019_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00019_00001_U (
.fgallag_sel( Ic655e213ab81f5d61a018d3ed7016b12[fgallag_SEL-1:0]),
.fgallag( fgallag_00019_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00019_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00019_00001 };

assign fgallag_final_00019_00001 = (Ic655e213ab81f5d61a018d3ed7016b12[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00019_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00019_00002_U (
.fgallag_sel( I2ffc4a604025a2f5c4e273c1d070a725[fgallag_SEL-1:0]),
.fgallag( fgallag_00019_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00019_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00019_00002 };

assign fgallag_final_00019_00002 = (I2ffc4a604025a2f5c4e273c1d070a725[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00019_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00019_00003_U (
.fgallag_sel( I1c76818a9a3b688ca897aa479f7d807f[fgallag_SEL-1:0]),
.fgallag( fgallag_00019_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00019_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00019_00003 };

assign fgallag_final_00019_00003 = (I1c76818a9a3b688ca897aa479f7d807f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00019_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00020_00000_U (
.fgallag_sel( I3bfee9d3d88f0569010a4e0101200c19[fgallag_SEL-1:0]),
.fgallag( fgallag_00020_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00020_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00020_00000 };

assign fgallag_final_00020_00000 = (I3bfee9d3d88f0569010a4e0101200c19[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00020_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00020_00001_U (
.fgallag_sel( I5d4738755a26beb6d0f61dd3dec0f804[fgallag_SEL-1:0]),
.fgallag( fgallag_00020_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00020_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00020_00001 };

assign fgallag_final_00020_00001 = (I5d4738755a26beb6d0f61dd3dec0f804[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00020_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00020_00002_U (
.fgallag_sel( I2f3c800091275bcb72d1a2a38fba53f3[fgallag_SEL-1:0]),
.fgallag( fgallag_00020_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00020_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00020_00002 };

assign fgallag_final_00020_00002 = (I2f3c800091275bcb72d1a2a38fba53f3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00020_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00020_00003_U (
.fgallag_sel( I378e67cca7c4ff6325683f8346963210[fgallag_SEL-1:0]),
.fgallag( fgallag_00020_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00020_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00020_00003 };

assign fgallag_final_00020_00003 = (I378e67cca7c4ff6325683f8346963210[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00020_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00020_00004_U (
.fgallag_sel( I04c8915a7f4bbde003f7facc84435c1a[fgallag_SEL-1:0]),
.fgallag( fgallag_00020_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00020_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00020_00004 };

assign fgallag_final_00020_00004 = (I04c8915a7f4bbde003f7facc84435c1a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00020_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00020_00005_U (
.fgallag_sel( I3f50b10072f38b6addee6845e6df9118[fgallag_SEL-1:0]),
.fgallag( fgallag_00020_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00020_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00020_00005 };

assign fgallag_final_00020_00005 = (I3f50b10072f38b6addee6845e6df9118[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00020_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00021_00000_U (
.fgallag_sel( Icc60eb18ba740036d2a17f98f15cfb98[fgallag_SEL-1:0]),
.fgallag( fgallag_00021_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00021_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00021_00000 };

assign fgallag_final_00021_00000 = (Icc60eb18ba740036d2a17f98f15cfb98[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00021_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00021_00001_U (
.fgallag_sel( I1677daa18aa8b226753b1a887b9420d1[fgallag_SEL-1:0]),
.fgallag( fgallag_00021_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00021_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00021_00001 };

assign fgallag_final_00021_00001 = (I1677daa18aa8b226753b1a887b9420d1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00021_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00021_00002_U (
.fgallag_sel( I36bc2d4c9a4480daa9b0944c08b50738[fgallag_SEL-1:0]),
.fgallag( fgallag_00021_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00021_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00021_00002 };

assign fgallag_final_00021_00002 = (I36bc2d4c9a4480daa9b0944c08b50738[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00021_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00021_00003_U (
.fgallag_sel( I38419a6905f50135a6783aacca0384dd[fgallag_SEL-1:0]),
.fgallag( fgallag_00021_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00021_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00021_00003 };

assign fgallag_final_00021_00003 = (I38419a6905f50135a6783aacca0384dd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00021_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00021_00004_U (
.fgallag_sel( Ib48892dcb0715987289662a14672611e[fgallag_SEL-1:0]),
.fgallag( fgallag_00021_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00021_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00021_00004 };

assign fgallag_final_00021_00004 = (Ib48892dcb0715987289662a14672611e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00021_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00021_00005_U (
.fgallag_sel( Icd9c94f929dbc71c9b836fda3019630b[fgallag_SEL-1:0]),
.fgallag( fgallag_00021_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00021_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00021_00005 };

assign fgallag_final_00021_00005 = (Icd9c94f929dbc71c9b836fda3019630b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00021_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00022_00000_U (
.fgallag_sel( I5d0249d9a772805b3fba3f3c7f5d35bd[fgallag_SEL-1:0]),
.fgallag( fgallag_00022_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00022_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00022_00000 };

assign fgallag_final_00022_00000 = (I5d0249d9a772805b3fba3f3c7f5d35bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00022_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00022_00001_U (
.fgallag_sel( Ie97341deb6fb24d49eb8b96bd0fd3f35[fgallag_SEL-1:0]),
.fgallag( fgallag_00022_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00022_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00022_00001 };

assign fgallag_final_00022_00001 = (Ie97341deb6fb24d49eb8b96bd0fd3f35[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00022_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00022_00002_U (
.fgallag_sel( I17dd788f9d8e91307b6b1ab7488f9ce2[fgallag_SEL-1:0]),
.fgallag( fgallag_00022_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00022_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00022_00002 };

assign fgallag_final_00022_00002 = (I17dd788f9d8e91307b6b1ab7488f9ce2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00022_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00022_00003_U (
.fgallag_sel( I92ae370022ed107b152b10fd0aa3d2b7[fgallag_SEL-1:0]),
.fgallag( fgallag_00022_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00022_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00022_00003 };

assign fgallag_final_00022_00003 = (I92ae370022ed107b152b10fd0aa3d2b7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00022_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00022_00004_U (
.fgallag_sel( Iebb39f0d19ec1208bbfba6cf67a3bfc7[fgallag_SEL-1:0]),
.fgallag( fgallag_00022_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00022_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00022_00004 };

assign fgallag_final_00022_00004 = (Iebb39f0d19ec1208bbfba6cf67a3bfc7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00022_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00022_00005_U (
.fgallag_sel( I81861f6bb8bbbab6e93407cfb4a852b8[fgallag_SEL-1:0]),
.fgallag( fgallag_00022_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00022_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00022_00005 };

assign fgallag_final_00022_00005 = (I81861f6bb8bbbab6e93407cfb4a852b8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00022_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00023_00000_U (
.fgallag_sel( I217b2e3ca0a534fc5b1910adf3c1b57d[fgallag_SEL-1:0]),
.fgallag( fgallag_00023_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00023_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00023_00000 };

assign fgallag_final_00023_00000 = (I217b2e3ca0a534fc5b1910adf3c1b57d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00023_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00023_00001_U (
.fgallag_sel( I8429b08891dc56af24c72ce1b7725457[fgallag_SEL-1:0]),
.fgallag( fgallag_00023_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00023_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00023_00001 };

assign fgallag_final_00023_00001 = (I8429b08891dc56af24c72ce1b7725457[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00023_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00023_00002_U (
.fgallag_sel( If96747262303f6c5c6b129e39224bd23[fgallag_SEL-1:0]),
.fgallag( fgallag_00023_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00023_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00023_00002 };

assign fgallag_final_00023_00002 = (If96747262303f6c5c6b129e39224bd23[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00023_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00023_00003_U (
.fgallag_sel( If7012457af15c405baeaa1710319b541[fgallag_SEL-1:0]),
.fgallag( fgallag_00023_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00023_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00023_00003 };

assign fgallag_final_00023_00003 = (If7012457af15c405baeaa1710319b541[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00023_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00023_00004_U (
.fgallag_sel( Ia0a0229ef71b85195352bb664ea4e4e3[fgallag_SEL-1:0]),
.fgallag( fgallag_00023_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00023_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00023_00004 };

assign fgallag_final_00023_00004 = (Ia0a0229ef71b85195352bb664ea4e4e3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00023_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00023_00005_U (
.fgallag_sel( I42aeb7c23accc2ca874c7f8221c3af93[fgallag_SEL-1:0]),
.fgallag( fgallag_00023_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00023_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00023_00005 };

assign fgallag_final_00023_00005 = (I42aeb7c23accc2ca874c7f8221c3af93[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00023_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00024_00000_U (
.fgallag_sel( I7df6a95bf51f40693c439c6df36510d4[fgallag_SEL-1:0]),
.fgallag( fgallag_00024_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00024_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00024_00000 };

assign fgallag_final_00024_00000 = (I7df6a95bf51f40693c439c6df36510d4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00024_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00024_00001_U (
.fgallag_sel( I8fe65f9c344d7ec8657f192abefc3fb6[fgallag_SEL-1:0]),
.fgallag( fgallag_00024_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00024_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00024_00001 };

assign fgallag_final_00024_00001 = (I8fe65f9c344d7ec8657f192abefc3fb6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00024_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00024_00002_U (
.fgallag_sel( I4d75c95d34d8d8aeeb528456bbe136e1[fgallag_SEL-1:0]),
.fgallag( fgallag_00024_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00024_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00024_00002 };

assign fgallag_final_00024_00002 = (I4d75c95d34d8d8aeeb528456bbe136e1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00024_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00024_00003_U (
.fgallag_sel( I43746054a38c9521f8da9db9d0e91f99[fgallag_SEL-1:0]),
.fgallag( fgallag_00024_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00024_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00024_00003 };

assign fgallag_final_00024_00003 = (I43746054a38c9521f8da9db9d0e91f99[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00024_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00024_00004_U (
.fgallag_sel( I0430ac2a4b2b2e2fc7f8154bf946553c[fgallag_SEL-1:0]),
.fgallag( fgallag_00024_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00024_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00024_00004 };

assign fgallag_final_00024_00004 = (I0430ac2a4b2b2e2fc7f8154bf946553c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00024_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00024_00005_U (
.fgallag_sel( I25dc807fd55b81c9f24fd0d1edcaa758[fgallag_SEL-1:0]),
.fgallag( fgallag_00024_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00024_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00024_00005 };

assign fgallag_final_00024_00005 = (I25dc807fd55b81c9f24fd0d1edcaa758[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00024_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00025_00000_U (
.fgallag_sel( I7881184f1779b9fd4fdf329c5f7664da[fgallag_SEL-1:0]),
.fgallag( fgallag_00025_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00025_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00025_00000 };

assign fgallag_final_00025_00000 = (I7881184f1779b9fd4fdf329c5f7664da[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00025_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00025_00001_U (
.fgallag_sel( I8e6de2d692a307ee8a5a4b2a9265a633[fgallag_SEL-1:0]),
.fgallag( fgallag_00025_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00025_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00025_00001 };

assign fgallag_final_00025_00001 = (I8e6de2d692a307ee8a5a4b2a9265a633[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00025_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00025_00002_U (
.fgallag_sel( I54b2b18ab051b468808a3d0fc4bc893f[fgallag_SEL-1:0]),
.fgallag( fgallag_00025_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00025_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00025_00002 };

assign fgallag_final_00025_00002 = (I54b2b18ab051b468808a3d0fc4bc893f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00025_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00025_00003_U (
.fgallag_sel( I37ee86e2ca32832862cb57efe76bbedf[fgallag_SEL-1:0]),
.fgallag( fgallag_00025_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00025_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00025_00003 };

assign fgallag_final_00025_00003 = (I37ee86e2ca32832862cb57efe76bbedf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00025_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00025_00004_U (
.fgallag_sel( Ic95f2fc697574803c0f7fa35c2609f0c[fgallag_SEL-1:0]),
.fgallag( fgallag_00025_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00025_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00025_00004 };

assign fgallag_final_00025_00004 = (Ic95f2fc697574803c0f7fa35c2609f0c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00025_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00025_00005_U (
.fgallag_sel( I933a30c52c9bec5172530b2d739a3b63[fgallag_SEL-1:0]),
.fgallag( fgallag_00025_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00025_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00025_00005 };

assign fgallag_final_00025_00005 = (I933a30c52c9bec5172530b2d739a3b63[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00025_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00026_00000_U (
.fgallag_sel( I7bbd7df18f85197c22fe8cfe37312af6[fgallag_SEL-1:0]),
.fgallag( fgallag_00026_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00026_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00026_00000 };

assign fgallag_final_00026_00000 = (I7bbd7df18f85197c22fe8cfe37312af6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00026_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00026_00001_U (
.fgallag_sel( I50d5ada7c91c7af16492c6b41151b68f[fgallag_SEL-1:0]),
.fgallag( fgallag_00026_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00026_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00026_00001 };

assign fgallag_final_00026_00001 = (I50d5ada7c91c7af16492c6b41151b68f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00026_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00026_00002_U (
.fgallag_sel( I32c8e7996b3473d4906c40018799a16b[fgallag_SEL-1:0]),
.fgallag( fgallag_00026_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00026_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00026_00002 };

assign fgallag_final_00026_00002 = (I32c8e7996b3473d4906c40018799a16b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00026_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00026_00003_U (
.fgallag_sel( Ic0eacd5a4812ad7ae3fa251ab2db4694[fgallag_SEL-1:0]),
.fgallag( fgallag_00026_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00026_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00026_00003 };

assign fgallag_final_00026_00003 = (Ic0eacd5a4812ad7ae3fa251ab2db4694[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00026_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00026_00004_U (
.fgallag_sel( Ideecf8ab87d28a840cd93851169ab05b[fgallag_SEL-1:0]),
.fgallag( fgallag_00026_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00026_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00026_00004 };

assign fgallag_final_00026_00004 = (Ideecf8ab87d28a840cd93851169ab05b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00026_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00026_00005_U (
.fgallag_sel( I1ac6775eb38457b7962241d2e7336b0d[fgallag_SEL-1:0]),
.fgallag( fgallag_00026_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00026_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00026_00005 };

assign fgallag_final_00026_00005 = (I1ac6775eb38457b7962241d2e7336b0d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00026_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00027_00000_U (
.fgallag_sel( I2ecaa89698604fddd863d7e28d643a57[fgallag_SEL-1:0]),
.fgallag( fgallag_00027_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00027_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00027_00000 };

assign fgallag_final_00027_00000 = (I2ecaa89698604fddd863d7e28d643a57[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00027_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00027_00001_U (
.fgallag_sel( I273e0fe9c51c8549c8dfff393ca2e4e1[fgallag_SEL-1:0]),
.fgallag( fgallag_00027_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00027_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00027_00001 };

assign fgallag_final_00027_00001 = (I273e0fe9c51c8549c8dfff393ca2e4e1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00027_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00027_00002_U (
.fgallag_sel( Ifb1fc76002f6920a1f44c7b1bbcd0020[fgallag_SEL-1:0]),
.fgallag( fgallag_00027_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00027_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00027_00002 };

assign fgallag_final_00027_00002 = (Ifb1fc76002f6920a1f44c7b1bbcd0020[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00027_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00027_00003_U (
.fgallag_sel( Idf6d4e3aa753aa396a9bffb27732f851[fgallag_SEL-1:0]),
.fgallag( fgallag_00027_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00027_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00027_00003 };

assign fgallag_final_00027_00003 = (Idf6d4e3aa753aa396a9bffb27732f851[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00027_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00027_00004_U (
.fgallag_sel( If14ca1f5d1c2977f9da79eaebaad1bf9[fgallag_SEL-1:0]),
.fgallag( fgallag_00027_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00027_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00027_00004 };

assign fgallag_final_00027_00004 = (If14ca1f5d1c2977f9da79eaebaad1bf9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00027_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00027_00005_U (
.fgallag_sel( If8f1505d9f10e30bd3320f500d34932f[fgallag_SEL-1:0]),
.fgallag( fgallag_00027_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00027_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00027_00005 };

assign fgallag_final_00027_00005 = (If8f1505d9f10e30bd3320f500d34932f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00027_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00028_00000_U (
.fgallag_sel( Id32aa77c6406b35a00168bb5452b12fb[fgallag_SEL-1:0]),
.fgallag( fgallag_00028_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00028_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00028_00000 };

assign fgallag_final_00028_00000 = (Id32aa77c6406b35a00168bb5452b12fb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00028_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00028_00001_U (
.fgallag_sel( I9a73686acefeb361337511f6943b036b[fgallag_SEL-1:0]),
.fgallag( fgallag_00028_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00028_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00028_00001 };

assign fgallag_final_00028_00001 = (I9a73686acefeb361337511f6943b036b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00028_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00028_00002_U (
.fgallag_sel( Ib6eb7ce5a070f3a87bcf0e18be8c855d[fgallag_SEL-1:0]),
.fgallag( fgallag_00028_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00028_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00028_00002 };

assign fgallag_final_00028_00002 = (Ib6eb7ce5a070f3a87bcf0e18be8c855d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00028_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00028_00003_U (
.fgallag_sel( If69b0b717c35d33fc8c0e59b07eb9edc[fgallag_SEL-1:0]),
.fgallag( fgallag_00028_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00028_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00028_00003 };

assign fgallag_final_00028_00003 = (If69b0b717c35d33fc8c0e59b07eb9edc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00028_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00028_00004_U (
.fgallag_sel( Ibb0d73078b779585e6b0e228391ecb96[fgallag_SEL-1:0]),
.fgallag( fgallag_00028_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00028_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00028_00004 };

assign fgallag_final_00028_00004 = (Ibb0d73078b779585e6b0e228391ecb96[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00028_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00028_00005_U (
.fgallag_sel( I2894546e399fe3e33d7579772a1310df[fgallag_SEL-1:0]),
.fgallag( fgallag_00028_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00028_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00028_00005 };

assign fgallag_final_00028_00005 = (I2894546e399fe3e33d7579772a1310df[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00028_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00029_00000_U (
.fgallag_sel( I97f99a266267859aed199b278a430417[fgallag_SEL-1:0]),
.fgallag( fgallag_00029_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00029_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00029_00000 };

assign fgallag_final_00029_00000 = (I97f99a266267859aed199b278a430417[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00029_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00029_00001_U (
.fgallag_sel( Ie18cc792329941a3654322376a937d8d[fgallag_SEL-1:0]),
.fgallag( fgallag_00029_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00029_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00029_00001 };

assign fgallag_final_00029_00001 = (Ie18cc792329941a3654322376a937d8d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00029_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00029_00002_U (
.fgallag_sel( Ie914a99f08d60b74c3c36a632a4ca9b0[fgallag_SEL-1:0]),
.fgallag( fgallag_00029_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00029_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00029_00002 };

assign fgallag_final_00029_00002 = (Ie914a99f08d60b74c3c36a632a4ca9b0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00029_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00029_00003_U (
.fgallag_sel( I82916e9dc3894ad88e12de01a68d6aa5[fgallag_SEL-1:0]),
.fgallag( fgallag_00029_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00029_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00029_00003 };

assign fgallag_final_00029_00003 = (I82916e9dc3894ad88e12de01a68d6aa5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00029_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00029_00004_U (
.fgallag_sel( I6cbf576b3d652e34c0221f8316b5a392[fgallag_SEL-1:0]),
.fgallag( fgallag_00029_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00029_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00029_00004 };

assign fgallag_final_00029_00004 = (I6cbf576b3d652e34c0221f8316b5a392[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00029_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00029_00005_U (
.fgallag_sel( I9141b2516d7f855cd186472780af7b67[fgallag_SEL-1:0]),
.fgallag( fgallag_00029_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00029_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00029_00005 };

assign fgallag_final_00029_00005 = (I9141b2516d7f855cd186472780af7b67[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00029_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00030_00000_U (
.fgallag_sel( I07bf32ed72de9c02abf700c64853af61[fgallag_SEL-1:0]),
.fgallag( fgallag_00030_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00030_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00030_00000 };

assign fgallag_final_00030_00000 = (I07bf32ed72de9c02abf700c64853af61[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00030_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00030_00001_U (
.fgallag_sel( I52663a2999fb9571834d517538691b6f[fgallag_SEL-1:0]),
.fgallag( fgallag_00030_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00030_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00030_00001 };

assign fgallag_final_00030_00001 = (I52663a2999fb9571834d517538691b6f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00030_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00030_00002_U (
.fgallag_sel( I8dcb88c94506367aabe8d7ed62cc56c2[fgallag_SEL-1:0]),
.fgallag( fgallag_00030_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00030_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00030_00002 };

assign fgallag_final_00030_00002 = (I8dcb88c94506367aabe8d7ed62cc56c2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00030_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00030_00003_U (
.fgallag_sel( Ie676a4bee61154145391d9cc473fe91d[fgallag_SEL-1:0]),
.fgallag( fgallag_00030_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00030_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00030_00003 };

assign fgallag_final_00030_00003 = (Ie676a4bee61154145391d9cc473fe91d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00030_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00030_00004_U (
.fgallag_sel( I9502c8fbf6b48749bf9f84a89a937dfe[fgallag_SEL-1:0]),
.fgallag( fgallag_00030_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00030_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00030_00004 };

assign fgallag_final_00030_00004 = (I9502c8fbf6b48749bf9f84a89a937dfe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00030_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00030_00005_U (
.fgallag_sel( I0c91e540e7106f32ae59491d8ed1853e[fgallag_SEL-1:0]),
.fgallag( fgallag_00030_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00030_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00030_00005 };

assign fgallag_final_00030_00005 = (I0c91e540e7106f32ae59491d8ed1853e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00030_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00031_00000_U (
.fgallag_sel( Iddfb8a8e261389eb4a2a10880c19446a[fgallag_SEL-1:0]),
.fgallag( fgallag_00031_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00031_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00031_00000 };

assign fgallag_final_00031_00000 = (Iddfb8a8e261389eb4a2a10880c19446a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00031_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00031_00001_U (
.fgallag_sel( If0d55f861d4b3f0970c529024ca142d5[fgallag_SEL-1:0]),
.fgallag( fgallag_00031_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00031_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00031_00001 };

assign fgallag_final_00031_00001 = (If0d55f861d4b3f0970c529024ca142d5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00031_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00031_00002_U (
.fgallag_sel( Ib054f5d3f5cbb29a053d0e50c23cb3a8[fgallag_SEL-1:0]),
.fgallag( fgallag_00031_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00031_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00031_00002 };

assign fgallag_final_00031_00002 = (Ib054f5d3f5cbb29a053d0e50c23cb3a8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00031_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00031_00003_U (
.fgallag_sel( I1d65e9f97e93de8cc2a5dd532f8e482a[fgallag_SEL-1:0]),
.fgallag( fgallag_00031_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00031_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00031_00003 };

assign fgallag_final_00031_00003 = (I1d65e9f97e93de8cc2a5dd532f8e482a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00031_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00031_00004_U (
.fgallag_sel( I3bdeab8c87325d46e45d9e2d44756934[fgallag_SEL-1:0]),
.fgallag( fgallag_00031_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00031_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00031_00004 };

assign fgallag_final_00031_00004 = (I3bdeab8c87325d46e45d9e2d44756934[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00031_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00031_00005_U (
.fgallag_sel( If9228f7ecf19c41f4bbd8dabd0d5816c[fgallag_SEL-1:0]),
.fgallag( fgallag_00031_00005 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00031_00005 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00031_00005 };

assign fgallag_final_00031_00005 = (If9228f7ecf19c41f4bbd8dabd0d5816c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00031_00005 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00032_00000_U (
.fgallag_sel( I9e3edee214c4937d2aa462d3cffa624b[fgallag_SEL-1:0]),
.fgallag( fgallag_00032_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00032_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00032_00000 };

assign fgallag_final_00032_00000 = (I9e3edee214c4937d2aa462d3cffa624b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00032_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00032_00001_U (
.fgallag_sel( I9fcbbd2e81b006b50e2d35ed2627bf83[fgallag_SEL-1:0]),
.fgallag( fgallag_00032_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00032_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00032_00001 };

assign fgallag_final_00032_00001 = (I9fcbbd2e81b006b50e2d35ed2627bf83[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00032_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00032_00002_U (
.fgallag_sel( Ie16f3d50ad5e5581ca099549db7232d2[fgallag_SEL-1:0]),
.fgallag( fgallag_00032_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00032_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00032_00002 };

assign fgallag_final_00032_00002 = (Ie16f3d50ad5e5581ca099549db7232d2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00032_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00032_00003_U (
.fgallag_sel( I6345e93f3fa7f5eb2008dd41742afc2d[fgallag_SEL-1:0]),
.fgallag( fgallag_00032_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00032_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00032_00003 };

assign fgallag_final_00032_00003 = (I6345e93f3fa7f5eb2008dd41742afc2d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00032_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00033_00000_U (
.fgallag_sel( I698b93e10073b5d29357cde4bcac9dbe[fgallag_SEL-1:0]),
.fgallag( fgallag_00033_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00033_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00033_00000 };

assign fgallag_final_00033_00000 = (I698b93e10073b5d29357cde4bcac9dbe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00033_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00033_00001_U (
.fgallag_sel( Ie7ced910d84655790823e6173a5a314a[fgallag_SEL-1:0]),
.fgallag( fgallag_00033_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00033_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00033_00001 };

assign fgallag_final_00033_00001 = (Ie7ced910d84655790823e6173a5a314a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00033_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00033_00002_U (
.fgallag_sel( If6e3b6fd1810f6964e9024329d7cb3e3[fgallag_SEL-1:0]),
.fgallag( fgallag_00033_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00033_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00033_00002 };

assign fgallag_final_00033_00002 = (If6e3b6fd1810f6964e9024329d7cb3e3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00033_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00033_00003_U (
.fgallag_sel( If1045908c6d7476bd5507e57d08c406c[fgallag_SEL-1:0]),
.fgallag( fgallag_00033_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00033_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00033_00003 };

assign fgallag_final_00033_00003 = (If1045908c6d7476bd5507e57d08c406c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00033_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00034_00000_U (
.fgallag_sel( I4d4f6705ed77a16ff31b34bae0d8b6d9[fgallag_SEL-1:0]),
.fgallag( fgallag_00034_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00034_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00034_00000 };

assign fgallag_final_00034_00000 = (I4d4f6705ed77a16ff31b34bae0d8b6d9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00034_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00034_00001_U (
.fgallag_sel( I70a492396580ac1143d8a2f4b181e873[fgallag_SEL-1:0]),
.fgallag( fgallag_00034_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00034_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00034_00001 };

assign fgallag_final_00034_00001 = (I70a492396580ac1143d8a2f4b181e873[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00034_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00034_00002_U (
.fgallag_sel( I2fade32b5bdf245fa15289620dae2670[fgallag_SEL-1:0]),
.fgallag( fgallag_00034_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00034_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00034_00002 };

assign fgallag_final_00034_00002 = (I2fade32b5bdf245fa15289620dae2670[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00034_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00034_00003_U (
.fgallag_sel( Ie0dc166f57fea074496241a32cdb6015[fgallag_SEL-1:0]),
.fgallag( fgallag_00034_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00034_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00034_00003 };

assign fgallag_final_00034_00003 = (Ie0dc166f57fea074496241a32cdb6015[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00034_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00035_00000_U (
.fgallag_sel( If6a2518891412caa6d6d507082501f1e[fgallag_SEL-1:0]),
.fgallag( fgallag_00035_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00035_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00035_00000 };

assign fgallag_final_00035_00000 = (If6a2518891412caa6d6d507082501f1e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00035_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00035_00001_U (
.fgallag_sel( Ic9912e5a838a377b26a19d22148a64df[fgallag_SEL-1:0]),
.fgallag( fgallag_00035_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00035_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00035_00001 };

assign fgallag_final_00035_00001 = (Ic9912e5a838a377b26a19d22148a64df[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00035_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00035_00002_U (
.fgallag_sel( Ibc0fca22d16444bc17877106ca772c31[fgallag_SEL-1:0]),
.fgallag( fgallag_00035_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00035_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00035_00002 };

assign fgallag_final_00035_00002 = (Ibc0fca22d16444bc17877106ca772c31[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00035_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00035_00003_U (
.fgallag_sel( Ie4291d233597d5d676a80fd62d9bd208[fgallag_SEL-1:0]),
.fgallag( fgallag_00035_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00035_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00035_00003 };

assign fgallag_final_00035_00003 = (Ie4291d233597d5d676a80fd62d9bd208[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00035_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00036_00000_U (
.fgallag_sel( Ifc13b798d76aa70ec1877c275fb31d36[fgallag_SEL-1:0]),
.fgallag( fgallag_00036_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00036_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00036_00000 };

assign fgallag_final_00036_00000 = (Ifc13b798d76aa70ec1877c275fb31d36[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00036_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00036_00001_U (
.fgallag_sel( I57d6637f0bdab578a790e4a12ccaa16b[fgallag_SEL-1:0]),
.fgallag( fgallag_00036_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00036_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00036_00001 };

assign fgallag_final_00036_00001 = (I57d6637f0bdab578a790e4a12ccaa16b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00036_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00036_00002_U (
.fgallag_sel( If8ea04fe685b4f20cdaf9a84984d56fe[fgallag_SEL-1:0]),
.fgallag( fgallag_00036_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00036_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00036_00002 };

assign fgallag_final_00036_00002 = (If8ea04fe685b4f20cdaf9a84984d56fe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00036_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00036_00003_U (
.fgallag_sel( Ie0c86f20c28bcbe410b191b90d29bf76[fgallag_SEL-1:0]),
.fgallag( fgallag_00036_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00036_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00036_00003 };

assign fgallag_final_00036_00003 = (Ie0c86f20c28bcbe410b191b90d29bf76[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00036_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00036_00004_U (
.fgallag_sel( I3dc5d3f66726e15968a70cbf3d3b656a[fgallag_SEL-1:0]),
.fgallag( fgallag_00036_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00036_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00036_00004 };

assign fgallag_final_00036_00004 = (I3dc5d3f66726e15968a70cbf3d3b656a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00036_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00037_00000_U (
.fgallag_sel( Id674686e7ac37fd6f63846f9a9cede19[fgallag_SEL-1:0]),
.fgallag( fgallag_00037_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00037_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00037_00000 };

assign fgallag_final_00037_00000 = (Id674686e7ac37fd6f63846f9a9cede19[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00037_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00037_00001_U (
.fgallag_sel( Ie2ed9668d13d219c60f2e0614488cd42[fgallag_SEL-1:0]),
.fgallag( fgallag_00037_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00037_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00037_00001 };

assign fgallag_final_00037_00001 = (Ie2ed9668d13d219c60f2e0614488cd42[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00037_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00037_00002_U (
.fgallag_sel( I98abc995ff89934534543be93c6e3ffa[fgallag_SEL-1:0]),
.fgallag( fgallag_00037_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00037_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00037_00002 };

assign fgallag_final_00037_00002 = (I98abc995ff89934534543be93c6e3ffa[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00037_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00037_00003_U (
.fgallag_sel( I579cf9386ab7b08efa204d735335e462[fgallag_SEL-1:0]),
.fgallag( fgallag_00037_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00037_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00037_00003 };

assign fgallag_final_00037_00003 = (I579cf9386ab7b08efa204d735335e462[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00037_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00037_00004_U (
.fgallag_sel( I9efa4d729d10a6b7cc335fb765ed032c[fgallag_SEL-1:0]),
.fgallag( fgallag_00037_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00037_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00037_00004 };

assign fgallag_final_00037_00004 = (I9efa4d729d10a6b7cc335fb765ed032c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00037_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00038_00000_U (
.fgallag_sel( If9191ebc8e88d4e75f0f35897ebb1421[fgallag_SEL-1:0]),
.fgallag( fgallag_00038_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00038_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00038_00000 };

assign fgallag_final_00038_00000 = (If9191ebc8e88d4e75f0f35897ebb1421[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00038_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00038_00001_U (
.fgallag_sel( I3511287cfe69d5cedc5a8fbcad708437[fgallag_SEL-1:0]),
.fgallag( fgallag_00038_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00038_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00038_00001 };

assign fgallag_final_00038_00001 = (I3511287cfe69d5cedc5a8fbcad708437[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00038_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00038_00002_U (
.fgallag_sel( I91812179d44cb675b90d477f33ec48ad[fgallag_SEL-1:0]),
.fgallag( fgallag_00038_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00038_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00038_00002 };

assign fgallag_final_00038_00002 = (I91812179d44cb675b90d477f33ec48ad[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00038_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00038_00003_U (
.fgallag_sel( Idb04a1aae91fdc477ca38ed66789ee88[fgallag_SEL-1:0]),
.fgallag( fgallag_00038_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00038_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00038_00003 };

assign fgallag_final_00038_00003 = (Idb04a1aae91fdc477ca38ed66789ee88[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00038_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00038_00004_U (
.fgallag_sel( I566054aece562960590ee28b157e4a3e[fgallag_SEL-1:0]),
.fgallag( fgallag_00038_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00038_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00038_00004 };

assign fgallag_final_00038_00004 = (I566054aece562960590ee28b157e4a3e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00038_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00039_00000_U (
.fgallag_sel( I7b2ffb762cd9ef7aa8ba224efb75c46c[fgallag_SEL-1:0]),
.fgallag( fgallag_00039_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00039_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00039_00000 };

assign fgallag_final_00039_00000 = (I7b2ffb762cd9ef7aa8ba224efb75c46c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00039_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00039_00001_U (
.fgallag_sel( Id90bbb642b0f4434d8a148a28b6b2f65[fgallag_SEL-1:0]),
.fgallag( fgallag_00039_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00039_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00039_00001 };

assign fgallag_final_00039_00001 = (Id90bbb642b0f4434d8a148a28b6b2f65[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00039_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00039_00002_U (
.fgallag_sel( Ia4e297e35d484b15adce7e1d67f582b0[fgallag_SEL-1:0]),
.fgallag( fgallag_00039_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00039_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00039_00002 };

assign fgallag_final_00039_00002 = (Ia4e297e35d484b15adce7e1d67f582b0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00039_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00039_00003_U (
.fgallag_sel( I84996b1d03b692f6f736fb04c7f91e83[fgallag_SEL-1:0]),
.fgallag( fgallag_00039_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00039_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00039_00003 };

assign fgallag_final_00039_00003 = (I84996b1d03b692f6f736fb04c7f91e83[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00039_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00039_00004_U (
.fgallag_sel( I83078cc7857fc17b30f640854a4d6be5[fgallag_SEL-1:0]),
.fgallag( fgallag_00039_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00039_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00039_00004 };

assign fgallag_final_00039_00004 = (I83078cc7857fc17b30f640854a4d6be5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00039_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00040_00000_U (
.fgallag_sel( I94bb467129904032736fb13dd636c600[fgallag_SEL-1:0]),
.fgallag( fgallag_00040_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00040_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00040_00000 };

assign fgallag_final_00040_00000 = (I94bb467129904032736fb13dd636c600[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00040_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00040_00001_U (
.fgallag_sel( Ifa76758b50f439170ecd6d86ff898bc4[fgallag_SEL-1:0]),
.fgallag( fgallag_00040_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00040_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00040_00001 };

assign fgallag_final_00040_00001 = (Ifa76758b50f439170ecd6d86ff898bc4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00040_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00040_00002_U (
.fgallag_sel( I9d831dd976e8cd5d8f6a6818601e6424[fgallag_SEL-1:0]),
.fgallag( fgallag_00040_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00040_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00040_00002 };

assign fgallag_final_00040_00002 = (I9d831dd976e8cd5d8f6a6818601e6424[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00040_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00040_00003_U (
.fgallag_sel( I474774ae149804412ed4aaf1cdcaba88[fgallag_SEL-1:0]),
.fgallag( fgallag_00040_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00040_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00040_00003 };

assign fgallag_final_00040_00003 = (I474774ae149804412ed4aaf1cdcaba88[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00040_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00040_00004_U (
.fgallag_sel( I964cdcb4e6b49a62d30c2a2540851317[fgallag_SEL-1:0]),
.fgallag( fgallag_00040_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00040_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00040_00004 };

assign fgallag_final_00040_00004 = (I964cdcb4e6b49a62d30c2a2540851317[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00040_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00041_00000_U (
.fgallag_sel( I6df268bc9f85ce88674a9165664ea84a[fgallag_SEL-1:0]),
.fgallag( fgallag_00041_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00041_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00041_00000 };

assign fgallag_final_00041_00000 = (I6df268bc9f85ce88674a9165664ea84a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00041_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00041_00001_U (
.fgallag_sel( I74fdcbe9f49f7bce1f5e31d956c5883c[fgallag_SEL-1:0]),
.fgallag( fgallag_00041_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00041_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00041_00001 };

assign fgallag_final_00041_00001 = (I74fdcbe9f49f7bce1f5e31d956c5883c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00041_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00041_00002_U (
.fgallag_sel( I4a1b8453cb7a21745d5f74ad05653ed2[fgallag_SEL-1:0]),
.fgallag( fgallag_00041_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00041_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00041_00002 };

assign fgallag_final_00041_00002 = (I4a1b8453cb7a21745d5f74ad05653ed2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00041_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00041_00003_U (
.fgallag_sel( I9c53b478b2011fac0615a152fe60d5b6[fgallag_SEL-1:0]),
.fgallag( fgallag_00041_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00041_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00041_00003 };

assign fgallag_final_00041_00003 = (I9c53b478b2011fac0615a152fe60d5b6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00041_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00041_00004_U (
.fgallag_sel( Id75dbed8f1a5befda32c60b994681013[fgallag_SEL-1:0]),
.fgallag( fgallag_00041_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00041_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00041_00004 };

assign fgallag_final_00041_00004 = (Id75dbed8f1a5befda32c60b994681013[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00041_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00042_00000_U (
.fgallag_sel( I378a59323b74623c5524f854d6e11226[fgallag_SEL-1:0]),
.fgallag( fgallag_00042_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00042_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00042_00000 };

assign fgallag_final_00042_00000 = (I378a59323b74623c5524f854d6e11226[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00042_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00042_00001_U (
.fgallag_sel( I080bf885464a0cc948a4450e9f7d1d26[fgallag_SEL-1:0]),
.fgallag( fgallag_00042_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00042_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00042_00001 };

assign fgallag_final_00042_00001 = (I080bf885464a0cc948a4450e9f7d1d26[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00042_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00042_00002_U (
.fgallag_sel( If769e73adea227de1fd85c2e89d0ba08[fgallag_SEL-1:0]),
.fgallag( fgallag_00042_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00042_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00042_00002 };

assign fgallag_final_00042_00002 = (If769e73adea227de1fd85c2e89d0ba08[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00042_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00042_00003_U (
.fgallag_sel( Ifa6a34b83225e9d9b28b14874c4444e3[fgallag_SEL-1:0]),
.fgallag( fgallag_00042_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00042_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00042_00003 };

assign fgallag_final_00042_00003 = (Ifa6a34b83225e9d9b28b14874c4444e3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00042_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00042_00004_U (
.fgallag_sel( I584b1d4d6fb7ee4f20ad9c96715cdf90[fgallag_SEL-1:0]),
.fgallag( fgallag_00042_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00042_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00042_00004 };

assign fgallag_final_00042_00004 = (I584b1d4d6fb7ee4f20ad9c96715cdf90[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00042_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00043_00000_U (
.fgallag_sel( I265f9b91fbb62164e589dcf96818c4f5[fgallag_SEL-1:0]),
.fgallag( fgallag_00043_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00043_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00043_00000 };

assign fgallag_final_00043_00000 = (I265f9b91fbb62164e589dcf96818c4f5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00043_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00043_00001_U (
.fgallag_sel( I3d59a47c88227734cf6fc0d6fd30db11[fgallag_SEL-1:0]),
.fgallag( fgallag_00043_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00043_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00043_00001 };

assign fgallag_final_00043_00001 = (I3d59a47c88227734cf6fc0d6fd30db11[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00043_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00043_00002_U (
.fgallag_sel( I6144b6df2c87ea0948d730343b42129f[fgallag_SEL-1:0]),
.fgallag( fgallag_00043_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00043_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00043_00002 };

assign fgallag_final_00043_00002 = (I6144b6df2c87ea0948d730343b42129f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00043_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00043_00003_U (
.fgallag_sel( Ia7ca7400e36ea572fba8e19bcc81ecbd[fgallag_SEL-1:0]),
.fgallag( fgallag_00043_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00043_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00043_00003 };

assign fgallag_final_00043_00003 = (Ia7ca7400e36ea572fba8e19bcc81ecbd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00043_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00043_00004_U (
.fgallag_sel( I302e61b49accf5db556b87517f2341f5[fgallag_SEL-1:0]),
.fgallag( fgallag_00043_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00043_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00043_00004 };

assign fgallag_final_00043_00004 = (I302e61b49accf5db556b87517f2341f5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00043_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00044_00000_U (
.fgallag_sel( I5d9af1abff6efe3a55c6568d936b6ec7[fgallag_SEL-1:0]),
.fgallag( fgallag_00044_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00044_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00044_00000 };

assign fgallag_final_00044_00000 = (I5d9af1abff6efe3a55c6568d936b6ec7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00044_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00044_00001_U (
.fgallag_sel( I8cde0aa611c476b5112edeb8f17f15bf[fgallag_SEL-1:0]),
.fgallag( fgallag_00044_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00044_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00044_00001 };

assign fgallag_final_00044_00001 = (I8cde0aa611c476b5112edeb8f17f15bf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00044_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00044_00002_U (
.fgallag_sel( Icaa40ec40d6d26cdf70bb5ae7d492e47[fgallag_SEL-1:0]),
.fgallag( fgallag_00044_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00044_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00044_00002 };

assign fgallag_final_00044_00002 = (Icaa40ec40d6d26cdf70bb5ae7d492e47[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00044_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00044_00003_U (
.fgallag_sel( I8346f15d822cacfeecbe5d75412cb53f[fgallag_SEL-1:0]),
.fgallag( fgallag_00044_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00044_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00044_00003 };

assign fgallag_final_00044_00003 = (I8346f15d822cacfeecbe5d75412cb53f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00044_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00044_00004_U (
.fgallag_sel( I5ee364aab320ab40c0f65feda6f53b18[fgallag_SEL-1:0]),
.fgallag( fgallag_00044_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00044_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00044_00004 };

assign fgallag_final_00044_00004 = (I5ee364aab320ab40c0f65feda6f53b18[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00044_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00045_00000_U (
.fgallag_sel( I1f0ecba054900f96cd7100741191c5f4[fgallag_SEL-1:0]),
.fgallag( fgallag_00045_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00045_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00045_00000 };

assign fgallag_final_00045_00000 = (I1f0ecba054900f96cd7100741191c5f4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00045_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00045_00001_U (
.fgallag_sel( I4faf2caf62966416118a54015908c889[fgallag_SEL-1:0]),
.fgallag( fgallag_00045_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00045_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00045_00001 };

assign fgallag_final_00045_00001 = (I4faf2caf62966416118a54015908c889[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00045_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00045_00002_U (
.fgallag_sel( Idd0329980a36f87859150530ab44b52d[fgallag_SEL-1:0]),
.fgallag( fgallag_00045_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00045_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00045_00002 };

assign fgallag_final_00045_00002 = (Idd0329980a36f87859150530ab44b52d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00045_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00045_00003_U (
.fgallag_sel( Ie66bc10dde27f08813d4d347fd7cf6ce[fgallag_SEL-1:0]),
.fgallag( fgallag_00045_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00045_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00045_00003 };

assign fgallag_final_00045_00003 = (Ie66bc10dde27f08813d4d347fd7cf6ce[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00045_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00045_00004_U (
.fgallag_sel( Ie1d8b3ea7c6603cebf2f9adb776910b7[fgallag_SEL-1:0]),
.fgallag( fgallag_00045_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00045_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00045_00004 };

assign fgallag_final_00045_00004 = (Ie1d8b3ea7c6603cebf2f9adb776910b7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00045_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00046_00000_U (
.fgallag_sel( Ia37488e9a50cf5cc08de74ade676db96[fgallag_SEL-1:0]),
.fgallag( fgallag_00046_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00046_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00046_00000 };

assign fgallag_final_00046_00000 = (Ia37488e9a50cf5cc08de74ade676db96[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00046_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00046_00001_U (
.fgallag_sel( I08aa45211cab01d567cd5eb172fd2f0c[fgallag_SEL-1:0]),
.fgallag( fgallag_00046_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00046_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00046_00001 };

assign fgallag_final_00046_00001 = (I08aa45211cab01d567cd5eb172fd2f0c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00046_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00046_00002_U (
.fgallag_sel( If4ff0c63ec1deb46412858e496451a01[fgallag_SEL-1:0]),
.fgallag( fgallag_00046_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00046_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00046_00002 };

assign fgallag_final_00046_00002 = (If4ff0c63ec1deb46412858e496451a01[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00046_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00046_00003_U (
.fgallag_sel( Ife7bfd15fc4c392b5d2288d9a4e879b3[fgallag_SEL-1:0]),
.fgallag( fgallag_00046_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00046_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00046_00003 };

assign fgallag_final_00046_00003 = (Ife7bfd15fc4c392b5d2288d9a4e879b3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00046_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00046_00004_U (
.fgallag_sel( I24ac26debafd03c7333d174e8725afd6[fgallag_SEL-1:0]),
.fgallag( fgallag_00046_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00046_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00046_00004 };

assign fgallag_final_00046_00004 = (I24ac26debafd03c7333d174e8725afd6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00046_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00047_00000_U (
.fgallag_sel( I99d80ad68e2563d0f78a0e3bb82c5328[fgallag_SEL-1:0]),
.fgallag( fgallag_00047_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00047_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00047_00000 };

assign fgallag_final_00047_00000 = (I99d80ad68e2563d0f78a0e3bb82c5328[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00047_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00047_00001_U (
.fgallag_sel( I9943733ef305983c629565c881054bbf[fgallag_SEL-1:0]),
.fgallag( fgallag_00047_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00047_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00047_00001 };

assign fgallag_final_00047_00001 = (I9943733ef305983c629565c881054bbf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00047_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00047_00002_U (
.fgallag_sel( I7cb4420bc55c03a6500f5228d31fe43c[fgallag_SEL-1:0]),
.fgallag( fgallag_00047_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00047_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00047_00002 };

assign fgallag_final_00047_00002 = (I7cb4420bc55c03a6500f5228d31fe43c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00047_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00047_00003_U (
.fgallag_sel( Ic4d19dec464359c0a9fa75148fe90c73[fgallag_SEL-1:0]),
.fgallag( fgallag_00047_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00047_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00047_00003 };

assign fgallag_final_00047_00003 = (Ic4d19dec464359c0a9fa75148fe90c73[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00047_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00047_00004_U (
.fgallag_sel( I44993416e1d22613dbd78402c37a934d[fgallag_SEL-1:0]),
.fgallag( fgallag_00047_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00047_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00047_00004 };

assign fgallag_final_00047_00004 = (I44993416e1d22613dbd78402c37a934d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00047_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00048_00000_U (
.fgallag_sel( Ibc9b94a9dea471805cb442ac6904bc97[fgallag_SEL-1:0]),
.fgallag( fgallag_00048_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00048_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00048_00000 };

assign fgallag_final_00048_00000 = (Ibc9b94a9dea471805cb442ac6904bc97[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00048_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00048_00001_U (
.fgallag_sel( I917d9f9b144d3bffafc77bddae7fba6b[fgallag_SEL-1:0]),
.fgallag( fgallag_00048_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00048_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00048_00001 };

assign fgallag_final_00048_00001 = (I917d9f9b144d3bffafc77bddae7fba6b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00048_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00048_00002_U (
.fgallag_sel( Ibc91c6c3d56bb8a14e22909c43ffec51[fgallag_SEL-1:0]),
.fgallag( fgallag_00048_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00048_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00048_00002 };

assign fgallag_final_00048_00002 = (Ibc91c6c3d56bb8a14e22909c43ffec51[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00048_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00048_00003_U (
.fgallag_sel( If7c2d3eddd96b47b6c2aea8b27c8c7f4[fgallag_SEL-1:0]),
.fgallag( fgallag_00048_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00048_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00048_00003 };

assign fgallag_final_00048_00003 = (If7c2d3eddd96b47b6c2aea8b27c8c7f4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00048_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00049_00000_U (
.fgallag_sel( I4df093ed94d26b058e97db550e347e3c[fgallag_SEL-1:0]),
.fgallag( fgallag_00049_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00049_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00049_00000 };

assign fgallag_final_00049_00000 = (I4df093ed94d26b058e97db550e347e3c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00049_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00049_00001_U (
.fgallag_sel( Ie90303b0326bee4ab203a8cf1e643da9[fgallag_SEL-1:0]),
.fgallag( fgallag_00049_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00049_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00049_00001 };

assign fgallag_final_00049_00001 = (Ie90303b0326bee4ab203a8cf1e643da9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00049_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00049_00002_U (
.fgallag_sel( I19030d352fd059156ee42c66f9270beb[fgallag_SEL-1:0]),
.fgallag( fgallag_00049_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00049_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00049_00002 };

assign fgallag_final_00049_00002 = (I19030d352fd059156ee42c66f9270beb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00049_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00049_00003_U (
.fgallag_sel( I36767a902c53a384128ae1443cf88963[fgallag_SEL-1:0]),
.fgallag( fgallag_00049_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00049_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00049_00003 };

assign fgallag_final_00049_00003 = (I36767a902c53a384128ae1443cf88963[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00049_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00050_00000_U (
.fgallag_sel( I868dffa3f07407f7996bb5bc596939b7[fgallag_SEL-1:0]),
.fgallag( fgallag_00050_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00050_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00050_00000 };

assign fgallag_final_00050_00000 = (I868dffa3f07407f7996bb5bc596939b7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00050_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00050_00001_U (
.fgallag_sel( I7d928be164d0dce8b1322ff230c053e9[fgallag_SEL-1:0]),
.fgallag( fgallag_00050_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00050_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00050_00001 };

assign fgallag_final_00050_00001 = (I7d928be164d0dce8b1322ff230c053e9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00050_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00050_00002_U (
.fgallag_sel( I98be4971a8a9a08abb3ebe474d7f0c6d[fgallag_SEL-1:0]),
.fgallag( fgallag_00050_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00050_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00050_00002 };

assign fgallag_final_00050_00002 = (I98be4971a8a9a08abb3ebe474d7f0c6d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00050_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00050_00003_U (
.fgallag_sel( I779e70dea33201e9237f29681ffd5e27[fgallag_SEL-1:0]),
.fgallag( fgallag_00050_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00050_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00050_00003 };

assign fgallag_final_00050_00003 = (I779e70dea33201e9237f29681ffd5e27[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00050_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00051_00000_U (
.fgallag_sel( Ie2262914042172ab7e08599278f36af5[fgallag_SEL-1:0]),
.fgallag( fgallag_00051_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00051_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00051_00000 };

assign fgallag_final_00051_00000 = (Ie2262914042172ab7e08599278f36af5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00051_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00051_00001_U (
.fgallag_sel( I4001323da8f7956cdd480ac2d56df929[fgallag_SEL-1:0]),
.fgallag( fgallag_00051_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00051_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00051_00001 };

assign fgallag_final_00051_00001 = (I4001323da8f7956cdd480ac2d56df929[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00051_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00051_00002_U (
.fgallag_sel( Ib1cd6731034887a0a55e405c9db3e8de[fgallag_SEL-1:0]),
.fgallag( fgallag_00051_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00051_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00051_00002 };

assign fgallag_final_00051_00002 = (Ib1cd6731034887a0a55e405c9db3e8de[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00051_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00051_00003_U (
.fgallag_sel( I51aa496e8c03944c28a908102514e6f8[fgallag_SEL-1:0]),
.fgallag( fgallag_00051_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00051_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00051_00003 };

assign fgallag_final_00051_00003 = (I51aa496e8c03944c28a908102514e6f8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00051_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00052_00000_U (
.fgallag_sel( I6415f3996318472532e161510ccc8ca3[fgallag_SEL-1:0]),
.fgallag( fgallag_00052_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00052_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00052_00000 };

assign fgallag_final_00052_00000 = (I6415f3996318472532e161510ccc8ca3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00052_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00052_00001_U (
.fgallag_sel( Ia11b671b59240988737979328c472812[fgallag_SEL-1:0]),
.fgallag( fgallag_00052_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00052_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00052_00001 };

assign fgallag_final_00052_00001 = (Ia11b671b59240988737979328c472812[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00052_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00052_00002_U (
.fgallag_sel( Id4fabe0165a117a402dc14f2f3ec626a[fgallag_SEL-1:0]),
.fgallag( fgallag_00052_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00052_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00052_00002 };

assign fgallag_final_00052_00002 = (Id4fabe0165a117a402dc14f2f3ec626a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00052_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00052_00003_U (
.fgallag_sel( I57238f501ab7278b308d76211ced8cf7[fgallag_SEL-1:0]),
.fgallag( fgallag_00052_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00052_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00052_00003 };

assign fgallag_final_00052_00003 = (I57238f501ab7278b308d76211ced8cf7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00052_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00052_00004_U (
.fgallag_sel( I9b257f8556ca4e5402637f01081b78e1[fgallag_SEL-1:0]),
.fgallag( fgallag_00052_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00052_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00052_00004 };

assign fgallag_final_00052_00004 = (I9b257f8556ca4e5402637f01081b78e1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00052_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00053_00000_U (
.fgallag_sel( I2e093412a9fa3972cea01664389d8c27[fgallag_SEL-1:0]),
.fgallag( fgallag_00053_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00053_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00053_00000 };

assign fgallag_final_00053_00000 = (I2e093412a9fa3972cea01664389d8c27[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00053_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00053_00001_U (
.fgallag_sel( I17907fd8c6975c8c642535ff929221a6[fgallag_SEL-1:0]),
.fgallag( fgallag_00053_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00053_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00053_00001 };

assign fgallag_final_00053_00001 = (I17907fd8c6975c8c642535ff929221a6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00053_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00053_00002_U (
.fgallag_sel( I3c6577b04ad56d864bbaa2c048323c11[fgallag_SEL-1:0]),
.fgallag( fgallag_00053_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00053_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00053_00002 };

assign fgallag_final_00053_00002 = (I3c6577b04ad56d864bbaa2c048323c11[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00053_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00053_00003_U (
.fgallag_sel( I6f0c341c05eaa8f35bbce4521f6e8f94[fgallag_SEL-1:0]),
.fgallag( fgallag_00053_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00053_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00053_00003 };

assign fgallag_final_00053_00003 = (I6f0c341c05eaa8f35bbce4521f6e8f94[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00053_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00053_00004_U (
.fgallag_sel( Ib72ba950ecf9ae2668374f6633a67ca7[fgallag_SEL-1:0]),
.fgallag( fgallag_00053_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00053_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00053_00004 };

assign fgallag_final_00053_00004 = (Ib72ba950ecf9ae2668374f6633a67ca7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00053_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00054_00000_U (
.fgallag_sel( I3d7c72d725f4563bb562e2992093cb02[fgallag_SEL-1:0]),
.fgallag( fgallag_00054_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00054_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00054_00000 };

assign fgallag_final_00054_00000 = (I3d7c72d725f4563bb562e2992093cb02[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00054_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00054_00001_U (
.fgallag_sel( I813c881ac61a59041be3be78f6a466c8[fgallag_SEL-1:0]),
.fgallag( fgallag_00054_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00054_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00054_00001 };

assign fgallag_final_00054_00001 = (I813c881ac61a59041be3be78f6a466c8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00054_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00054_00002_U (
.fgallag_sel( I866510e7dc721fa5aac312bc5ab5ba0a[fgallag_SEL-1:0]),
.fgallag( fgallag_00054_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00054_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00054_00002 };

assign fgallag_final_00054_00002 = (I866510e7dc721fa5aac312bc5ab5ba0a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00054_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00054_00003_U (
.fgallag_sel( Ib4432359f97849dff6ad3e0f044157bd[fgallag_SEL-1:0]),
.fgallag( fgallag_00054_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00054_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00054_00003 };

assign fgallag_final_00054_00003 = (Ib4432359f97849dff6ad3e0f044157bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00054_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00054_00004_U (
.fgallag_sel( Ic86aa6eb1b4dcc2520309089b43292e6[fgallag_SEL-1:0]),
.fgallag( fgallag_00054_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00054_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00054_00004 };

assign fgallag_final_00054_00004 = (Ic86aa6eb1b4dcc2520309089b43292e6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00054_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00055_00000_U (
.fgallag_sel( I0731115afe5c15bcf131f7ef4f05802b[fgallag_SEL-1:0]),
.fgallag( fgallag_00055_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00055_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00055_00000 };

assign fgallag_final_00055_00000 = (I0731115afe5c15bcf131f7ef4f05802b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00055_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00055_00001_U (
.fgallag_sel( Ib080b8fd34385aa7986dace4afd95267[fgallag_SEL-1:0]),
.fgallag( fgallag_00055_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00055_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00055_00001 };

assign fgallag_final_00055_00001 = (Ib080b8fd34385aa7986dace4afd95267[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00055_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00055_00002_U (
.fgallag_sel( I134890b77451d0b78afc7402a6a28048[fgallag_SEL-1:0]),
.fgallag( fgallag_00055_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00055_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00055_00002 };

assign fgallag_final_00055_00002 = (I134890b77451d0b78afc7402a6a28048[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00055_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00055_00003_U (
.fgallag_sel( I956da75f13433c1dd7a3cbd3b78922c1[fgallag_SEL-1:0]),
.fgallag( fgallag_00055_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00055_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00055_00003 };

assign fgallag_final_00055_00003 = (I956da75f13433c1dd7a3cbd3b78922c1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00055_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00055_00004_U (
.fgallag_sel( I440b26c9f1b9ccf70f97c9d5f732d38e[fgallag_SEL-1:0]),
.fgallag( fgallag_00055_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00055_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00055_00004 };

assign fgallag_final_00055_00004 = (I440b26c9f1b9ccf70f97c9d5f732d38e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00055_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00056_00000_U (
.fgallag_sel( I5e3a441faca44bffc4368d96d8fb0bfd[fgallag_SEL-1:0]),
.fgallag( fgallag_00056_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00056_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00056_00000 };

assign fgallag_final_00056_00000 = (I5e3a441faca44bffc4368d96d8fb0bfd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00056_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00056_00001_U (
.fgallag_sel( I21d7ba25247a87a1a9c245d0d1f553b0[fgallag_SEL-1:0]),
.fgallag( fgallag_00056_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00056_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00056_00001 };

assign fgallag_final_00056_00001 = (I21d7ba25247a87a1a9c245d0d1f553b0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00056_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00056_00002_U (
.fgallag_sel( I55aafa8162cfc4fccfae68cf78cd1c2b[fgallag_SEL-1:0]),
.fgallag( fgallag_00056_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00056_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00056_00002 };

assign fgallag_final_00056_00002 = (I55aafa8162cfc4fccfae68cf78cd1c2b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00056_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00056_00003_U (
.fgallag_sel( Ib99c25f0d8d6493cac4d5c816884c704[fgallag_SEL-1:0]),
.fgallag( fgallag_00056_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00056_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00056_00003 };

assign fgallag_final_00056_00003 = (Ib99c25f0d8d6493cac4d5c816884c704[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00056_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00056_00004_U (
.fgallag_sel( Iee7c9f0a0e8ca127efee008b4874edbd[fgallag_SEL-1:0]),
.fgallag( fgallag_00056_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00056_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00056_00004 };

assign fgallag_final_00056_00004 = (Iee7c9f0a0e8ca127efee008b4874edbd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00056_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00057_00000_U (
.fgallag_sel( I17b4a3baae65161387f472037ffc6fc4[fgallag_SEL-1:0]),
.fgallag( fgallag_00057_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00057_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00057_00000 };

assign fgallag_final_00057_00000 = (I17b4a3baae65161387f472037ffc6fc4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00057_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00057_00001_U (
.fgallag_sel( Ie7b7b202a968fe73f6b1e02a044414c5[fgallag_SEL-1:0]),
.fgallag( fgallag_00057_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00057_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00057_00001 };

assign fgallag_final_00057_00001 = (Ie7b7b202a968fe73f6b1e02a044414c5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00057_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00057_00002_U (
.fgallag_sel( I479ab5c0e483c36267d8248340006666[fgallag_SEL-1:0]),
.fgallag( fgallag_00057_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00057_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00057_00002 };

assign fgallag_final_00057_00002 = (I479ab5c0e483c36267d8248340006666[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00057_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00057_00003_U (
.fgallag_sel( I777bfe165e25d7fde4fc950f23db7b84[fgallag_SEL-1:0]),
.fgallag( fgallag_00057_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00057_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00057_00003 };

assign fgallag_final_00057_00003 = (I777bfe165e25d7fde4fc950f23db7b84[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00057_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00057_00004_U (
.fgallag_sel( I146d505a34ddb8d65e0a1769f623a7fd[fgallag_SEL-1:0]),
.fgallag( fgallag_00057_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00057_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00057_00004 };

assign fgallag_final_00057_00004 = (I146d505a34ddb8d65e0a1769f623a7fd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00057_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00058_00000_U (
.fgallag_sel( Ia85239bddc04bf50bcf037ed2f76d7ac[fgallag_SEL-1:0]),
.fgallag( fgallag_00058_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00058_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00058_00000 };

assign fgallag_final_00058_00000 = (Ia85239bddc04bf50bcf037ed2f76d7ac[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00058_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00058_00001_U (
.fgallag_sel( Ia7306bacf3c2b180d3261a5c1f0f4a30[fgallag_SEL-1:0]),
.fgallag( fgallag_00058_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00058_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00058_00001 };

assign fgallag_final_00058_00001 = (Ia7306bacf3c2b180d3261a5c1f0f4a30[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00058_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00058_00002_U (
.fgallag_sel( I2018147b86e47af5842c4f29d047d157[fgallag_SEL-1:0]),
.fgallag( fgallag_00058_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00058_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00058_00002 };

assign fgallag_final_00058_00002 = (I2018147b86e47af5842c4f29d047d157[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00058_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00058_00003_U (
.fgallag_sel( Id17a85459845f8a8be694c4bf1fc29c9[fgallag_SEL-1:0]),
.fgallag( fgallag_00058_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00058_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00058_00003 };

assign fgallag_final_00058_00003 = (Id17a85459845f8a8be694c4bf1fc29c9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00058_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00058_00004_U (
.fgallag_sel( Ic012b15584d9d25af38f83d0526503da[fgallag_SEL-1:0]),
.fgallag( fgallag_00058_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00058_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00058_00004 };

assign fgallag_final_00058_00004 = (Ic012b15584d9d25af38f83d0526503da[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00058_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00059_00000_U (
.fgallag_sel( I7f09bd4a45143a036ce04af11b9927f9[fgallag_SEL-1:0]),
.fgallag( fgallag_00059_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00059_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00059_00000 };

assign fgallag_final_00059_00000 = (I7f09bd4a45143a036ce04af11b9927f9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00059_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00059_00001_U (
.fgallag_sel( Ica32f94af6e6f3eaf2b724a2173fa463[fgallag_SEL-1:0]),
.fgallag( fgallag_00059_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00059_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00059_00001 };

assign fgallag_final_00059_00001 = (Ica32f94af6e6f3eaf2b724a2173fa463[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00059_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00059_00002_U (
.fgallag_sel( Ib750bb83ddfbbad2a2be8d1c8392b4ff[fgallag_SEL-1:0]),
.fgallag( fgallag_00059_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00059_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00059_00002 };

assign fgallag_final_00059_00002 = (Ib750bb83ddfbbad2a2be8d1c8392b4ff[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00059_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00059_00003_U (
.fgallag_sel( I3906ece39480f96020717c6243e8ba4c[fgallag_SEL-1:0]),
.fgallag( fgallag_00059_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00059_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00059_00003 };

assign fgallag_final_00059_00003 = (I3906ece39480f96020717c6243e8ba4c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00059_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00059_00004_U (
.fgallag_sel( Ie68ce21ade07fa53c30ebf27216b03f9[fgallag_SEL-1:0]),
.fgallag( fgallag_00059_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00059_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00059_00004 };

assign fgallag_final_00059_00004 = (Ie68ce21ade07fa53c30ebf27216b03f9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00059_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00060_00000_U (
.fgallag_sel( I6cc6fa167c0d2b4b62ddbeecea175ed2[fgallag_SEL-1:0]),
.fgallag( fgallag_00060_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00060_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00060_00000 };

assign fgallag_final_00060_00000 = (I6cc6fa167c0d2b4b62ddbeecea175ed2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00060_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00060_00001_U (
.fgallag_sel( Ibddf3468ae7c27d5a4b1388e524aa9c2[fgallag_SEL-1:0]),
.fgallag( fgallag_00060_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00060_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00060_00001 };

assign fgallag_final_00060_00001 = (Ibddf3468ae7c27d5a4b1388e524aa9c2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00060_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00060_00002_U (
.fgallag_sel( Iadcb2b3acaac2e1bb505c65d3cbe4235[fgallag_SEL-1:0]),
.fgallag( fgallag_00060_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00060_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00060_00002 };

assign fgallag_final_00060_00002 = (Iadcb2b3acaac2e1bb505c65d3cbe4235[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00060_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00060_00003_U (
.fgallag_sel( I37cd96b8b0a4939d9a70098fd8bcf452[fgallag_SEL-1:0]),
.fgallag( fgallag_00060_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00060_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00060_00003 };

assign fgallag_final_00060_00003 = (I37cd96b8b0a4939d9a70098fd8bcf452[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00060_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00061_00000_U (
.fgallag_sel( Ib34b169dcc76daee2d1aa2b2a7513af3[fgallag_SEL-1:0]),
.fgallag( fgallag_00061_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00061_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00061_00000 };

assign fgallag_final_00061_00000 = (Ib34b169dcc76daee2d1aa2b2a7513af3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00061_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00061_00001_U (
.fgallag_sel( If36fc316d6ec7c7e09eae77807b37099[fgallag_SEL-1:0]),
.fgallag( fgallag_00061_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00061_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00061_00001 };

assign fgallag_final_00061_00001 = (If36fc316d6ec7c7e09eae77807b37099[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00061_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00061_00002_U (
.fgallag_sel( Ifd214c332218ac5c0fe5aded4b952711[fgallag_SEL-1:0]),
.fgallag( fgallag_00061_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00061_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00061_00002 };

assign fgallag_final_00061_00002 = (Ifd214c332218ac5c0fe5aded4b952711[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00061_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00061_00003_U (
.fgallag_sel( Idcd0fc8f86e2b6f03606b818b8346e5a[fgallag_SEL-1:0]),
.fgallag( fgallag_00061_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00061_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00061_00003 };

assign fgallag_final_00061_00003 = (Idcd0fc8f86e2b6f03606b818b8346e5a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00061_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00062_00000_U (
.fgallag_sel( If486aa8ac2cfb46f936714812cc760df[fgallag_SEL-1:0]),
.fgallag( fgallag_00062_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00062_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00062_00000 };

assign fgallag_final_00062_00000 = (If486aa8ac2cfb46f936714812cc760df[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00062_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00062_00001_U (
.fgallag_sel( I2d8e5b5fdbda7d599423c38aaace6658[fgallag_SEL-1:0]),
.fgallag( fgallag_00062_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00062_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00062_00001 };

assign fgallag_final_00062_00001 = (I2d8e5b5fdbda7d599423c38aaace6658[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00062_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00062_00002_U (
.fgallag_sel( I6d0878fb7ec75c0a26be4dbba62f80dc[fgallag_SEL-1:0]),
.fgallag( fgallag_00062_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00062_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00062_00002 };

assign fgallag_final_00062_00002 = (I6d0878fb7ec75c0a26be4dbba62f80dc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00062_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00062_00003_U (
.fgallag_sel( I16a16ff0e8a6685a09803634da429fd2[fgallag_SEL-1:0]),
.fgallag( fgallag_00062_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00062_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00062_00003 };

assign fgallag_final_00062_00003 = (I16a16ff0e8a6685a09803634da429fd2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00062_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00063_00000_U (
.fgallag_sel( Idb211abaa54ac26e7379c64a63f7d07c[fgallag_SEL-1:0]),
.fgallag( fgallag_00063_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00063_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00063_00000 };

assign fgallag_final_00063_00000 = (Idb211abaa54ac26e7379c64a63f7d07c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00063_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00063_00001_U (
.fgallag_sel( I351205eb71acb31b59d2b4470f0ba28c[fgallag_SEL-1:0]),
.fgallag( fgallag_00063_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00063_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00063_00001 };

assign fgallag_final_00063_00001 = (I351205eb71acb31b59d2b4470f0ba28c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00063_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00063_00002_U (
.fgallag_sel( If5660c495bf7690252783d888d1ad6e8[fgallag_SEL-1:0]),
.fgallag( fgallag_00063_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00063_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00063_00002 };

assign fgallag_final_00063_00002 = (If5660c495bf7690252783d888d1ad6e8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00063_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00063_00003_U (
.fgallag_sel( I3a5229cb8e44a15560b5c7bef96e65cc[fgallag_SEL-1:0]),
.fgallag( fgallag_00063_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00063_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00063_00003 };

assign fgallag_final_00063_00003 = (I3a5229cb8e44a15560b5c7bef96e65cc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00063_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00064_00000_U (
.fgallag_sel( I889b9b0828e97fe44d8366c5ef71a8f2[fgallag_SEL-1:0]),
.fgallag( fgallag_00064_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00064_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00064_00000 };

assign fgallag_final_00064_00000 = (I889b9b0828e97fe44d8366c5ef71a8f2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00064_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00064_00001_U (
.fgallag_sel( Ie23062e00e39ead706f5b6ead233747d[fgallag_SEL-1:0]),
.fgallag( fgallag_00064_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00064_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00064_00001 };

assign fgallag_final_00064_00001 = (Ie23062e00e39ead706f5b6ead233747d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00064_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00064_00002_U (
.fgallag_sel( I8a2589544c75ecfdc31d28912c639695[fgallag_SEL-1:0]),
.fgallag( fgallag_00064_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00064_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00064_00002 };

assign fgallag_final_00064_00002 = (I8a2589544c75ecfdc31d28912c639695[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00064_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00064_00003_U (
.fgallag_sel( I5c21c59147e9c3a74c7cbbb6f2a23919[fgallag_SEL-1:0]),
.fgallag( fgallag_00064_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00064_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00064_00003 };

assign fgallag_final_00064_00003 = (I5c21c59147e9c3a74c7cbbb6f2a23919[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00064_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00064_00004_U (
.fgallag_sel( Idacd78e24408e432abbbfb0c447fdde5[fgallag_SEL-1:0]),
.fgallag( fgallag_00064_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00064_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00064_00004 };

assign fgallag_final_00064_00004 = (Idacd78e24408e432abbbfb0c447fdde5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00064_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00065_00000_U (
.fgallag_sel( I0e8b171fe5080485a7f4fef83f1f1528[fgallag_SEL-1:0]),
.fgallag( fgallag_00065_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00065_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00065_00000 };

assign fgallag_final_00065_00000 = (I0e8b171fe5080485a7f4fef83f1f1528[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00065_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00065_00001_U (
.fgallag_sel( Ib22c2bd76e6c29cc2f1440885bf24b7b[fgallag_SEL-1:0]),
.fgallag( fgallag_00065_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00065_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00065_00001 };

assign fgallag_final_00065_00001 = (Ib22c2bd76e6c29cc2f1440885bf24b7b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00065_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00065_00002_U (
.fgallag_sel( I149559fccd9def4ec1ead1fdcff3c7fd[fgallag_SEL-1:0]),
.fgallag( fgallag_00065_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00065_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00065_00002 };

assign fgallag_final_00065_00002 = (I149559fccd9def4ec1ead1fdcff3c7fd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00065_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00065_00003_U (
.fgallag_sel( Icfa8fed3239748abca27a5fc17de79c0[fgallag_SEL-1:0]),
.fgallag( fgallag_00065_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00065_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00065_00003 };

assign fgallag_final_00065_00003 = (Icfa8fed3239748abca27a5fc17de79c0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00065_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00065_00004_U (
.fgallag_sel( I2ff115fa483f080d93bada49a9566b33[fgallag_SEL-1:0]),
.fgallag( fgallag_00065_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00065_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00065_00004 };

assign fgallag_final_00065_00004 = (I2ff115fa483f080d93bada49a9566b33[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00065_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00066_00000_U (
.fgallag_sel( Ibee4f3cd2f516c29ab68e07a640ab65e[fgallag_SEL-1:0]),
.fgallag( fgallag_00066_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00066_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00066_00000 };

assign fgallag_final_00066_00000 = (Ibee4f3cd2f516c29ab68e07a640ab65e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00066_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00066_00001_U (
.fgallag_sel( Ie495ab560f59ad038992c573de7d2f5b[fgallag_SEL-1:0]),
.fgallag( fgallag_00066_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00066_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00066_00001 };

assign fgallag_final_00066_00001 = (Ie495ab560f59ad038992c573de7d2f5b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00066_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00066_00002_U (
.fgallag_sel( Ibd812def78c3a9c02f9ba45cc0413711[fgallag_SEL-1:0]),
.fgallag( fgallag_00066_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00066_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00066_00002 };

assign fgallag_final_00066_00002 = (Ibd812def78c3a9c02f9ba45cc0413711[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00066_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00066_00003_U (
.fgallag_sel( I98166634dc80201b0cefb01d9559c228[fgallag_SEL-1:0]),
.fgallag( fgallag_00066_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00066_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00066_00003 };

assign fgallag_final_00066_00003 = (I98166634dc80201b0cefb01d9559c228[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00066_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00066_00004_U (
.fgallag_sel( Ic2f03a980b5f0b042853ca746abab22b[fgallag_SEL-1:0]),
.fgallag( fgallag_00066_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00066_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00066_00004 };

assign fgallag_final_00066_00004 = (Ic2f03a980b5f0b042853ca746abab22b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00066_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00067_00000_U (
.fgallag_sel( I2807a88097d2683ebdb9e0e785e3af02[fgallag_SEL-1:0]),
.fgallag( fgallag_00067_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00067_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00067_00000 };

assign fgallag_final_00067_00000 = (I2807a88097d2683ebdb9e0e785e3af02[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00067_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00067_00001_U (
.fgallag_sel( I8bebbb3a676c8506af0768516abcd740[fgallag_SEL-1:0]),
.fgallag( fgallag_00067_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00067_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00067_00001 };

assign fgallag_final_00067_00001 = (I8bebbb3a676c8506af0768516abcd740[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00067_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00067_00002_U (
.fgallag_sel( I31d380f34691c9fe9022035f233b77e2[fgallag_SEL-1:0]),
.fgallag( fgallag_00067_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00067_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00067_00002 };

assign fgallag_final_00067_00002 = (I31d380f34691c9fe9022035f233b77e2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00067_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00067_00003_U (
.fgallag_sel( I1ffb5675c98ab5b3c62b24eb23441473[fgallag_SEL-1:0]),
.fgallag( fgallag_00067_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00067_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00067_00003 };

assign fgallag_final_00067_00003 = (I1ffb5675c98ab5b3c62b24eb23441473[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00067_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00067_00004_U (
.fgallag_sel( If56424546ec4f3445853538207ea864e[fgallag_SEL-1:0]),
.fgallag( fgallag_00067_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00067_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00067_00004 };

assign fgallag_final_00067_00004 = (If56424546ec4f3445853538207ea864e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00067_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00068_00000_U (
.fgallag_sel( I31a49be4a34d9bac2e0d815097439772[fgallag_SEL-1:0]),
.fgallag( fgallag_00068_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00068_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00068_00000 };

assign fgallag_final_00068_00000 = (I31a49be4a34d9bac2e0d815097439772[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00068_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00068_00001_U (
.fgallag_sel( I6b96a2498078953e87de223aa2236d50[fgallag_SEL-1:0]),
.fgallag( fgallag_00068_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00068_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00068_00001 };

assign fgallag_final_00068_00001 = (I6b96a2498078953e87de223aa2236d50[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00068_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00068_00002_U (
.fgallag_sel( I79bf36e298a85a42c7432f877055f0b4[fgallag_SEL-1:0]),
.fgallag( fgallag_00068_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00068_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00068_00002 };

assign fgallag_final_00068_00002 = (I79bf36e298a85a42c7432f877055f0b4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00068_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00068_00003_U (
.fgallag_sel( I90c070b9bde5da05e8a5d25d2de3ba6b[fgallag_SEL-1:0]),
.fgallag( fgallag_00068_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00068_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00068_00003 };

assign fgallag_final_00068_00003 = (I90c070b9bde5da05e8a5d25d2de3ba6b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00068_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00068_00004_U (
.fgallag_sel( I28d0e4e6d772dd58d845d91952ada300[fgallag_SEL-1:0]),
.fgallag( fgallag_00068_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00068_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00068_00004 };

assign fgallag_final_00068_00004 = (I28d0e4e6d772dd58d845d91952ada300[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00068_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00069_00000_U (
.fgallag_sel( I7232b4e277acc6f1acefcb606ca24508[fgallag_SEL-1:0]),
.fgallag( fgallag_00069_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00069_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00069_00000 };

assign fgallag_final_00069_00000 = (I7232b4e277acc6f1acefcb606ca24508[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00069_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00069_00001_U (
.fgallag_sel( I32da124c433c55f692ffa4734d0dc8fc[fgallag_SEL-1:0]),
.fgallag( fgallag_00069_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00069_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00069_00001 };

assign fgallag_final_00069_00001 = (I32da124c433c55f692ffa4734d0dc8fc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00069_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00069_00002_U (
.fgallag_sel( I56e487db14eeb8d93f494d2f11b57a49[fgallag_SEL-1:0]),
.fgallag( fgallag_00069_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00069_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00069_00002 };

assign fgallag_final_00069_00002 = (I56e487db14eeb8d93f494d2f11b57a49[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00069_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00069_00003_U (
.fgallag_sel( I94d3c02bd5b8e84926d4b3c2f56efeac[fgallag_SEL-1:0]),
.fgallag( fgallag_00069_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00069_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00069_00003 };

assign fgallag_final_00069_00003 = (I94d3c02bd5b8e84926d4b3c2f56efeac[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00069_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00069_00004_U (
.fgallag_sel( I0c35b2e9176f9a06e26ca67d036411b4[fgallag_SEL-1:0]),
.fgallag( fgallag_00069_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00069_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00069_00004 };

assign fgallag_final_00069_00004 = (I0c35b2e9176f9a06e26ca67d036411b4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00069_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00070_00000_U (
.fgallag_sel( Ia6ee7b70d0b7fe7c346760b1784e50b9[fgallag_SEL-1:0]),
.fgallag( fgallag_00070_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00070_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00070_00000 };

assign fgallag_final_00070_00000 = (Ia6ee7b70d0b7fe7c346760b1784e50b9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00070_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00070_00001_U (
.fgallag_sel( I7ce57c278c683ad045526e49bcc47412[fgallag_SEL-1:0]),
.fgallag( fgallag_00070_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00070_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00070_00001 };

assign fgallag_final_00070_00001 = (I7ce57c278c683ad045526e49bcc47412[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00070_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00070_00002_U (
.fgallag_sel( Ie3d3e681cac0bb919946ac27057409e2[fgallag_SEL-1:0]),
.fgallag( fgallag_00070_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00070_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00070_00002 };

assign fgallag_final_00070_00002 = (Ie3d3e681cac0bb919946ac27057409e2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00070_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00070_00003_U (
.fgallag_sel( I8ea0a8cdd6506c982ad75f23136bcebe[fgallag_SEL-1:0]),
.fgallag( fgallag_00070_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00070_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00070_00003 };

assign fgallag_final_00070_00003 = (I8ea0a8cdd6506c982ad75f23136bcebe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00070_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00070_00004_U (
.fgallag_sel( Ic812f8bc775c5ee6a83e2b9aeb22b2a4[fgallag_SEL-1:0]),
.fgallag( fgallag_00070_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00070_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00070_00004 };

assign fgallag_final_00070_00004 = (Ic812f8bc775c5ee6a83e2b9aeb22b2a4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00070_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00071_00000_U (
.fgallag_sel( I0f0adf7fe957b9a68772bd8a1bc163d4[fgallag_SEL-1:0]),
.fgallag( fgallag_00071_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00071_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00071_00000 };

assign fgallag_final_00071_00000 = (I0f0adf7fe957b9a68772bd8a1bc163d4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00071_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00071_00001_U (
.fgallag_sel( If09562f8d82bc1dea7c38ed51523a889[fgallag_SEL-1:0]),
.fgallag( fgallag_00071_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00071_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00071_00001 };

assign fgallag_final_00071_00001 = (If09562f8d82bc1dea7c38ed51523a889[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00071_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00071_00002_U (
.fgallag_sel( Ib0fd21d66cd89c4e5c95fbc9c7680b62[fgallag_SEL-1:0]),
.fgallag( fgallag_00071_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00071_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00071_00002 };

assign fgallag_final_00071_00002 = (Ib0fd21d66cd89c4e5c95fbc9c7680b62[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00071_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00071_00003_U (
.fgallag_sel( I5a2b2bfadc638fe3fdc31136a8f09a8d[fgallag_SEL-1:0]),
.fgallag( fgallag_00071_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00071_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00071_00003 };

assign fgallag_final_00071_00003 = (I5a2b2bfadc638fe3fdc31136a8f09a8d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00071_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00071_00004_U (
.fgallag_sel( Ica914d8c556285d6b90b35747065a6e5[fgallag_SEL-1:0]),
.fgallag( fgallag_00071_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00071_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00071_00004 };

assign fgallag_final_00071_00004 = (Ica914d8c556285d6b90b35747065a6e5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00071_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00072_00000_U (
.fgallag_sel( I00c5d739bccb0ab6d05da70fe51aafea[fgallag_SEL-1:0]),
.fgallag( fgallag_00072_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00072_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00072_00000 };

assign fgallag_final_00072_00000 = (I00c5d739bccb0ab6d05da70fe51aafea[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00072_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00072_00001_U (
.fgallag_sel( I18e448761bc014ce490b766183350312[fgallag_SEL-1:0]),
.fgallag( fgallag_00072_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00072_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00072_00001 };

assign fgallag_final_00072_00001 = (I18e448761bc014ce490b766183350312[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00072_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00072_00002_U (
.fgallag_sel( I1b5920f488e9469bd416a6af3072a30b[fgallag_SEL-1:0]),
.fgallag( fgallag_00072_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00072_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00072_00002 };

assign fgallag_final_00072_00002 = (I1b5920f488e9469bd416a6af3072a30b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00072_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00072_00003_U (
.fgallag_sel( I70b41ffed4b6d88ddff219c567b8e968[fgallag_SEL-1:0]),
.fgallag( fgallag_00072_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00072_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00072_00003 };

assign fgallag_final_00072_00003 = (I70b41ffed4b6d88ddff219c567b8e968[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00072_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00073_00000_U (
.fgallag_sel( I935e083b4561da7d015e98ca7f02854e[fgallag_SEL-1:0]),
.fgallag( fgallag_00073_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00073_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00073_00000 };

assign fgallag_final_00073_00000 = (I935e083b4561da7d015e98ca7f02854e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00073_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00073_00001_U (
.fgallag_sel( Iaca9ef263bf220d786242b88c994fd21[fgallag_SEL-1:0]),
.fgallag( fgallag_00073_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00073_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00073_00001 };

assign fgallag_final_00073_00001 = (Iaca9ef263bf220d786242b88c994fd21[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00073_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00073_00002_U (
.fgallag_sel( I92169291959eb33452b79bfd32618cbc[fgallag_SEL-1:0]),
.fgallag( fgallag_00073_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00073_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00073_00002 };

assign fgallag_final_00073_00002 = (I92169291959eb33452b79bfd32618cbc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00073_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00073_00003_U (
.fgallag_sel( I126dabc3ebb9c4157adf62b57f217bd0[fgallag_SEL-1:0]),
.fgallag( fgallag_00073_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00073_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00073_00003 };

assign fgallag_final_00073_00003 = (I126dabc3ebb9c4157adf62b57f217bd0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00073_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00074_00000_U (
.fgallag_sel( If4433b1ef2eb963cd301946958b69884[fgallag_SEL-1:0]),
.fgallag( fgallag_00074_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00074_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00074_00000 };

assign fgallag_final_00074_00000 = (If4433b1ef2eb963cd301946958b69884[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00074_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00074_00001_U (
.fgallag_sel( I67ac5b9b794787b3c4738c3366689871[fgallag_SEL-1:0]),
.fgallag( fgallag_00074_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00074_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00074_00001 };

assign fgallag_final_00074_00001 = (I67ac5b9b794787b3c4738c3366689871[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00074_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00074_00002_U (
.fgallag_sel( I4f022d70078c412bdbef158f750d3da3[fgallag_SEL-1:0]),
.fgallag( fgallag_00074_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00074_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00074_00002 };

assign fgallag_final_00074_00002 = (I4f022d70078c412bdbef158f750d3da3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00074_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00074_00003_U (
.fgallag_sel( I6be6165385f6a77aeedb88f2baaa9cab[fgallag_SEL-1:0]),
.fgallag( fgallag_00074_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00074_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00074_00003 };

assign fgallag_final_00074_00003 = (I6be6165385f6a77aeedb88f2baaa9cab[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00074_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00075_00000_U (
.fgallag_sel( Id1f7fe91547e158e1d39edffb1421ff3[fgallag_SEL-1:0]),
.fgallag( fgallag_00075_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00075_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00075_00000 };

assign fgallag_final_00075_00000 = (Id1f7fe91547e158e1d39edffb1421ff3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00075_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00075_00001_U (
.fgallag_sel( I7a51924134902612db53941390891245[fgallag_SEL-1:0]),
.fgallag( fgallag_00075_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00075_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00075_00001 };

assign fgallag_final_00075_00001 = (I7a51924134902612db53941390891245[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00075_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00075_00002_U (
.fgallag_sel( I45128b9e29dd2fdd94a78fc5ffdff2b1[fgallag_SEL-1:0]),
.fgallag( fgallag_00075_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00075_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00075_00002 };

assign fgallag_final_00075_00002 = (I45128b9e29dd2fdd94a78fc5ffdff2b1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00075_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00075_00003_U (
.fgallag_sel( I7f1082408c8ebb5be18e8f71ff9510e5[fgallag_SEL-1:0]),
.fgallag( fgallag_00075_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00075_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00075_00003 };

assign fgallag_final_00075_00003 = (I7f1082408c8ebb5be18e8f71ff9510e5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00075_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00076_00000_U (
.fgallag_sel( I655ebf19c2f4b3dde716668f9ce12e59[fgallag_SEL-1:0]),
.fgallag( fgallag_00076_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00076_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00076_00000 };

assign fgallag_final_00076_00000 = (I655ebf19c2f4b3dde716668f9ce12e59[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00076_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00076_00001_U (
.fgallag_sel( Ibc9d493a507122d92af42d858cdc4c61[fgallag_SEL-1:0]),
.fgallag( fgallag_00076_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00076_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00076_00001 };

assign fgallag_final_00076_00001 = (Ibc9d493a507122d92af42d858cdc4c61[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00076_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00076_00002_U (
.fgallag_sel( Ib3d3103e5ee4feb160a97c7e26f7102b[fgallag_SEL-1:0]),
.fgallag( fgallag_00076_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00076_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00076_00002 };

assign fgallag_final_00076_00002 = (Ib3d3103e5ee4feb160a97c7e26f7102b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00076_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00076_00003_U (
.fgallag_sel( I6cc56b119e72175df3b7ce64dc3d9305[fgallag_SEL-1:0]),
.fgallag( fgallag_00076_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00076_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00076_00003 };

assign fgallag_final_00076_00003 = (I6cc56b119e72175df3b7ce64dc3d9305[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00076_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00077_00000_U (
.fgallag_sel( I57cf4a9378f1cdd94a1a5608dc57e05f[fgallag_SEL-1:0]),
.fgallag( fgallag_00077_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00077_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00077_00000 };

assign fgallag_final_00077_00000 = (I57cf4a9378f1cdd94a1a5608dc57e05f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00077_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00077_00001_U (
.fgallag_sel( I4160ab1aa18e8151c0a5c23b9edeb907[fgallag_SEL-1:0]),
.fgallag( fgallag_00077_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00077_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00077_00001 };

assign fgallag_final_00077_00001 = (I4160ab1aa18e8151c0a5c23b9edeb907[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00077_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00077_00002_U (
.fgallag_sel( Ia1f183f2d904d006e46399424e06c614[fgallag_SEL-1:0]),
.fgallag( fgallag_00077_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00077_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00077_00002 };

assign fgallag_final_00077_00002 = (Ia1f183f2d904d006e46399424e06c614[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00077_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00077_00003_U (
.fgallag_sel( If979702738671323995e56108bc9376c[fgallag_SEL-1:0]),
.fgallag( fgallag_00077_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00077_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00077_00003 };

assign fgallag_final_00077_00003 = (If979702738671323995e56108bc9376c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00077_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00078_00000_U (
.fgallag_sel( Ibc96fe0a6bf1f95036f97c7d44fab575[fgallag_SEL-1:0]),
.fgallag( fgallag_00078_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00078_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00078_00000 };

assign fgallag_final_00078_00000 = (Ibc96fe0a6bf1f95036f97c7d44fab575[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00078_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00078_00001_U (
.fgallag_sel( I755a38220a693ba43701d30e7e9508ad[fgallag_SEL-1:0]),
.fgallag( fgallag_00078_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00078_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00078_00001 };

assign fgallag_final_00078_00001 = (I755a38220a693ba43701d30e7e9508ad[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00078_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00078_00002_U (
.fgallag_sel( I896fb82baa9647a14f4b5b1ecfa70a15[fgallag_SEL-1:0]),
.fgallag( fgallag_00078_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00078_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00078_00002 };

assign fgallag_final_00078_00002 = (I896fb82baa9647a14f4b5b1ecfa70a15[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00078_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00078_00003_U (
.fgallag_sel( I23d1c973d7a2048353fbb68e4a294c08[fgallag_SEL-1:0]),
.fgallag( fgallag_00078_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00078_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00078_00003 };

assign fgallag_final_00078_00003 = (I23d1c973d7a2048353fbb68e4a294c08[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00078_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00079_00000_U (
.fgallag_sel( If9fd1e08af14f2fd4ca363383f48580a[fgallag_SEL-1:0]),
.fgallag( fgallag_00079_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00079_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00079_00000 };

assign fgallag_final_00079_00000 = (If9fd1e08af14f2fd4ca363383f48580a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00079_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00079_00001_U (
.fgallag_sel( I8f3782f78d88a5c3bc93709564999b30[fgallag_SEL-1:0]),
.fgallag( fgallag_00079_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00079_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00079_00001 };

assign fgallag_final_00079_00001 = (I8f3782f78d88a5c3bc93709564999b30[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00079_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00079_00002_U (
.fgallag_sel( I986d61d79ce31f4677f3293339db6ad2[fgallag_SEL-1:0]),
.fgallag( fgallag_00079_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00079_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00079_00002 };

assign fgallag_final_00079_00002 = (I986d61d79ce31f4677f3293339db6ad2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00079_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00079_00003_U (
.fgallag_sel( Ica4d93d9fad21316002008ade5106a9d[fgallag_SEL-1:0]),
.fgallag( fgallag_00079_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00079_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00079_00003 };

assign fgallag_final_00079_00003 = (Ica4d93d9fad21316002008ade5106a9d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00079_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00080_00000_U (
.fgallag_sel( If77592d5d8bed32477fd690341e543d0[fgallag_SEL-1:0]),
.fgallag( fgallag_00080_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00080_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00080_00000 };

assign fgallag_final_00080_00000 = (If77592d5d8bed32477fd690341e543d0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00080_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00080_00001_U (
.fgallag_sel( I25b70c6b830cbfe1b41d8f289c751924[fgallag_SEL-1:0]),
.fgallag( fgallag_00080_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00080_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00080_00001 };

assign fgallag_final_00080_00001 = (I25b70c6b830cbfe1b41d8f289c751924[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00080_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00080_00002_U (
.fgallag_sel( I2a5d65eeffa18dd9af9fe36463dafd7c[fgallag_SEL-1:0]),
.fgallag( fgallag_00080_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00080_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00080_00002 };

assign fgallag_final_00080_00002 = (I2a5d65eeffa18dd9af9fe36463dafd7c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00080_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00080_00003_U (
.fgallag_sel( Ibafa6e10bd4edf5d224fdeb2f9adbf98[fgallag_SEL-1:0]),
.fgallag( fgallag_00080_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00080_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00080_00003 };

assign fgallag_final_00080_00003 = (Ibafa6e10bd4edf5d224fdeb2f9adbf98[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00080_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00081_00000_U (
.fgallag_sel( Ifc25402bd879bc5c43b4945b60cd4540[fgallag_SEL-1:0]),
.fgallag( fgallag_00081_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00081_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00081_00000 };

assign fgallag_final_00081_00000 = (Ifc25402bd879bc5c43b4945b60cd4540[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00081_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00081_00001_U (
.fgallag_sel( Iec48da6882325d8a33e0e0e845eb18a0[fgallag_SEL-1:0]),
.fgallag( fgallag_00081_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00081_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00081_00001 };

assign fgallag_final_00081_00001 = (Iec48da6882325d8a33e0e0e845eb18a0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00081_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00081_00002_U (
.fgallag_sel( I0fd05e46862fdf8e614afaa3fd478602[fgallag_SEL-1:0]),
.fgallag( fgallag_00081_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00081_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00081_00002 };

assign fgallag_final_00081_00002 = (I0fd05e46862fdf8e614afaa3fd478602[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00081_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00081_00003_U (
.fgallag_sel( I6253a59dca81842d9ab6e58cf204abbf[fgallag_SEL-1:0]),
.fgallag( fgallag_00081_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00081_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00081_00003 };

assign fgallag_final_00081_00003 = (I6253a59dca81842d9ab6e58cf204abbf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00081_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00082_00000_U (
.fgallag_sel( Ib18d64bc58b354358ee6ac16785880e2[fgallag_SEL-1:0]),
.fgallag( fgallag_00082_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00082_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00082_00000 };

assign fgallag_final_00082_00000 = (Ib18d64bc58b354358ee6ac16785880e2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00082_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00082_00001_U (
.fgallag_sel( I28689b693a7a5f761a1f252aa3ef3b67[fgallag_SEL-1:0]),
.fgallag( fgallag_00082_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00082_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00082_00001 };

assign fgallag_final_00082_00001 = (I28689b693a7a5f761a1f252aa3ef3b67[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00082_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00082_00002_U (
.fgallag_sel( I1a4e6d12f9776d5e61094e0b5edf71d9[fgallag_SEL-1:0]),
.fgallag( fgallag_00082_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00082_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00082_00002 };

assign fgallag_final_00082_00002 = (I1a4e6d12f9776d5e61094e0b5edf71d9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00082_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00082_00003_U (
.fgallag_sel( I8e1ad23b7ac662bb827a83d3709f0adb[fgallag_SEL-1:0]),
.fgallag( fgallag_00082_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00082_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00082_00003 };

assign fgallag_final_00082_00003 = (I8e1ad23b7ac662bb827a83d3709f0adb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00082_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00083_00000_U (
.fgallag_sel( I000ad2287813072cc18dad933758f2ab[fgallag_SEL-1:0]),
.fgallag( fgallag_00083_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00083_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00083_00000 };

assign fgallag_final_00083_00000 = (I000ad2287813072cc18dad933758f2ab[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00083_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00083_00001_U (
.fgallag_sel( I7bc3698b51b89ac38ba5f4b5428a0c96[fgallag_SEL-1:0]),
.fgallag( fgallag_00083_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00083_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00083_00001 };

assign fgallag_final_00083_00001 = (I7bc3698b51b89ac38ba5f4b5428a0c96[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00083_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00083_00002_U (
.fgallag_sel( I78aea1705621e2845a331c3e61a8055b[fgallag_SEL-1:0]),
.fgallag( fgallag_00083_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00083_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00083_00002 };

assign fgallag_final_00083_00002 = (I78aea1705621e2845a331c3e61a8055b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00083_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00083_00003_U (
.fgallag_sel( I0a31314c3580f5f9e61e79c133e5d794[fgallag_SEL-1:0]),
.fgallag( fgallag_00083_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00083_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00083_00003 };

assign fgallag_final_00083_00003 = (I0a31314c3580f5f9e61e79c133e5d794[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00083_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00084_00000_U (
.fgallag_sel( I0e274fd7bfc0388fef95a8ceb939ee91[fgallag_SEL-1:0]),
.fgallag( fgallag_00084_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00084_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00084_00000 };

assign fgallag_final_00084_00000 = (I0e274fd7bfc0388fef95a8ceb939ee91[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00084_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00084_00001_U (
.fgallag_sel( Id6f39ddcb73d3f4ec081a365d11d1ef4[fgallag_SEL-1:0]),
.fgallag( fgallag_00084_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00084_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00084_00001 };

assign fgallag_final_00084_00001 = (Id6f39ddcb73d3f4ec081a365d11d1ef4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00084_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00084_00002_U (
.fgallag_sel( I807770bfa86d160459d6ec3c0f4d6a0b[fgallag_SEL-1:0]),
.fgallag( fgallag_00084_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00084_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00084_00002 };

assign fgallag_final_00084_00002 = (I807770bfa86d160459d6ec3c0f4d6a0b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00084_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00084_00003_U (
.fgallag_sel( I31c89b8a11a3090bfd74b112cbc474bb[fgallag_SEL-1:0]),
.fgallag( fgallag_00084_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00084_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00084_00003 };

assign fgallag_final_00084_00003 = (I31c89b8a11a3090bfd74b112cbc474bb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00084_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00085_00000_U (
.fgallag_sel( I79b82cb1bfc72bd5a9d313b9e9c9203c[fgallag_SEL-1:0]),
.fgallag( fgallag_00085_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00085_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00085_00000 };

assign fgallag_final_00085_00000 = (I79b82cb1bfc72bd5a9d313b9e9c9203c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00085_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00085_00001_U (
.fgallag_sel( Ib1046ae03c9a77fd2c0b3e9838e9af87[fgallag_SEL-1:0]),
.fgallag( fgallag_00085_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00085_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00085_00001 };

assign fgallag_final_00085_00001 = (Ib1046ae03c9a77fd2c0b3e9838e9af87[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00085_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00085_00002_U (
.fgallag_sel( Ic63723fd43cbbbde51c233a3cca15d3f[fgallag_SEL-1:0]),
.fgallag( fgallag_00085_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00085_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00085_00002 };

assign fgallag_final_00085_00002 = (Ic63723fd43cbbbde51c233a3cca15d3f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00085_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00085_00003_U (
.fgallag_sel( I3abbb59abada1aec6941185f95f738bd[fgallag_SEL-1:0]),
.fgallag( fgallag_00085_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00085_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00085_00003 };

assign fgallag_final_00085_00003 = (I3abbb59abada1aec6941185f95f738bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00085_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00086_00000_U (
.fgallag_sel( I8d5bd7039a77ce82ce0f6cbba9c2a076[fgallag_SEL-1:0]),
.fgallag( fgallag_00086_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00086_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00086_00000 };

assign fgallag_final_00086_00000 = (I8d5bd7039a77ce82ce0f6cbba9c2a076[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00086_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00086_00001_U (
.fgallag_sel( I527ad0b9382dd7b6e657dc1a32d8e472[fgallag_SEL-1:0]),
.fgallag( fgallag_00086_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00086_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00086_00001 };

assign fgallag_final_00086_00001 = (I527ad0b9382dd7b6e657dc1a32d8e472[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00086_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00086_00002_U (
.fgallag_sel( I8de02f32e14e719f4930d99743c04a20[fgallag_SEL-1:0]),
.fgallag( fgallag_00086_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00086_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00086_00002 };

assign fgallag_final_00086_00002 = (I8de02f32e14e719f4930d99743c04a20[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00086_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00086_00003_U (
.fgallag_sel( I7614dd5e9628c761dd9b2a512cb1da98[fgallag_SEL-1:0]),
.fgallag( fgallag_00086_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00086_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00086_00003 };

assign fgallag_final_00086_00003 = (I7614dd5e9628c761dd9b2a512cb1da98[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00086_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00087_00000_U (
.fgallag_sel( Icae7efa4742dd0ad943ee1f67b0c9b14[fgallag_SEL-1:0]),
.fgallag( fgallag_00087_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00087_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00087_00000 };

assign fgallag_final_00087_00000 = (Icae7efa4742dd0ad943ee1f67b0c9b14[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00087_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00087_00001_U (
.fgallag_sel( Ieb1854b79e9a2bc6cf5aa1c319e8e753[fgallag_SEL-1:0]),
.fgallag( fgallag_00087_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00087_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00087_00001 };

assign fgallag_final_00087_00001 = (Ieb1854b79e9a2bc6cf5aa1c319e8e753[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00087_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00087_00002_U (
.fgallag_sel( Iff50b77f300183ca59a67ccbcc9573c4[fgallag_SEL-1:0]),
.fgallag( fgallag_00087_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00087_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00087_00002 };

assign fgallag_final_00087_00002 = (Iff50b77f300183ca59a67ccbcc9573c4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00087_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00087_00003_U (
.fgallag_sel( I4868604f8178663de759d4c63dc6c4bd[fgallag_SEL-1:0]),
.fgallag( fgallag_00087_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00087_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00087_00003 };

assign fgallag_final_00087_00003 = (I4868604f8178663de759d4c63dc6c4bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00087_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00088_00000_U (
.fgallag_sel( Ife992a151986c58df4cba79b6bc4ac0a[fgallag_SEL-1:0]),
.fgallag( fgallag_00088_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00088_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00088_00000 };

assign fgallag_final_00088_00000 = (Ife992a151986c58df4cba79b6bc4ac0a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00088_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00088_00001_U (
.fgallag_sel( I9ab973fb74d9fac5d78eb8fc2c7ecf36[fgallag_SEL-1:0]),
.fgallag( fgallag_00088_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00088_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00088_00001 };

assign fgallag_final_00088_00001 = (I9ab973fb74d9fac5d78eb8fc2c7ecf36[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00088_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00088_00002_U (
.fgallag_sel( I5ee7916e859b86a98538659401685016[fgallag_SEL-1:0]),
.fgallag( fgallag_00088_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00088_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00088_00002 };

assign fgallag_final_00088_00002 = (I5ee7916e859b86a98538659401685016[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00088_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00089_00000_U (
.fgallag_sel( I48c284cefb8cfb5a938a8f23ce4d7f03[fgallag_SEL-1:0]),
.fgallag( fgallag_00089_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00089_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00089_00000 };

assign fgallag_final_00089_00000 = (I48c284cefb8cfb5a938a8f23ce4d7f03[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00089_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00089_00001_U (
.fgallag_sel( I5c1fc666b77a689478654dd29519f458[fgallag_SEL-1:0]),
.fgallag( fgallag_00089_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00089_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00089_00001 };

assign fgallag_final_00089_00001 = (I5c1fc666b77a689478654dd29519f458[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00089_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00089_00002_U (
.fgallag_sel( I38bba98b59184c75ba3b27e1dcf52182[fgallag_SEL-1:0]),
.fgallag( fgallag_00089_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00089_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00089_00002 };

assign fgallag_final_00089_00002 = (I38bba98b59184c75ba3b27e1dcf52182[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00089_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00090_00000_U (
.fgallag_sel( I6905b65403c16b0211643227ece536f6[fgallag_SEL-1:0]),
.fgallag( fgallag_00090_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00090_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00090_00000 };

assign fgallag_final_00090_00000 = (I6905b65403c16b0211643227ece536f6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00090_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00090_00001_U (
.fgallag_sel( I3ed34401bba9d5f229bc98480aedd9a5[fgallag_SEL-1:0]),
.fgallag( fgallag_00090_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00090_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00090_00001 };

assign fgallag_final_00090_00001 = (I3ed34401bba9d5f229bc98480aedd9a5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00090_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00090_00002_U (
.fgallag_sel( Ib4d05804277cddc7f00ac17ac14f5325[fgallag_SEL-1:0]),
.fgallag( fgallag_00090_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00090_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00090_00002 };

assign fgallag_final_00090_00002 = (Ib4d05804277cddc7f00ac17ac14f5325[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00090_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00091_00000_U (
.fgallag_sel( I41babdca6d3fa462849592d37b0a7998[fgallag_SEL-1:0]),
.fgallag( fgallag_00091_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00091_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00091_00000 };

assign fgallag_final_00091_00000 = (I41babdca6d3fa462849592d37b0a7998[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00091_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00091_00001_U (
.fgallag_sel( I58cfec706dc929ebfdeaca6e01b00c0a[fgallag_SEL-1:0]),
.fgallag( fgallag_00091_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00091_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00091_00001 };

assign fgallag_final_00091_00001 = (I58cfec706dc929ebfdeaca6e01b00c0a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00091_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00091_00002_U (
.fgallag_sel( I7efe3c5b2fc69840a79545e0399ce749[fgallag_SEL-1:0]),
.fgallag( fgallag_00091_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00091_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00091_00002 };

assign fgallag_final_00091_00002 = (I7efe3c5b2fc69840a79545e0399ce749[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00091_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00092_00000_U (
.fgallag_sel( I70e3eeb2b3966676d16a6aa4c85753ab[fgallag_SEL-1:0]),
.fgallag( fgallag_00092_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00092_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00092_00000 };

assign fgallag_final_00092_00000 = (I70e3eeb2b3966676d16a6aa4c85753ab[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00092_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00092_00001_U (
.fgallag_sel( I2a32d545d1e7beecc7531174c7e8dfbc[fgallag_SEL-1:0]),
.fgallag( fgallag_00092_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00092_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00092_00001 };

assign fgallag_final_00092_00001 = (I2a32d545d1e7beecc7531174c7e8dfbc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00092_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00092_00002_U (
.fgallag_sel( Ib8fb40e4ba0ba1f5e9f5a99d1271ed06[fgallag_SEL-1:0]),
.fgallag( fgallag_00092_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00092_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00092_00002 };

assign fgallag_final_00092_00002 = (Ib8fb40e4ba0ba1f5e9f5a99d1271ed06[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00092_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00092_00003_U (
.fgallag_sel( Ica792cb9850a61fa4a8bd8a4b6c6ca05[fgallag_SEL-1:0]),
.fgallag( fgallag_00092_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00092_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00092_00003 };

assign fgallag_final_00092_00003 = (Ica792cb9850a61fa4a8bd8a4b6c6ca05[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00092_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00093_00000_U (
.fgallag_sel( I779e5997c66649d6d54fd7f0514c47bd[fgallag_SEL-1:0]),
.fgallag( fgallag_00093_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00093_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00093_00000 };

assign fgallag_final_00093_00000 = (I779e5997c66649d6d54fd7f0514c47bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00093_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00093_00001_U (
.fgallag_sel( I5aa578b0c2831453683fa44af1878cb8[fgallag_SEL-1:0]),
.fgallag( fgallag_00093_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00093_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00093_00001 };

assign fgallag_final_00093_00001 = (I5aa578b0c2831453683fa44af1878cb8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00093_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00093_00002_U (
.fgallag_sel( I735d6229ef1a4ecda0a1f1dbdfb53fc1[fgallag_SEL-1:0]),
.fgallag( fgallag_00093_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00093_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00093_00002 };

assign fgallag_final_00093_00002 = (I735d6229ef1a4ecda0a1f1dbdfb53fc1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00093_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00093_00003_U (
.fgallag_sel( I62affd47512c5e8f0979244115624d97[fgallag_SEL-1:0]),
.fgallag( fgallag_00093_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00093_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00093_00003 };

assign fgallag_final_00093_00003 = (I62affd47512c5e8f0979244115624d97[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00093_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00094_00000_U (
.fgallag_sel( I14fe27afb3df5531b18dc9604e8dbe65[fgallag_SEL-1:0]),
.fgallag( fgallag_00094_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00094_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00094_00000 };

assign fgallag_final_00094_00000 = (I14fe27afb3df5531b18dc9604e8dbe65[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00094_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00094_00001_U (
.fgallag_sel( Ib1b1626c84dad8ad13c058f921ffd57d[fgallag_SEL-1:0]),
.fgallag( fgallag_00094_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00094_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00094_00001 };

assign fgallag_final_00094_00001 = (Ib1b1626c84dad8ad13c058f921ffd57d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00094_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00094_00002_U (
.fgallag_sel( Idf4a4bdddb88c21c5afe10a02373a6eb[fgallag_SEL-1:0]),
.fgallag( fgallag_00094_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00094_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00094_00002 };

assign fgallag_final_00094_00002 = (Idf4a4bdddb88c21c5afe10a02373a6eb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00094_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00094_00003_U (
.fgallag_sel( Iadefc2a3d07ed4b2c3c46b2ab5dec252[fgallag_SEL-1:0]),
.fgallag( fgallag_00094_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00094_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00094_00003 };

assign fgallag_final_00094_00003 = (Iadefc2a3d07ed4b2c3c46b2ab5dec252[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00094_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00095_00000_U (
.fgallag_sel( I19315957077b037ffc6415dbb06ef789[fgallag_SEL-1:0]),
.fgallag( fgallag_00095_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00095_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00095_00000 };

assign fgallag_final_00095_00000 = (I19315957077b037ffc6415dbb06ef789[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00095_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00095_00001_U (
.fgallag_sel( I1f9be09334407fc86c83a7c127e17bbe[fgallag_SEL-1:0]),
.fgallag( fgallag_00095_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00095_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00095_00001 };

assign fgallag_final_00095_00001 = (I1f9be09334407fc86c83a7c127e17bbe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00095_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00095_00002_U (
.fgallag_sel( I28e17a5af7a7286a2643100d6d058dc0[fgallag_SEL-1:0]),
.fgallag( fgallag_00095_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00095_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00095_00002 };

assign fgallag_final_00095_00002 = (I28e17a5af7a7286a2643100d6d058dc0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00095_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00095_00003_U (
.fgallag_sel( Icb2297c397bfe56be251ffb6b249a020[fgallag_SEL-1:0]),
.fgallag( fgallag_00095_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00095_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00095_00003 };

assign fgallag_final_00095_00003 = (Icb2297c397bfe56be251ffb6b249a020[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00095_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00096_00000_U (
.fgallag_sel( I64a48984527d660002f1f82c376c7a84[fgallag_SEL-1:0]),
.fgallag( fgallag_00096_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00096_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00096_00000 };

assign fgallag_final_00096_00000 = (I64a48984527d660002f1f82c376c7a84[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00096_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00096_00001_U (
.fgallag_sel( I238b5fc70ce9f05b6322a2691b3a0207[fgallag_SEL-1:0]),
.fgallag( fgallag_00096_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00096_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00096_00001 };

assign fgallag_final_00096_00001 = (I238b5fc70ce9f05b6322a2691b3a0207[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00096_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00096_00002_U (
.fgallag_sel( I00c16e7ad3821981032a42d5baa767b3[fgallag_SEL-1:0]),
.fgallag( fgallag_00096_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00096_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00096_00002 };

assign fgallag_final_00096_00002 = (I00c16e7ad3821981032a42d5baa767b3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00096_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00096_00003_U (
.fgallag_sel( I42fd5b094da200b33036e6cb8c7d0286[fgallag_SEL-1:0]),
.fgallag( fgallag_00096_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00096_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00096_00003 };

assign fgallag_final_00096_00003 = (I42fd5b094da200b33036e6cb8c7d0286[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00096_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00097_00000_U (
.fgallag_sel( I98b7e26a0e9ec9ad750ff87cc0641a73[fgallag_SEL-1:0]),
.fgallag( fgallag_00097_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00097_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00097_00000 };

assign fgallag_final_00097_00000 = (I98b7e26a0e9ec9ad750ff87cc0641a73[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00097_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00097_00001_U (
.fgallag_sel( I3ec904916870171bf837e162d1030052[fgallag_SEL-1:0]),
.fgallag( fgallag_00097_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00097_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00097_00001 };

assign fgallag_final_00097_00001 = (I3ec904916870171bf837e162d1030052[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00097_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00097_00002_U (
.fgallag_sel( Iedb11b97900b7dd769d31f8a89521975[fgallag_SEL-1:0]),
.fgallag( fgallag_00097_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00097_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00097_00002 };

assign fgallag_final_00097_00002 = (Iedb11b97900b7dd769d31f8a89521975[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00097_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00097_00003_U (
.fgallag_sel( Id0dceec6497c9f13ada07138986d4145[fgallag_SEL-1:0]),
.fgallag( fgallag_00097_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00097_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00097_00003 };

assign fgallag_final_00097_00003 = (Id0dceec6497c9f13ada07138986d4145[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00097_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00098_00000_U (
.fgallag_sel( Ibfe7d9bac29b8838f20cdcfe8ef7da0c[fgallag_SEL-1:0]),
.fgallag( fgallag_00098_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00098_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00098_00000 };

assign fgallag_final_00098_00000 = (Ibfe7d9bac29b8838f20cdcfe8ef7da0c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00098_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00098_00001_U (
.fgallag_sel( I4d6c95605595942a34573d6ed55eb326[fgallag_SEL-1:0]),
.fgallag( fgallag_00098_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00098_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00098_00001 };

assign fgallag_final_00098_00001 = (I4d6c95605595942a34573d6ed55eb326[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00098_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00098_00002_U (
.fgallag_sel( Id6d8f32958dfa1a98958a84e7f1aed02[fgallag_SEL-1:0]),
.fgallag( fgallag_00098_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00098_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00098_00002 };

assign fgallag_final_00098_00002 = (Id6d8f32958dfa1a98958a84e7f1aed02[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00098_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00098_00003_U (
.fgallag_sel( I971cdf9ddd1bfff5664eec35f22da335[fgallag_SEL-1:0]),
.fgallag( fgallag_00098_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00098_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00098_00003 };

assign fgallag_final_00098_00003 = (I971cdf9ddd1bfff5664eec35f22da335[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00098_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00099_00000_U (
.fgallag_sel( Idd8bc1412a0dc5f489ef253a6164ceea[fgallag_SEL-1:0]),
.fgallag( fgallag_00099_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00099_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00099_00000 };

assign fgallag_final_00099_00000 = (Idd8bc1412a0dc5f489ef253a6164ceea[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00099_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00099_00001_U (
.fgallag_sel( Idbeec36de0128e5924e214877c82bf11[fgallag_SEL-1:0]),
.fgallag( fgallag_00099_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00099_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00099_00001 };

assign fgallag_final_00099_00001 = (Idbeec36de0128e5924e214877c82bf11[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00099_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00099_00002_U (
.fgallag_sel( I50a9cd240979bc56421bf85011ae99ed[fgallag_SEL-1:0]),
.fgallag( fgallag_00099_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00099_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00099_00002 };

assign fgallag_final_00099_00002 = (I50a9cd240979bc56421bf85011ae99ed[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00099_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00099_00003_U (
.fgallag_sel( I6437095f6bad2d4fb2fbe0361f60bba1[fgallag_SEL-1:0]),
.fgallag( fgallag_00099_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00099_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00099_00003 };

assign fgallag_final_00099_00003 = (I6437095f6bad2d4fb2fbe0361f60bba1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00099_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00100_00000_U (
.fgallag_sel( Ie9b6eb3bbac26635aa00c38110958d46[fgallag_SEL-1:0]),
.fgallag( fgallag_00100_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00100_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00100_00000 };

assign fgallag_final_00100_00000 = (Ie9b6eb3bbac26635aa00c38110958d46[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00100_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00100_00001_U (
.fgallag_sel( I9f34e81e3ffb85539a6273babc2a732e[fgallag_SEL-1:0]),
.fgallag( fgallag_00100_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00100_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00100_00001 };

assign fgallag_final_00100_00001 = (I9f34e81e3ffb85539a6273babc2a732e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00100_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00100_00002_U (
.fgallag_sel( Id0a1ab8472d704001e0eba0317b117d6[fgallag_SEL-1:0]),
.fgallag( fgallag_00100_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00100_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00100_00002 };

assign fgallag_final_00100_00002 = (Id0a1ab8472d704001e0eba0317b117d6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00100_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00101_00000_U (
.fgallag_sel( I9e632217cd0561d8faa28e4b8850d995[fgallag_SEL-1:0]),
.fgallag( fgallag_00101_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00101_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00101_00000 };

assign fgallag_final_00101_00000 = (I9e632217cd0561d8faa28e4b8850d995[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00101_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00101_00001_U (
.fgallag_sel( Iedeb5b7b2fa8acf1ea083102678710ea[fgallag_SEL-1:0]),
.fgallag( fgallag_00101_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00101_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00101_00001 };

assign fgallag_final_00101_00001 = (Iedeb5b7b2fa8acf1ea083102678710ea[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00101_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00101_00002_U (
.fgallag_sel( I972431d1f5af0bdf4828e4f85591e358[fgallag_SEL-1:0]),
.fgallag( fgallag_00101_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00101_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00101_00002 };

assign fgallag_final_00101_00002 = (I972431d1f5af0bdf4828e4f85591e358[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00101_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00102_00000_U (
.fgallag_sel( I1f41024b715d8312944ccbf70e95bb40[fgallag_SEL-1:0]),
.fgallag( fgallag_00102_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00102_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00102_00000 };

assign fgallag_final_00102_00000 = (I1f41024b715d8312944ccbf70e95bb40[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00102_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00102_00001_U (
.fgallag_sel( Ia6bb5ca05f5d0af452c994dd50004e1d[fgallag_SEL-1:0]),
.fgallag( fgallag_00102_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00102_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00102_00001 };

assign fgallag_final_00102_00001 = (Ia6bb5ca05f5d0af452c994dd50004e1d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00102_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00102_00002_U (
.fgallag_sel( I9a1d1d1c862808f9a769cbdb3bc634e1[fgallag_SEL-1:0]),
.fgallag( fgallag_00102_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00102_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00102_00002 };

assign fgallag_final_00102_00002 = (I9a1d1d1c862808f9a769cbdb3bc634e1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00102_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00103_00000_U (
.fgallag_sel( I9734eb86f4e73ba217739baf5cb1b13c[fgallag_SEL-1:0]),
.fgallag( fgallag_00103_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00103_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00103_00000 };

assign fgallag_final_00103_00000 = (I9734eb86f4e73ba217739baf5cb1b13c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00103_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00103_00001_U (
.fgallag_sel( Ifc0fe00f86569956df72d8a960337e8c[fgallag_SEL-1:0]),
.fgallag( fgallag_00103_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00103_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00103_00001 };

assign fgallag_final_00103_00001 = (Ifc0fe00f86569956df72d8a960337e8c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00103_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00103_00002_U (
.fgallag_sel( I223341a807a1d555f759632f67815159[fgallag_SEL-1:0]),
.fgallag( fgallag_00103_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00103_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00103_00002 };

assign fgallag_final_00103_00002 = (I223341a807a1d555f759632f67815159[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00103_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00104_00000_U (
.fgallag_sel( I6c1f5cdf5f2917118941f4af14d67fef[fgallag_SEL-1:0]),
.fgallag( fgallag_00104_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00104_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00104_00000 };

assign fgallag_final_00104_00000 = (I6c1f5cdf5f2917118941f4af14d67fef[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00104_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00104_00001_U (
.fgallag_sel( Ie84e88fd1aa2a0b90aa1715fcd27a329[fgallag_SEL-1:0]),
.fgallag( fgallag_00104_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00104_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00104_00001 };

assign fgallag_final_00104_00001 = (Ie84e88fd1aa2a0b90aa1715fcd27a329[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00104_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00104_00002_U (
.fgallag_sel( I558f70d7039a8bb58d8ea3f72e43dac0[fgallag_SEL-1:0]),
.fgallag( fgallag_00104_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00104_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00104_00002 };

assign fgallag_final_00104_00002 = (I558f70d7039a8bb58d8ea3f72e43dac0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00104_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00104_00003_U (
.fgallag_sel( I9924269ed3de12f1f2a28893c7f95292[fgallag_SEL-1:0]),
.fgallag( fgallag_00104_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00104_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00104_00003 };

assign fgallag_final_00104_00003 = (I9924269ed3de12f1f2a28893c7f95292[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00104_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00104_00004_U (
.fgallag_sel( If1153befd1396be2798cc14535ddeb8a[fgallag_SEL-1:0]),
.fgallag( fgallag_00104_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00104_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00104_00004 };

assign fgallag_final_00104_00004 = (If1153befd1396be2798cc14535ddeb8a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00104_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00105_00000_U (
.fgallag_sel( I9bc447b20687fb3e7eff45792bd4dc3a[fgallag_SEL-1:0]),
.fgallag( fgallag_00105_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00105_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00105_00000 };

assign fgallag_final_00105_00000 = (I9bc447b20687fb3e7eff45792bd4dc3a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00105_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00105_00001_U (
.fgallag_sel( If590520f01e452db9867a8d6d5dab29b[fgallag_SEL-1:0]),
.fgallag( fgallag_00105_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00105_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00105_00001 };

assign fgallag_final_00105_00001 = (If590520f01e452db9867a8d6d5dab29b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00105_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00105_00002_U (
.fgallag_sel( Id93ee7d283016ab9b0aaa21237237c54[fgallag_SEL-1:0]),
.fgallag( fgallag_00105_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00105_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00105_00002 };

assign fgallag_final_00105_00002 = (Id93ee7d283016ab9b0aaa21237237c54[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00105_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00105_00003_U (
.fgallag_sel( Ic1cf03baabaed466fe532e4db3a9ea78[fgallag_SEL-1:0]),
.fgallag( fgallag_00105_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00105_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00105_00003 };

assign fgallag_final_00105_00003 = (Ic1cf03baabaed466fe532e4db3a9ea78[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00105_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00105_00004_U (
.fgallag_sel( If3031f9aa8f6eba90eac12db7839fefd[fgallag_SEL-1:0]),
.fgallag( fgallag_00105_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00105_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00105_00004 };

assign fgallag_final_00105_00004 = (If3031f9aa8f6eba90eac12db7839fefd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00105_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00106_00000_U (
.fgallag_sel( I0dc2708970ca2b6c092273b6626bacd6[fgallag_SEL-1:0]),
.fgallag( fgallag_00106_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00106_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00106_00000 };

assign fgallag_final_00106_00000 = (I0dc2708970ca2b6c092273b6626bacd6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00106_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00106_00001_U (
.fgallag_sel( Ia58944aebf0b4f0a7d76a1444fced9de[fgallag_SEL-1:0]),
.fgallag( fgallag_00106_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00106_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00106_00001 };

assign fgallag_final_00106_00001 = (Ia58944aebf0b4f0a7d76a1444fced9de[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00106_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00106_00002_U (
.fgallag_sel( Iedd8e69679d10e05f2889f1d71cf0e7b[fgallag_SEL-1:0]),
.fgallag( fgallag_00106_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00106_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00106_00002 };

assign fgallag_final_00106_00002 = (Iedd8e69679d10e05f2889f1d71cf0e7b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00106_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00106_00003_U (
.fgallag_sel( I90f0d471914a2333b9dc14d6d01cf927[fgallag_SEL-1:0]),
.fgallag( fgallag_00106_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00106_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00106_00003 };

assign fgallag_final_00106_00003 = (I90f0d471914a2333b9dc14d6d01cf927[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00106_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00106_00004_U (
.fgallag_sel( Idceeb22013af64b6bb9f0d773e9ffe9a[fgallag_SEL-1:0]),
.fgallag( fgallag_00106_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00106_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00106_00004 };

assign fgallag_final_00106_00004 = (Idceeb22013af64b6bb9f0d773e9ffe9a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00106_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00107_00000_U (
.fgallag_sel( If43574342e60a625fb6bee5a495e88f3[fgallag_SEL-1:0]),
.fgallag( fgallag_00107_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00107_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00107_00000 };

assign fgallag_final_00107_00000 = (If43574342e60a625fb6bee5a495e88f3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00107_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00107_00001_U (
.fgallag_sel( Id285f055275014d9f23d35f91879afa1[fgallag_SEL-1:0]),
.fgallag( fgallag_00107_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00107_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00107_00001 };

assign fgallag_final_00107_00001 = (Id285f055275014d9f23d35f91879afa1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00107_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00107_00002_U (
.fgallag_sel( I8c803ab08db372802117de4fa4e2a187[fgallag_SEL-1:0]),
.fgallag( fgallag_00107_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00107_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00107_00002 };

assign fgallag_final_00107_00002 = (I8c803ab08db372802117de4fa4e2a187[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00107_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00107_00003_U (
.fgallag_sel( I13ba48a6b360f3cff5f37ce60cb735c6[fgallag_SEL-1:0]),
.fgallag( fgallag_00107_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00107_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00107_00003 };

assign fgallag_final_00107_00003 = (I13ba48a6b360f3cff5f37ce60cb735c6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00107_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00107_00004_U (
.fgallag_sel( I4547cd1dad45dfd01e335e8cf20eadd6[fgallag_SEL-1:0]),
.fgallag( fgallag_00107_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00107_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00107_00004 };

assign fgallag_final_00107_00004 = (I4547cd1dad45dfd01e335e8cf20eadd6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00107_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00108_00000_U (
.fgallag_sel( I0a305655b815b0cc159ac1c5f4ce30f8[fgallag_SEL-1:0]),
.fgallag( fgallag_00108_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00108_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00108_00000 };

assign fgallag_final_00108_00000 = (I0a305655b815b0cc159ac1c5f4ce30f8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00108_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00108_00001_U (
.fgallag_sel( I3633737da6b74284b0ea9a06c3f5875f[fgallag_SEL-1:0]),
.fgallag( fgallag_00108_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00108_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00108_00001 };

assign fgallag_final_00108_00001 = (I3633737da6b74284b0ea9a06c3f5875f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00108_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00108_00002_U (
.fgallag_sel( Ia949c1b338d1cba07cf6bb6572c3e322[fgallag_SEL-1:0]),
.fgallag( fgallag_00108_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00108_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00108_00002 };

assign fgallag_final_00108_00002 = (Ia949c1b338d1cba07cf6bb6572c3e322[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00108_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00109_00000_U (
.fgallag_sel( I9a0185f8400159415bc0ad6c38284041[fgallag_SEL-1:0]),
.fgallag( fgallag_00109_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00109_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00109_00000 };

assign fgallag_final_00109_00000 = (I9a0185f8400159415bc0ad6c38284041[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00109_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00109_00001_U (
.fgallag_sel( I3eeffe43e7deed7ee77a7f5a3bce3cd2[fgallag_SEL-1:0]),
.fgallag( fgallag_00109_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00109_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00109_00001 };

assign fgallag_final_00109_00001 = (I3eeffe43e7deed7ee77a7f5a3bce3cd2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00109_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00109_00002_U (
.fgallag_sel( I85af0c31ca7002ae569d9f5ce39943f7[fgallag_SEL-1:0]),
.fgallag( fgallag_00109_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00109_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00109_00002 };

assign fgallag_final_00109_00002 = (I85af0c31ca7002ae569d9f5ce39943f7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00109_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00110_00000_U (
.fgallag_sel( I3dfb8d2fad83fbd807fbfc6330c5b857[fgallag_SEL-1:0]),
.fgallag( fgallag_00110_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00110_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00110_00000 };

assign fgallag_final_00110_00000 = (I3dfb8d2fad83fbd807fbfc6330c5b857[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00110_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00110_00001_U (
.fgallag_sel( Ic12be21bcba5fa49437cc44dd8a7f064[fgallag_SEL-1:0]),
.fgallag( fgallag_00110_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00110_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00110_00001 };

assign fgallag_final_00110_00001 = (Ic12be21bcba5fa49437cc44dd8a7f064[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00110_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00110_00002_U (
.fgallag_sel( I713a384d022d3012e3d0019f5c4ac077[fgallag_SEL-1:0]),
.fgallag( fgallag_00110_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00110_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00110_00002 };

assign fgallag_final_00110_00002 = (I713a384d022d3012e3d0019f5c4ac077[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00110_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00111_00000_U (
.fgallag_sel( I80550019479d0323d0dd7e7d0f767d83[fgallag_SEL-1:0]),
.fgallag( fgallag_00111_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00111_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00111_00000 };

assign fgallag_final_00111_00000 = (I80550019479d0323d0dd7e7d0f767d83[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00111_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00111_00001_U (
.fgallag_sel( Ib8a866f080dd997e0b6c93b6c844d1bc[fgallag_SEL-1:0]),
.fgallag( fgallag_00111_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00111_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00111_00001 };

assign fgallag_final_00111_00001 = (Ib8a866f080dd997e0b6c93b6c844d1bc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00111_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00111_00002_U (
.fgallag_sel( Id542de206d736ee3769ea0bd037cb627[fgallag_SEL-1:0]),
.fgallag( fgallag_00111_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00111_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00111_00002 };

assign fgallag_final_00111_00002 = (Id542de206d736ee3769ea0bd037cb627[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00111_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00112_00000_U (
.fgallag_sel( I77e6cdb09c92492c3303d0213de9c291[fgallag_SEL-1:0]),
.fgallag( fgallag_00112_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00112_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00112_00000 };

assign fgallag_final_00112_00000 = (I77e6cdb09c92492c3303d0213de9c291[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00112_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00112_00001_U (
.fgallag_sel( I788c33a9f94b26f4ce0f515891d06f90[fgallag_SEL-1:0]),
.fgallag( fgallag_00112_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00112_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00112_00001 };

assign fgallag_final_00112_00001 = (I788c33a9f94b26f4ce0f515891d06f90[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00112_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00112_00002_U (
.fgallag_sel( Iaf7074c2b570a296fe2ea8a5a7097ca0[fgallag_SEL-1:0]),
.fgallag( fgallag_00112_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00112_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00112_00002 };

assign fgallag_final_00112_00002 = (Iaf7074c2b570a296fe2ea8a5a7097ca0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00112_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00112_00003_U (
.fgallag_sel( I8964c6d3f8e02866a6ad86553ab05d99[fgallag_SEL-1:0]),
.fgallag( fgallag_00112_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00112_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00112_00003 };

assign fgallag_final_00112_00003 = (I8964c6d3f8e02866a6ad86553ab05d99[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00112_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00113_00000_U (
.fgallag_sel( I2aa25edaca90c9dae8ed63b48d333c17[fgallag_SEL-1:0]),
.fgallag( fgallag_00113_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00113_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00113_00000 };

assign fgallag_final_00113_00000 = (I2aa25edaca90c9dae8ed63b48d333c17[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00113_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00113_00001_U (
.fgallag_sel( I51a440917c7ae23339bec6f8a745c103[fgallag_SEL-1:0]),
.fgallag( fgallag_00113_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00113_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00113_00001 };

assign fgallag_final_00113_00001 = (I51a440917c7ae23339bec6f8a745c103[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00113_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00113_00002_U (
.fgallag_sel( I56ce875e4619d4d8d6ca2fa0ddee91b1[fgallag_SEL-1:0]),
.fgallag( fgallag_00113_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00113_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00113_00002 };

assign fgallag_final_00113_00002 = (I56ce875e4619d4d8d6ca2fa0ddee91b1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00113_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00113_00003_U (
.fgallag_sel( I80607da8f92f5a5d2e4798a62a7b1c5c[fgallag_SEL-1:0]),
.fgallag( fgallag_00113_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00113_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00113_00003 };

assign fgallag_final_00113_00003 = (I80607da8f92f5a5d2e4798a62a7b1c5c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00113_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00114_00000_U (
.fgallag_sel( Ic4dcaa520e26bac40b3876f02074f856[fgallag_SEL-1:0]),
.fgallag( fgallag_00114_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00114_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00114_00000 };

assign fgallag_final_00114_00000 = (Ic4dcaa520e26bac40b3876f02074f856[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00114_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00114_00001_U (
.fgallag_sel( I3b2714d34081a3b6cccc47fa1638e72e[fgallag_SEL-1:0]),
.fgallag( fgallag_00114_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00114_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00114_00001 };

assign fgallag_final_00114_00001 = (I3b2714d34081a3b6cccc47fa1638e72e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00114_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00114_00002_U (
.fgallag_sel( I2db1d1ee8f546c00e512875ce2e13cee[fgallag_SEL-1:0]),
.fgallag( fgallag_00114_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00114_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00114_00002 };

assign fgallag_final_00114_00002 = (I2db1d1ee8f546c00e512875ce2e13cee[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00114_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00114_00003_U (
.fgallag_sel( If80a6bb104ff3b2020e909103c104063[fgallag_SEL-1:0]),
.fgallag( fgallag_00114_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00114_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00114_00003 };

assign fgallag_final_00114_00003 = (If80a6bb104ff3b2020e909103c104063[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00114_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00115_00000_U (
.fgallag_sel( Iadb72cc5444816fbd132256493930bb4[fgallag_SEL-1:0]),
.fgallag( fgallag_00115_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00115_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00115_00000 };

assign fgallag_final_00115_00000 = (Iadb72cc5444816fbd132256493930bb4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00115_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00115_00001_U (
.fgallag_sel( I3a8ec1ad07bfada3d2c6ffca88b8b678[fgallag_SEL-1:0]),
.fgallag( fgallag_00115_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00115_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00115_00001 };

assign fgallag_final_00115_00001 = (I3a8ec1ad07bfada3d2c6ffca88b8b678[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00115_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00115_00002_U (
.fgallag_sel( I0aa042b86d9f68d22a49b4eb480a9088[fgallag_SEL-1:0]),
.fgallag( fgallag_00115_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00115_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00115_00002 };

assign fgallag_final_00115_00002 = (I0aa042b86d9f68d22a49b4eb480a9088[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00115_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00115_00003_U (
.fgallag_sel( I89a387374771b68d87d7ff2dcc810829[fgallag_SEL-1:0]),
.fgallag( fgallag_00115_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00115_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00115_00003 };

assign fgallag_final_00115_00003 = (I89a387374771b68d87d7ff2dcc810829[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00115_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00116_00000_U (
.fgallag_sel( I2935b3d5c3bba4dddfc7ae03fa77b229[fgallag_SEL-1:0]),
.fgallag( fgallag_00116_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00116_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00116_00000 };

assign fgallag_final_00116_00000 = (I2935b3d5c3bba4dddfc7ae03fa77b229[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00116_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00116_00001_U (
.fgallag_sel( I4e0c0248f4aa97d263d64dfec36e3aa2[fgallag_SEL-1:0]),
.fgallag( fgallag_00116_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00116_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00116_00001 };

assign fgallag_final_00116_00001 = (I4e0c0248f4aa97d263d64dfec36e3aa2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00116_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00116_00002_U (
.fgallag_sel( Ia2871d7493b2727d2cb2fbab596b7e6a[fgallag_SEL-1:0]),
.fgallag( fgallag_00116_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00116_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00116_00002 };

assign fgallag_final_00116_00002 = (Ia2871d7493b2727d2cb2fbab596b7e6a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00116_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00117_00000_U (
.fgallag_sel( Ie57adae8873946d6c706074b52a49786[fgallag_SEL-1:0]),
.fgallag( fgallag_00117_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00117_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00117_00000 };

assign fgallag_final_00117_00000 = (Ie57adae8873946d6c706074b52a49786[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00117_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00117_00001_U (
.fgallag_sel( If5ac85646e4b339a19af658f01d0a17f[fgallag_SEL-1:0]),
.fgallag( fgallag_00117_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00117_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00117_00001 };

assign fgallag_final_00117_00001 = (If5ac85646e4b339a19af658f01d0a17f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00117_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00117_00002_U (
.fgallag_sel( I1c092426f34be030b3e020f40517b0e1[fgallag_SEL-1:0]),
.fgallag( fgallag_00117_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00117_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00117_00002 };

assign fgallag_final_00117_00002 = (I1c092426f34be030b3e020f40517b0e1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00117_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00118_00000_U (
.fgallag_sel( Ic719b72ad271bc7c077067518e6bbb98[fgallag_SEL-1:0]),
.fgallag( fgallag_00118_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00118_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00118_00000 };

assign fgallag_final_00118_00000 = (Ic719b72ad271bc7c077067518e6bbb98[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00118_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00118_00001_U (
.fgallag_sel( Ib87362230682c88d68a0ba70e25f3c20[fgallag_SEL-1:0]),
.fgallag( fgallag_00118_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00118_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00118_00001 };

assign fgallag_final_00118_00001 = (Ib87362230682c88d68a0ba70e25f3c20[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00118_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00118_00002_U (
.fgallag_sel( Ifcf097a102f8dc1f912022fed893d222[fgallag_SEL-1:0]),
.fgallag( fgallag_00118_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00118_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00118_00002 };

assign fgallag_final_00118_00002 = (Ifcf097a102f8dc1f912022fed893d222[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00118_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00119_00000_U (
.fgallag_sel( I56483ca3fa550dc59bfa347780cfef7b[fgallag_SEL-1:0]),
.fgallag( fgallag_00119_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00119_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00119_00000 };

assign fgallag_final_00119_00000 = (I56483ca3fa550dc59bfa347780cfef7b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00119_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00119_00001_U (
.fgallag_sel( I4aa9f61be376458185c3235442c8fda0[fgallag_SEL-1:0]),
.fgallag( fgallag_00119_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00119_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00119_00001 };

assign fgallag_final_00119_00001 = (I4aa9f61be376458185c3235442c8fda0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00119_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00119_00002_U (
.fgallag_sel( Id91fde1007d47258273299de80721390[fgallag_SEL-1:0]),
.fgallag( fgallag_00119_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00119_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00119_00002 };

assign fgallag_final_00119_00002 = (Id91fde1007d47258273299de80721390[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00119_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00120_00000_U (
.fgallag_sel( Id58498c34aff2e1216c189b9df88822c[fgallag_SEL-1:0]),
.fgallag( fgallag_00120_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00120_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00120_00000 };

assign fgallag_final_00120_00000 = (Id58498c34aff2e1216c189b9df88822c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00120_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00120_00001_U (
.fgallag_sel( Ib52e0c68caadcf4dd9636a84f5460e53[fgallag_SEL-1:0]),
.fgallag( fgallag_00120_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00120_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00120_00001 };

assign fgallag_final_00120_00001 = (Ib52e0c68caadcf4dd9636a84f5460e53[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00120_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00120_00002_U (
.fgallag_sel( Ie19679053b289bb5a0aad570cc81bd14[fgallag_SEL-1:0]),
.fgallag( fgallag_00120_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00120_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00120_00002 };

assign fgallag_final_00120_00002 = (Ie19679053b289bb5a0aad570cc81bd14[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00120_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00120_00003_U (
.fgallag_sel( I8862c5ef45b723c9abf5d0ab6854a900[fgallag_SEL-1:0]),
.fgallag( fgallag_00120_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00120_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00120_00003 };

assign fgallag_final_00120_00003 = (I8862c5ef45b723c9abf5d0ab6854a900[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00120_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00120_00004_U (
.fgallag_sel( I30db951a07af96a8ddf59360141b9a6a[fgallag_SEL-1:0]),
.fgallag( fgallag_00120_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00120_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00120_00004 };

assign fgallag_final_00120_00004 = (I30db951a07af96a8ddf59360141b9a6a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00120_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00121_00000_U (
.fgallag_sel( I4855a0a0c6426d33014ce6a4c96965ce[fgallag_SEL-1:0]),
.fgallag( fgallag_00121_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00121_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00121_00000 };

assign fgallag_final_00121_00000 = (I4855a0a0c6426d33014ce6a4c96965ce[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00121_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00121_00001_U (
.fgallag_sel( I362e8db1791718290bd33a79b4fc0855[fgallag_SEL-1:0]),
.fgallag( fgallag_00121_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00121_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00121_00001 };

assign fgallag_final_00121_00001 = (I362e8db1791718290bd33a79b4fc0855[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00121_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00121_00002_U (
.fgallag_sel( I773f0508440fb71d73fd82a372cc0a00[fgallag_SEL-1:0]),
.fgallag( fgallag_00121_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00121_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00121_00002 };

assign fgallag_final_00121_00002 = (I773f0508440fb71d73fd82a372cc0a00[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00121_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00121_00003_U (
.fgallag_sel( I792891cecae468d7a87e12f2da62a718[fgallag_SEL-1:0]),
.fgallag( fgallag_00121_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00121_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00121_00003 };

assign fgallag_final_00121_00003 = (I792891cecae468d7a87e12f2da62a718[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00121_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00121_00004_U (
.fgallag_sel( I33303820ad094d7a0ab53bca722fc609[fgallag_SEL-1:0]),
.fgallag( fgallag_00121_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00121_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00121_00004 };

assign fgallag_final_00121_00004 = (I33303820ad094d7a0ab53bca722fc609[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00121_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00122_00000_U (
.fgallag_sel( Iff98739de575e25104c0dc30f08912a5[fgallag_SEL-1:0]),
.fgallag( fgallag_00122_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00122_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00122_00000 };

assign fgallag_final_00122_00000 = (Iff98739de575e25104c0dc30f08912a5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00122_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00122_00001_U (
.fgallag_sel( I1952614b64ea451e9d0646dcce5dd1cd[fgallag_SEL-1:0]),
.fgallag( fgallag_00122_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00122_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00122_00001 };

assign fgallag_final_00122_00001 = (I1952614b64ea451e9d0646dcce5dd1cd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00122_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00122_00002_U (
.fgallag_sel( I49c1a7d1c20a25496821ad80c7eff790[fgallag_SEL-1:0]),
.fgallag( fgallag_00122_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00122_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00122_00002 };

assign fgallag_final_00122_00002 = (I49c1a7d1c20a25496821ad80c7eff790[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00122_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00122_00003_U (
.fgallag_sel( Ie2be17a55e79ca76350e033f227800de[fgallag_SEL-1:0]),
.fgallag( fgallag_00122_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00122_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00122_00003 };

assign fgallag_final_00122_00003 = (Ie2be17a55e79ca76350e033f227800de[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00122_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00122_00004_U (
.fgallag_sel( I737a5b06f848cacf0c8da4985c73c66b[fgallag_SEL-1:0]),
.fgallag( fgallag_00122_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00122_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00122_00004 };

assign fgallag_final_00122_00004 = (I737a5b06f848cacf0c8da4985c73c66b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00122_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00123_00000_U (
.fgallag_sel( Iab160609bb21501aa55b662d2010357b[fgallag_SEL-1:0]),
.fgallag( fgallag_00123_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00123_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00123_00000 };

assign fgallag_final_00123_00000 = (Iab160609bb21501aa55b662d2010357b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00123_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00123_00001_U (
.fgallag_sel( Ief74f1a9d4a43ee5c9def7b83369bb21[fgallag_SEL-1:0]),
.fgallag( fgallag_00123_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00123_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00123_00001 };

assign fgallag_final_00123_00001 = (Ief74f1a9d4a43ee5c9def7b83369bb21[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00123_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00123_00002_U (
.fgallag_sel( Id144423f50751e661db3860a8487d004[fgallag_SEL-1:0]),
.fgallag( fgallag_00123_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00123_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00123_00002 };

assign fgallag_final_00123_00002 = (Id144423f50751e661db3860a8487d004[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00123_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00123_00003_U (
.fgallag_sel( I623352a4f6705b21d461d6b32e85c12b[fgallag_SEL-1:0]),
.fgallag( fgallag_00123_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00123_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00123_00003 };

assign fgallag_final_00123_00003 = (I623352a4f6705b21d461d6b32e85c12b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00123_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00123_00004_U (
.fgallag_sel( I28d1dc8dc594977b5058b5bb9f6bfc66[fgallag_SEL-1:0]),
.fgallag( fgallag_00123_00004 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00123_00004 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00123_00004 };

assign fgallag_final_00123_00004 = (I28d1dc8dc594977b5058b5bb9f6bfc66[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00123_00004 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00124_00000_U (
.fgallag_sel( I5371a83bf9d6f334cf8d1c5b082527e9[fgallag_SEL-1:0]),
.fgallag( fgallag_00124_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00124_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00124_00000 };

assign fgallag_final_00124_00000 = (I5371a83bf9d6f334cf8d1c5b082527e9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00124_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00124_00001_U (
.fgallag_sel( If1605d6646fd267e701668a7245b3b44[fgallag_SEL-1:0]),
.fgallag( fgallag_00124_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00124_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00124_00001 };

assign fgallag_final_00124_00001 = (If1605d6646fd267e701668a7245b3b44[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00124_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00124_00002_U (
.fgallag_sel( Idf5eb1ac2c5bd92fa08ed935ae298255[fgallag_SEL-1:0]),
.fgallag( fgallag_00124_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00124_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00124_00002 };

assign fgallag_final_00124_00002 = (Idf5eb1ac2c5bd92fa08ed935ae298255[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00124_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00125_00000_U (
.fgallag_sel( I44ce30330c4d2d6033a0a970dd2bdd68[fgallag_SEL-1:0]),
.fgallag( fgallag_00125_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00125_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00125_00000 };

assign fgallag_final_00125_00000 = (I44ce30330c4d2d6033a0a970dd2bdd68[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00125_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00125_00001_U (
.fgallag_sel( Ic101b8f56ea1e25c6b752583a1b01242[fgallag_SEL-1:0]),
.fgallag( fgallag_00125_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00125_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00125_00001 };

assign fgallag_final_00125_00001 = (Ic101b8f56ea1e25c6b752583a1b01242[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00125_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00125_00002_U (
.fgallag_sel( Ib7cf44e681881e55d2d353280a6319d6[fgallag_SEL-1:0]),
.fgallag( fgallag_00125_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00125_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00125_00002 };

assign fgallag_final_00125_00002 = (Ib7cf44e681881e55d2d353280a6319d6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00125_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00126_00000_U (
.fgallag_sel( I35690f724e964248dbb1e80fb1ea49f8[fgallag_SEL-1:0]),
.fgallag( fgallag_00126_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00126_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00126_00000 };

assign fgallag_final_00126_00000 = (I35690f724e964248dbb1e80fb1ea49f8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00126_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00126_00001_U (
.fgallag_sel( I5affa2759148a6baf5b9f0cd3122348c[fgallag_SEL-1:0]),
.fgallag( fgallag_00126_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00126_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00126_00001 };

assign fgallag_final_00126_00001 = (I5affa2759148a6baf5b9f0cd3122348c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00126_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00126_00002_U (
.fgallag_sel( Iaeea1f06ff0c6e9cfa43ba14420c3adc[fgallag_SEL-1:0]),
.fgallag( fgallag_00126_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00126_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00126_00002 };

assign fgallag_final_00126_00002 = (Iaeea1f06ff0c6e9cfa43ba14420c3adc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00126_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00127_00000_U (
.fgallag_sel( Iac5a23266c3b038b4b54a916dccdf3a8[fgallag_SEL-1:0]),
.fgallag( fgallag_00127_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00127_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00127_00000 };

assign fgallag_final_00127_00000 = (Iac5a23266c3b038b4b54a916dccdf3a8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00127_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00127_00001_U (
.fgallag_sel( Icdfb7f52cc27b1cfcde90a100d29af13[fgallag_SEL-1:0]),
.fgallag( fgallag_00127_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00127_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00127_00001 };

assign fgallag_final_00127_00001 = (Icdfb7f52cc27b1cfcde90a100d29af13[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00127_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00127_00002_U (
.fgallag_sel( I71484d7e00efa02a08b54a1405f2902c[fgallag_SEL-1:0]),
.fgallag( fgallag_00127_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00127_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00127_00002 };

assign fgallag_final_00127_00002 = (I71484d7e00efa02a08b54a1405f2902c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00127_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00128_00000_U (
.fgallag_sel( I68a9b0607e69e8b3dae64689eb288a33[fgallag_SEL-1:0]),
.fgallag( fgallag_00128_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00128_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00128_00000 };

assign fgallag_final_00128_00000 = (I68a9b0607e69e8b3dae64689eb288a33[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00128_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00128_00001_U (
.fgallag_sel( I2598c48aad48072a7f216b2ab56ee532[fgallag_SEL-1:0]),
.fgallag( fgallag_00128_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00128_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00128_00001 };

assign fgallag_final_00128_00001 = (I2598c48aad48072a7f216b2ab56ee532[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00128_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00128_00002_U (
.fgallag_sel( I796e3a193b1b66fa9a04ca60aee11ea1[fgallag_SEL-1:0]),
.fgallag( fgallag_00128_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00128_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00128_00002 };

assign fgallag_final_00128_00002 = (I796e3a193b1b66fa9a04ca60aee11ea1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00128_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00128_00003_U (
.fgallag_sel( Ic96be7e69faf0f43b92618131cf0c98a[fgallag_SEL-1:0]),
.fgallag( fgallag_00128_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00128_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00128_00003 };

assign fgallag_final_00128_00003 = (Ic96be7e69faf0f43b92618131cf0c98a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00128_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00129_00000_U (
.fgallag_sel( I648afe4114ce435bf1d13e0ad54425cf[fgallag_SEL-1:0]),
.fgallag( fgallag_00129_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00129_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00129_00000 };

assign fgallag_final_00129_00000 = (I648afe4114ce435bf1d13e0ad54425cf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00129_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00129_00001_U (
.fgallag_sel( If05d7e30b4717e0a1bfd20b90d0539bd[fgallag_SEL-1:0]),
.fgallag( fgallag_00129_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00129_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00129_00001 };

assign fgallag_final_00129_00001 = (If05d7e30b4717e0a1bfd20b90d0539bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00129_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00129_00002_U (
.fgallag_sel( I5fc356af8a62a1d739cb375fb851e90f[fgallag_SEL-1:0]),
.fgallag( fgallag_00129_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00129_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00129_00002 };

assign fgallag_final_00129_00002 = (I5fc356af8a62a1d739cb375fb851e90f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00129_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00129_00003_U (
.fgallag_sel( I22f4c5403fbe33d18f97cf21786cdd80[fgallag_SEL-1:0]),
.fgallag( fgallag_00129_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00129_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00129_00003 };

assign fgallag_final_00129_00003 = (I22f4c5403fbe33d18f97cf21786cdd80[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00129_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00130_00000_U (
.fgallag_sel( I9a1b2b9f924099f1e57fa501ba2e33ba[fgallag_SEL-1:0]),
.fgallag( fgallag_00130_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00130_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00130_00000 };

assign fgallag_final_00130_00000 = (I9a1b2b9f924099f1e57fa501ba2e33ba[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00130_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00130_00001_U (
.fgallag_sel( If6253af4ebc430e4937269a5f4989b29[fgallag_SEL-1:0]),
.fgallag( fgallag_00130_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00130_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00130_00001 };

assign fgallag_final_00130_00001 = (If6253af4ebc430e4937269a5f4989b29[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00130_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00130_00002_U (
.fgallag_sel( I0427d17423548dbb33cf792883b4be8c[fgallag_SEL-1:0]),
.fgallag( fgallag_00130_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00130_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00130_00002 };

assign fgallag_final_00130_00002 = (I0427d17423548dbb33cf792883b4be8c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00130_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00130_00003_U (
.fgallag_sel( Ie539faf01ae85253e399308fef98afd6[fgallag_SEL-1:0]),
.fgallag( fgallag_00130_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00130_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00130_00003 };

assign fgallag_final_00130_00003 = (Ie539faf01ae85253e399308fef98afd6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00130_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00131_00000_U (
.fgallag_sel( Iae6e7c42f250cd9223f18f8830fb177d[fgallag_SEL-1:0]),
.fgallag( fgallag_00131_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00131_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00131_00000 };

assign fgallag_final_00131_00000 = (Iae6e7c42f250cd9223f18f8830fb177d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00131_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00131_00001_U (
.fgallag_sel( Iff47ec1743b59d7f90e9042af7ce44cb[fgallag_SEL-1:0]),
.fgallag( fgallag_00131_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00131_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00131_00001 };

assign fgallag_final_00131_00001 = (Iff47ec1743b59d7f90e9042af7ce44cb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00131_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00131_00002_U (
.fgallag_sel( I1cf4a55ebab332defa32d2922b885285[fgallag_SEL-1:0]),
.fgallag( fgallag_00131_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00131_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00131_00002 };

assign fgallag_final_00131_00002 = (I1cf4a55ebab332defa32d2922b885285[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00131_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00131_00003_U (
.fgallag_sel( I284913858691ad5724073b73a820047a[fgallag_SEL-1:0]),
.fgallag( fgallag_00131_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00131_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00131_00003 };

assign fgallag_final_00131_00003 = (I284913858691ad5724073b73a820047a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00131_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00132_00000_U (
.fgallag_sel( I35626ca53adbbf0a3a71cc6fcf43bcb1[fgallag_SEL-1:0]),
.fgallag( fgallag_00132_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00132_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00132_00000 };

assign fgallag_final_00132_00000 = (I35626ca53adbbf0a3a71cc6fcf43bcb1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00132_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00132_00001_U (
.fgallag_sel( I0d74ef22d31abcec73c7c582310b1e6d[fgallag_SEL-1:0]),
.fgallag( fgallag_00132_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00132_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00132_00001 };

assign fgallag_final_00132_00001 = (I0d74ef22d31abcec73c7c582310b1e6d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00132_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00132_00002_U (
.fgallag_sel( I15f4cf1aa0ad5ce2bda52df338e677e3[fgallag_SEL-1:0]),
.fgallag( fgallag_00132_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00132_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00132_00002 };

assign fgallag_final_00132_00002 = (I15f4cf1aa0ad5ce2bda52df338e677e3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00132_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00132_00003_U (
.fgallag_sel( I6c5ca5e68c8844bb1617a2288b5bbc37[fgallag_SEL-1:0]),
.fgallag( fgallag_00132_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00132_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00132_00003 };

assign fgallag_final_00132_00003 = (I6c5ca5e68c8844bb1617a2288b5bbc37[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00132_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00133_00000_U (
.fgallag_sel( I44343a9491069c3c8ea4fbd6255a5a6c[fgallag_SEL-1:0]),
.fgallag( fgallag_00133_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00133_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00133_00000 };

assign fgallag_final_00133_00000 = (I44343a9491069c3c8ea4fbd6255a5a6c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00133_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00133_00001_U (
.fgallag_sel( I1d8318b94d86e1fd28323a5e5684a37b[fgallag_SEL-1:0]),
.fgallag( fgallag_00133_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00133_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00133_00001 };

assign fgallag_final_00133_00001 = (I1d8318b94d86e1fd28323a5e5684a37b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00133_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00133_00002_U (
.fgallag_sel( I825e83bd88575868f4fcc9a8b8729663[fgallag_SEL-1:0]),
.fgallag( fgallag_00133_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00133_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00133_00002 };

assign fgallag_final_00133_00002 = (I825e83bd88575868f4fcc9a8b8729663[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00133_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00133_00003_U (
.fgallag_sel( I3184a16c71cff80c8c90b40e45f114b8[fgallag_SEL-1:0]),
.fgallag( fgallag_00133_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00133_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00133_00003 };

assign fgallag_final_00133_00003 = (I3184a16c71cff80c8c90b40e45f114b8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00133_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00134_00000_U (
.fgallag_sel( Iae133550f8bad8357a73e7de1372faa3[fgallag_SEL-1:0]),
.fgallag( fgallag_00134_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00134_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00134_00000 };

assign fgallag_final_00134_00000 = (Iae133550f8bad8357a73e7de1372faa3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00134_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00134_00001_U (
.fgallag_sel( Ibccb4a43c410f698e0fff68553326a77[fgallag_SEL-1:0]),
.fgallag( fgallag_00134_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00134_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00134_00001 };

assign fgallag_final_00134_00001 = (Ibccb4a43c410f698e0fff68553326a77[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00134_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00134_00002_U (
.fgallag_sel( I72dc7aa294a3af89101ea62a4223170e[fgallag_SEL-1:0]),
.fgallag( fgallag_00134_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00134_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00134_00002 };

assign fgallag_final_00134_00002 = (I72dc7aa294a3af89101ea62a4223170e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00134_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00134_00003_U (
.fgallag_sel( I91eb3e70921e0b141a344bc57dfbc934[fgallag_SEL-1:0]),
.fgallag( fgallag_00134_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00134_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00134_00003 };

assign fgallag_final_00134_00003 = (I91eb3e70921e0b141a344bc57dfbc934[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00134_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00135_00000_U (
.fgallag_sel( I1986f22f2269cc135c6ed28d35fb0bd1[fgallag_SEL-1:0]),
.fgallag( fgallag_00135_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00135_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00135_00000 };

assign fgallag_final_00135_00000 = (I1986f22f2269cc135c6ed28d35fb0bd1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00135_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00135_00001_U (
.fgallag_sel( Ibef24017bc71de9c002aafa7ce9a784c[fgallag_SEL-1:0]),
.fgallag( fgallag_00135_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00135_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00135_00001 };

assign fgallag_final_00135_00001 = (Ibef24017bc71de9c002aafa7ce9a784c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00135_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00135_00002_U (
.fgallag_sel( Ieae3ed78fa2c45507066f4e20d96e956[fgallag_SEL-1:0]),
.fgallag( fgallag_00135_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00135_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00135_00002 };

assign fgallag_final_00135_00002 = (Ieae3ed78fa2c45507066f4e20d96e956[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00135_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00135_00003_U (
.fgallag_sel( I730fd25ffc7778fd4bb02d33cb3870d6[fgallag_SEL-1:0]),
.fgallag( fgallag_00135_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00135_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00135_00003 };

assign fgallag_final_00135_00003 = (I730fd25ffc7778fd4bb02d33cb3870d6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00135_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00136_00000_U (
.fgallag_sel( I9a32313f2911b797fb0848f7d97e62b9[fgallag_SEL-1:0]),
.fgallag( fgallag_00136_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00136_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00136_00000 };

assign fgallag_final_00136_00000 = (I9a32313f2911b797fb0848f7d97e62b9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00136_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00136_00001_U (
.fgallag_sel( I6373e2d64fdb5dd77733b3e4bb405121[fgallag_SEL-1:0]),
.fgallag( fgallag_00136_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00136_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00136_00001 };

assign fgallag_final_00136_00001 = (I6373e2d64fdb5dd77733b3e4bb405121[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00136_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00136_00002_U (
.fgallag_sel( Ib437aa67ab7c13b45d7a4d56ce9e79b8[fgallag_SEL-1:0]),
.fgallag( fgallag_00136_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00136_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00136_00002 };

assign fgallag_final_00136_00002 = (Ib437aa67ab7c13b45d7a4d56ce9e79b8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00136_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00136_00003_U (
.fgallag_sel( I0cb5c7a759f4c75d4a675f9777f15c5f[fgallag_SEL-1:0]),
.fgallag( fgallag_00136_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00136_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00136_00003 };

assign fgallag_final_00136_00003 = (I0cb5c7a759f4c75d4a675f9777f15c5f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00136_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00137_00000_U (
.fgallag_sel( I0ca91c1426ba14a7b47a081cb3becd19[fgallag_SEL-1:0]),
.fgallag( fgallag_00137_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00137_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00137_00000 };

assign fgallag_final_00137_00000 = (I0ca91c1426ba14a7b47a081cb3becd19[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00137_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00137_00001_U (
.fgallag_sel( I0737e0cc7453e328efab2277bb712ea8[fgallag_SEL-1:0]),
.fgallag( fgallag_00137_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00137_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00137_00001 };

assign fgallag_final_00137_00001 = (I0737e0cc7453e328efab2277bb712ea8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00137_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00137_00002_U (
.fgallag_sel( I456af863661122cc303fccb235f3c7a1[fgallag_SEL-1:0]),
.fgallag( fgallag_00137_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00137_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00137_00002 };

assign fgallag_final_00137_00002 = (I456af863661122cc303fccb235f3c7a1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00137_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00137_00003_U (
.fgallag_sel( Idc5916c4800e9f647d51c52444ab6fff[fgallag_SEL-1:0]),
.fgallag( fgallag_00137_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00137_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00137_00003 };

assign fgallag_final_00137_00003 = (Idc5916c4800e9f647d51c52444ab6fff[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00137_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00138_00000_U (
.fgallag_sel( I57aca70e2b8d126c120736b2606ed333[fgallag_SEL-1:0]),
.fgallag( fgallag_00138_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00138_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00138_00000 };

assign fgallag_final_00138_00000 = (I57aca70e2b8d126c120736b2606ed333[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00138_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00138_00001_U (
.fgallag_sel( Ic6650a6d092b749b4498c08d69cf815e[fgallag_SEL-1:0]),
.fgallag( fgallag_00138_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00138_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00138_00001 };

assign fgallag_final_00138_00001 = (Ic6650a6d092b749b4498c08d69cf815e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00138_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00138_00002_U (
.fgallag_sel( Ic2e3b8f91eb218650c7b9c515c7efe97[fgallag_SEL-1:0]),
.fgallag( fgallag_00138_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00138_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00138_00002 };

assign fgallag_final_00138_00002 = (Ic2e3b8f91eb218650c7b9c515c7efe97[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00138_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00138_00003_U (
.fgallag_sel( I93a084aa1e6881ab8dc905dcdcdfd7ee[fgallag_SEL-1:0]),
.fgallag( fgallag_00138_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00138_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00138_00003 };

assign fgallag_final_00138_00003 = (I93a084aa1e6881ab8dc905dcdcdfd7ee[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00138_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00139_00000_U (
.fgallag_sel( I8cba172573be52c5a90bd40e6f40a508[fgallag_SEL-1:0]),
.fgallag( fgallag_00139_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00139_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00139_00000 };

assign fgallag_final_00139_00000 = (I8cba172573be52c5a90bd40e6f40a508[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00139_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00139_00001_U (
.fgallag_sel( I1cccfd1516af59265731121dde878116[fgallag_SEL-1:0]),
.fgallag( fgallag_00139_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00139_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00139_00001 };

assign fgallag_final_00139_00001 = (I1cccfd1516af59265731121dde878116[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00139_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00139_00002_U (
.fgallag_sel( Ia171bbefe2d20b4c058126c33ef28eb8[fgallag_SEL-1:0]),
.fgallag( fgallag_00139_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00139_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00139_00002 };

assign fgallag_final_00139_00002 = (Ia171bbefe2d20b4c058126c33ef28eb8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00139_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00139_00003_U (
.fgallag_sel( I84bc44a5d53a8f66b985b70c7ec1ae7c[fgallag_SEL-1:0]),
.fgallag( fgallag_00139_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00139_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00139_00003 };

assign fgallag_final_00139_00003 = (I84bc44a5d53a8f66b985b70c7ec1ae7c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00139_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00140_00000_U (
.fgallag_sel( I321b104ca3c818018d4b03adfe1110b9[fgallag_SEL-1:0]),
.fgallag( fgallag_00140_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00140_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00140_00000 };

assign fgallag_final_00140_00000 = (I321b104ca3c818018d4b03adfe1110b9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00140_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00140_00001_U (
.fgallag_sel( Ia79b8994da536c86634bf6f54a21145d[fgallag_SEL-1:0]),
.fgallag( fgallag_00140_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00140_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00140_00001 };

assign fgallag_final_00140_00001 = (Ia79b8994da536c86634bf6f54a21145d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00140_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00140_00002_U (
.fgallag_sel( I4df55ce80eec5fee295b5a0ae92bd6c8[fgallag_SEL-1:0]),
.fgallag( fgallag_00140_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00140_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00140_00002 };

assign fgallag_final_00140_00002 = (I4df55ce80eec5fee295b5a0ae92bd6c8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00140_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00140_00003_U (
.fgallag_sel( I46593a7956590d870fe680228081a6d2[fgallag_SEL-1:0]),
.fgallag( fgallag_00140_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00140_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00140_00003 };

assign fgallag_final_00140_00003 = (I46593a7956590d870fe680228081a6d2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00140_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00141_00000_U (
.fgallag_sel( I906e9da31de73ae45579607a014e8b54[fgallag_SEL-1:0]),
.fgallag( fgallag_00141_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00141_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00141_00000 };

assign fgallag_final_00141_00000 = (I906e9da31de73ae45579607a014e8b54[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00141_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00141_00001_U (
.fgallag_sel( If5dd1a1b9e3fc0e67a85da3183480aed[fgallag_SEL-1:0]),
.fgallag( fgallag_00141_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00141_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00141_00001 };

assign fgallag_final_00141_00001 = (If5dd1a1b9e3fc0e67a85da3183480aed[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00141_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00141_00002_U (
.fgallag_sel( Iadfb1571c78c3f0c05e4ef498267df24[fgallag_SEL-1:0]),
.fgallag( fgallag_00141_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00141_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00141_00002 };

assign fgallag_final_00141_00002 = (Iadfb1571c78c3f0c05e4ef498267df24[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00141_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00141_00003_U (
.fgallag_sel( Icebb43b184c2745cc9da9d01b06bc62f[fgallag_SEL-1:0]),
.fgallag( fgallag_00141_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00141_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00141_00003 };

assign fgallag_final_00141_00003 = (Icebb43b184c2745cc9da9d01b06bc62f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00141_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00142_00000_U (
.fgallag_sel( I6e4b0489ec7333abf2245a1b72a8923d[fgallag_SEL-1:0]),
.fgallag( fgallag_00142_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00142_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00142_00000 };

assign fgallag_final_00142_00000 = (I6e4b0489ec7333abf2245a1b72a8923d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00142_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00142_00001_U (
.fgallag_sel( I24ac5dd30526c1d3bc7b941103a66804[fgallag_SEL-1:0]),
.fgallag( fgallag_00142_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00142_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00142_00001 };

assign fgallag_final_00142_00001 = (I24ac5dd30526c1d3bc7b941103a66804[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00142_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00142_00002_U (
.fgallag_sel( I33681b2292c086fe536dae2aec70903a[fgallag_SEL-1:0]),
.fgallag( fgallag_00142_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00142_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00142_00002 };

assign fgallag_final_00142_00002 = (I33681b2292c086fe536dae2aec70903a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00142_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00142_00003_U (
.fgallag_sel( Ia373ca76c3b15a4148532b3822f82ba5[fgallag_SEL-1:0]),
.fgallag( fgallag_00142_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00142_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00142_00003 };

assign fgallag_final_00142_00003 = (Ia373ca76c3b15a4148532b3822f82ba5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00142_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00143_00000_U (
.fgallag_sel( I7d08adbaf66cea04be4891db610bca3f[fgallag_SEL-1:0]),
.fgallag( fgallag_00143_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00143_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00143_00000 };

assign fgallag_final_00143_00000 = (I7d08adbaf66cea04be4891db610bca3f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00143_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00143_00001_U (
.fgallag_sel( Ic09ed51b20f411683a801eaad61657a3[fgallag_SEL-1:0]),
.fgallag( fgallag_00143_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00143_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00143_00001 };

assign fgallag_final_00143_00001 = (Ic09ed51b20f411683a801eaad61657a3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00143_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00143_00002_U (
.fgallag_sel( I6a9af8c9009b5de47ebe9ee8b79d3831[fgallag_SEL-1:0]),
.fgallag( fgallag_00143_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00143_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00143_00002 };

assign fgallag_final_00143_00002 = (I6a9af8c9009b5de47ebe9ee8b79d3831[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00143_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00143_00003_U (
.fgallag_sel( Ife18e8a16d4437161b75a93e3dff1b5b[fgallag_SEL-1:0]),
.fgallag( fgallag_00143_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00143_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00143_00003 };

assign fgallag_final_00143_00003 = (Ife18e8a16d4437161b75a93e3dff1b5b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00143_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00144_00000_U (
.fgallag_sel( I0cde86532c8db1a32d9fbe38a40b91b8[fgallag_SEL-1:0]),
.fgallag( fgallag_00144_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00144_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00144_00000 };

assign fgallag_final_00144_00000 = (I0cde86532c8db1a32d9fbe38a40b91b8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00144_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00144_00001_U (
.fgallag_sel( I49c8ec4cd33e6caed8ed7dab779e7ebb[fgallag_SEL-1:0]),
.fgallag( fgallag_00144_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00144_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00144_00001 };

assign fgallag_final_00144_00001 = (I49c8ec4cd33e6caed8ed7dab779e7ebb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00144_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00144_00002_U (
.fgallag_sel( Idb86f95570587a0711d796aac7004c25[fgallag_SEL-1:0]),
.fgallag( fgallag_00144_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00144_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00144_00002 };

assign fgallag_final_00144_00002 = (Idb86f95570587a0711d796aac7004c25[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00144_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00144_00003_U (
.fgallag_sel( I2d1373d0b18992fa46a9607a86d21520[fgallag_SEL-1:0]),
.fgallag( fgallag_00144_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00144_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00144_00003 };

assign fgallag_final_00144_00003 = (I2d1373d0b18992fa46a9607a86d21520[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00144_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00145_00000_U (
.fgallag_sel( I30f26e090ab14551cbac41883ad8a152[fgallag_SEL-1:0]),
.fgallag( fgallag_00145_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00145_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00145_00000 };

assign fgallag_final_00145_00000 = (I30f26e090ab14551cbac41883ad8a152[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00145_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00145_00001_U (
.fgallag_sel( Ib1b4e41ab25733d1d6dd54e1fe81a419[fgallag_SEL-1:0]),
.fgallag( fgallag_00145_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00145_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00145_00001 };

assign fgallag_final_00145_00001 = (Ib1b4e41ab25733d1d6dd54e1fe81a419[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00145_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00145_00002_U (
.fgallag_sel( I146c0d5154a6de44c0536de873904ccf[fgallag_SEL-1:0]),
.fgallag( fgallag_00145_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00145_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00145_00002 };

assign fgallag_final_00145_00002 = (I146c0d5154a6de44c0536de873904ccf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00145_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00145_00003_U (
.fgallag_sel( I8eb9d4839a478a4e28b45a549b5682a4[fgallag_SEL-1:0]),
.fgallag( fgallag_00145_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00145_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00145_00003 };

assign fgallag_final_00145_00003 = (I8eb9d4839a478a4e28b45a549b5682a4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00145_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00146_00000_U (
.fgallag_sel( I2501ef991a59512c43693ba9d7db8571[fgallag_SEL-1:0]),
.fgallag( fgallag_00146_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00146_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00146_00000 };

assign fgallag_final_00146_00000 = (I2501ef991a59512c43693ba9d7db8571[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00146_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00146_00001_U (
.fgallag_sel( I38213f78fd4dc52f9d2c9b7b22136c1c[fgallag_SEL-1:0]),
.fgallag( fgallag_00146_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00146_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00146_00001 };

assign fgallag_final_00146_00001 = (I38213f78fd4dc52f9d2c9b7b22136c1c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00146_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00146_00002_U (
.fgallag_sel( I49ce91ac152279af421bbc6c4d9b8087[fgallag_SEL-1:0]),
.fgallag( fgallag_00146_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00146_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00146_00002 };

assign fgallag_final_00146_00002 = (I49ce91ac152279af421bbc6c4d9b8087[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00146_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00146_00003_U (
.fgallag_sel( I6a2b7bb2cb3ca2ab932c211a68dded55[fgallag_SEL-1:0]),
.fgallag( fgallag_00146_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00146_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00146_00003 };

assign fgallag_final_00146_00003 = (I6a2b7bb2cb3ca2ab932c211a68dded55[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00146_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00147_00000_U (
.fgallag_sel( Idaae6ba9da8754615a2c34ef859492db[fgallag_SEL-1:0]),
.fgallag( fgallag_00147_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00147_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00147_00000 };

assign fgallag_final_00147_00000 = (Idaae6ba9da8754615a2c34ef859492db[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00147_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00147_00001_U (
.fgallag_sel( Icaca9fc70a3ec6c48c0e41f8168e2bb9[fgallag_SEL-1:0]),
.fgallag( fgallag_00147_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00147_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00147_00001 };

assign fgallag_final_00147_00001 = (Icaca9fc70a3ec6c48c0e41f8168e2bb9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00147_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00147_00002_U (
.fgallag_sel( I4f69b8ff834c7ab3194bc9390ce0f5f6[fgallag_SEL-1:0]),
.fgallag( fgallag_00147_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00147_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00147_00002 };

assign fgallag_final_00147_00002 = (I4f69b8ff834c7ab3194bc9390ce0f5f6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00147_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00147_00003_U (
.fgallag_sel( I037cb596cd48c5533ed22bc32518d992[fgallag_SEL-1:0]),
.fgallag( fgallag_00147_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00147_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00147_00003 };

assign fgallag_final_00147_00003 = (I037cb596cd48c5533ed22bc32518d992[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00147_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00148_00000_U (
.fgallag_sel( I94a89577951de90edc4f73b281ad7364[fgallag_SEL-1:0]),
.fgallag( fgallag_00148_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00148_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00148_00000 };

assign fgallag_final_00148_00000 = (I94a89577951de90edc4f73b281ad7364[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00148_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00148_00001_U (
.fgallag_sel( Ib7493a1a384aebaa7999ff1fb867fc6b[fgallag_SEL-1:0]),
.fgallag( fgallag_00148_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00148_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00148_00001 };

assign fgallag_final_00148_00001 = (Ib7493a1a384aebaa7999ff1fb867fc6b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00148_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00148_00002_U (
.fgallag_sel( I2ceb9e423696539135c5bae5cc2d8d98[fgallag_SEL-1:0]),
.fgallag( fgallag_00148_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00148_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00148_00002 };

assign fgallag_final_00148_00002 = (I2ceb9e423696539135c5bae5cc2d8d98[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00148_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00149_00000_U (
.fgallag_sel( Ia6bbf236436b2ed22bbaae3b8849de6d[fgallag_SEL-1:0]),
.fgallag( fgallag_00149_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00149_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00149_00000 };

assign fgallag_final_00149_00000 = (Ia6bbf236436b2ed22bbaae3b8849de6d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00149_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00149_00001_U (
.fgallag_sel( I33cdaee4676d546dd5507df4704ea1f8[fgallag_SEL-1:0]),
.fgallag( fgallag_00149_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00149_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00149_00001 };

assign fgallag_final_00149_00001 = (I33cdaee4676d546dd5507df4704ea1f8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00149_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00149_00002_U (
.fgallag_sel( Ia44daa9ddc3e4d377267333813d4675f[fgallag_SEL-1:0]),
.fgallag( fgallag_00149_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00149_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00149_00002 };

assign fgallag_final_00149_00002 = (Ia44daa9ddc3e4d377267333813d4675f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00149_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00150_00000_U (
.fgallag_sel( Ie1f8fff3f43426d6bc39e45322a532ca[fgallag_SEL-1:0]),
.fgallag( fgallag_00150_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00150_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00150_00000 };

assign fgallag_final_00150_00000 = (Ie1f8fff3f43426d6bc39e45322a532ca[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00150_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00150_00001_U (
.fgallag_sel( I4ee181895efc22862b6e85802a944095[fgallag_SEL-1:0]),
.fgallag( fgallag_00150_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00150_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00150_00001 };

assign fgallag_final_00150_00001 = (I4ee181895efc22862b6e85802a944095[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00150_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00150_00002_U (
.fgallag_sel( I5c24ea83cabbb6be089ac084732cb9d6[fgallag_SEL-1:0]),
.fgallag( fgallag_00150_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00150_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00150_00002 };

assign fgallag_final_00150_00002 = (I5c24ea83cabbb6be089ac084732cb9d6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00150_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00151_00000_U (
.fgallag_sel( Ifee2342449a3b3d0036ce2ecbc9ae189[fgallag_SEL-1:0]),
.fgallag( fgallag_00151_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00151_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00151_00000 };

assign fgallag_final_00151_00000 = (Ifee2342449a3b3d0036ce2ecbc9ae189[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00151_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00151_00001_U (
.fgallag_sel( I70a9a9b8f25066612a50e411ad68e6c4[fgallag_SEL-1:0]),
.fgallag( fgallag_00151_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00151_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00151_00001 };

assign fgallag_final_00151_00001 = (I70a9a9b8f25066612a50e411ad68e6c4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00151_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00151_00002_U (
.fgallag_sel( I1870059af857c79d444bef948bb536ef[fgallag_SEL-1:0]),
.fgallag( fgallag_00151_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00151_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00151_00002 };

assign fgallag_final_00151_00002 = (I1870059af857c79d444bef948bb536ef[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00151_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00152_00000_U (
.fgallag_sel( Iafe61ab12e232a1090123a0f16eefaca[fgallag_SEL-1:0]),
.fgallag( fgallag_00152_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00152_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00152_00000 };

assign fgallag_final_00152_00000 = (Iafe61ab12e232a1090123a0f16eefaca[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00152_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00152_00001_U (
.fgallag_sel( I10ca809fe9a04eaf5d7784ba69314178[fgallag_SEL-1:0]),
.fgallag( fgallag_00152_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00152_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00152_00001 };

assign fgallag_final_00152_00001 = (I10ca809fe9a04eaf5d7784ba69314178[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00152_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00152_00002_U (
.fgallag_sel( I7a1bd0a115b3a1f85cb9c54840f5bf9b[fgallag_SEL-1:0]),
.fgallag( fgallag_00152_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00152_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00152_00002 };

assign fgallag_final_00152_00002 = (I7a1bd0a115b3a1f85cb9c54840f5bf9b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00152_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00152_00003_U (
.fgallag_sel( I986a564393d944d7d202414431c6d165[fgallag_SEL-1:0]),
.fgallag( fgallag_00152_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00152_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00152_00003 };

assign fgallag_final_00152_00003 = (I986a564393d944d7d202414431c6d165[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00152_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00153_00000_U (
.fgallag_sel( I464042aaa60a41c7e1faf3d16eeb121d[fgallag_SEL-1:0]),
.fgallag( fgallag_00153_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00153_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00153_00000 };

assign fgallag_final_00153_00000 = (I464042aaa60a41c7e1faf3d16eeb121d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00153_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00153_00001_U (
.fgallag_sel( I34b9a0bf2b6b562fb36291022ddf5179[fgallag_SEL-1:0]),
.fgallag( fgallag_00153_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00153_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00153_00001 };

assign fgallag_final_00153_00001 = (I34b9a0bf2b6b562fb36291022ddf5179[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00153_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00153_00002_U (
.fgallag_sel( I17dd8612b5c7f9dcc90f17e584aab2d3[fgallag_SEL-1:0]),
.fgallag( fgallag_00153_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00153_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00153_00002 };

assign fgallag_final_00153_00002 = (I17dd8612b5c7f9dcc90f17e584aab2d3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00153_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00153_00003_U (
.fgallag_sel( Id77cf7c05844d83e808a694971145261[fgallag_SEL-1:0]),
.fgallag( fgallag_00153_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00153_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00153_00003 };

assign fgallag_final_00153_00003 = (Id77cf7c05844d83e808a694971145261[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00153_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00154_00000_U (
.fgallag_sel( I276c1155d766437253f12b25066b84e4[fgallag_SEL-1:0]),
.fgallag( fgallag_00154_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00154_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00154_00000 };

assign fgallag_final_00154_00000 = (I276c1155d766437253f12b25066b84e4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00154_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00154_00001_U (
.fgallag_sel( Id75b386d8076893cb73baca69c3eff59[fgallag_SEL-1:0]),
.fgallag( fgallag_00154_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00154_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00154_00001 };

assign fgallag_final_00154_00001 = (Id75b386d8076893cb73baca69c3eff59[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00154_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00154_00002_U (
.fgallag_sel( If62ddbe87274965cfd83189c6666401e[fgallag_SEL-1:0]),
.fgallag( fgallag_00154_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00154_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00154_00002 };

assign fgallag_final_00154_00002 = (If62ddbe87274965cfd83189c6666401e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00154_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00154_00003_U (
.fgallag_sel( I4f73a07452638a610b31e3ee52cb5639[fgallag_SEL-1:0]),
.fgallag( fgallag_00154_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00154_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00154_00003 };

assign fgallag_final_00154_00003 = (I4f73a07452638a610b31e3ee52cb5639[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00154_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00155_00000_U (
.fgallag_sel( I2a4faf3344d9bf4ee71da0be8994788a[fgallag_SEL-1:0]),
.fgallag( fgallag_00155_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00155_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00155_00000 };

assign fgallag_final_00155_00000 = (I2a4faf3344d9bf4ee71da0be8994788a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00155_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00155_00001_U (
.fgallag_sel( I7d7ad0cbb962a47e229fe9d8406e6fe1[fgallag_SEL-1:0]),
.fgallag( fgallag_00155_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00155_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00155_00001 };

assign fgallag_final_00155_00001 = (I7d7ad0cbb962a47e229fe9d8406e6fe1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00155_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00155_00002_U (
.fgallag_sel( I82988dc2dc83ac61380d2a5cb6551768[fgallag_SEL-1:0]),
.fgallag( fgallag_00155_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00155_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00155_00002 };

assign fgallag_final_00155_00002 = (I82988dc2dc83ac61380d2a5cb6551768[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00155_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00155_00003_U (
.fgallag_sel( I058c3a9848fd30010e4742d8682081ac[fgallag_SEL-1:0]),
.fgallag( fgallag_00155_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00155_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00155_00003 };

assign fgallag_final_00155_00003 = (I058c3a9848fd30010e4742d8682081ac[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00155_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00156_00000_U (
.fgallag_sel( I368121c2534820a7147858c06e58b3fc[fgallag_SEL-1:0]),
.fgallag( fgallag_00156_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00156_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00156_00000 };

assign fgallag_final_00156_00000 = (I368121c2534820a7147858c06e58b3fc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00156_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00156_00001_U (
.fgallag_sel( I03d4541eeb1440aa72ee490c49977e32[fgallag_SEL-1:0]),
.fgallag( fgallag_00156_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00156_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00156_00001 };

assign fgallag_final_00156_00001 = (I03d4541eeb1440aa72ee490c49977e32[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00156_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00156_00002_U (
.fgallag_sel( I75fdf5a355949a87b768b1e67db674e4[fgallag_SEL-1:0]),
.fgallag( fgallag_00156_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00156_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00156_00002 };

assign fgallag_final_00156_00002 = (I75fdf5a355949a87b768b1e67db674e4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00156_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00156_00003_U (
.fgallag_sel( I088f4a0af0239602d422324549cb9799[fgallag_SEL-1:0]),
.fgallag( fgallag_00156_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00156_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00156_00003 };

assign fgallag_final_00156_00003 = (I088f4a0af0239602d422324549cb9799[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00156_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00157_00000_U (
.fgallag_sel( I787fe66b38237caf805ec14970d154c7[fgallag_SEL-1:0]),
.fgallag( fgallag_00157_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00157_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00157_00000 };

assign fgallag_final_00157_00000 = (I787fe66b38237caf805ec14970d154c7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00157_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00157_00001_U (
.fgallag_sel( Icef176cff3ae503dbbe2af9ecfc4c859[fgallag_SEL-1:0]),
.fgallag( fgallag_00157_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00157_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00157_00001 };

assign fgallag_final_00157_00001 = (Icef176cff3ae503dbbe2af9ecfc4c859[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00157_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00157_00002_U (
.fgallag_sel( Ie0a66e4871bfe94f6716279ecc9ef21c[fgallag_SEL-1:0]),
.fgallag( fgallag_00157_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00157_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00157_00002 };

assign fgallag_final_00157_00002 = (Ie0a66e4871bfe94f6716279ecc9ef21c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00157_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00157_00003_U (
.fgallag_sel( I474adf7a975b405c288058139a08be38[fgallag_SEL-1:0]),
.fgallag( fgallag_00157_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00157_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00157_00003 };

assign fgallag_final_00157_00003 = (I474adf7a975b405c288058139a08be38[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00157_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00158_00000_U (
.fgallag_sel( Iebeadb39658f41dcf8719ed413e46144[fgallag_SEL-1:0]),
.fgallag( fgallag_00158_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00158_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00158_00000 };

assign fgallag_final_00158_00000 = (Iebeadb39658f41dcf8719ed413e46144[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00158_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00158_00001_U (
.fgallag_sel( Ie018b0d9f05a86207ae09ca2efac54e2[fgallag_SEL-1:0]),
.fgallag( fgallag_00158_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00158_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00158_00001 };

assign fgallag_final_00158_00001 = (Ie018b0d9f05a86207ae09ca2efac54e2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00158_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00158_00002_U (
.fgallag_sel( I51ee69807609fca0f332c8bc31afd632[fgallag_SEL-1:0]),
.fgallag( fgallag_00158_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00158_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00158_00002 };

assign fgallag_final_00158_00002 = (I51ee69807609fca0f332c8bc31afd632[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00158_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00158_00003_U (
.fgallag_sel( Iee1cb471704b2a8718a68ef93fd2e356[fgallag_SEL-1:0]),
.fgallag( fgallag_00158_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00158_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00158_00003 };

assign fgallag_final_00158_00003 = (Iee1cb471704b2a8718a68ef93fd2e356[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00158_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00159_00000_U (
.fgallag_sel( I1731c0e3be86eec142c3732ee836e4d5[fgallag_SEL-1:0]),
.fgallag( fgallag_00159_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00159_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00159_00000 };

assign fgallag_final_00159_00000 = (I1731c0e3be86eec142c3732ee836e4d5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00159_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00159_00001_U (
.fgallag_sel( Id3b8c0ca32331f94fd98c8dae72bb15d[fgallag_SEL-1:0]),
.fgallag( fgallag_00159_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00159_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00159_00001 };

assign fgallag_final_00159_00001 = (Id3b8c0ca32331f94fd98c8dae72bb15d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00159_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00159_00002_U (
.fgallag_sel( I6a86b0a82441c6c14436a3e0af6b0fb7[fgallag_SEL-1:0]),
.fgallag( fgallag_00159_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00159_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00159_00002 };

assign fgallag_final_00159_00002 = (I6a86b0a82441c6c14436a3e0af6b0fb7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00159_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00159_00003_U (
.fgallag_sel( I8c92ff598084da7a50f7c68da96620b3[fgallag_SEL-1:0]),
.fgallag( fgallag_00159_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00159_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00159_00003 };

assign fgallag_final_00159_00003 = (I8c92ff598084da7a50f7c68da96620b3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00159_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00160_00000_U (
.fgallag_sel( I8bd1862e7bc2e83e9863389d532e6623[fgallag_SEL-1:0]),
.fgallag( fgallag_00160_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00160_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00160_00000 };

assign fgallag_final_00160_00000 = (I8bd1862e7bc2e83e9863389d532e6623[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00160_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00160_00001_U (
.fgallag_sel( I8053269f8bd78a931878c8350693e1d6[fgallag_SEL-1:0]),
.fgallag( fgallag_00160_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00160_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00160_00001 };

assign fgallag_final_00160_00001 = (I8053269f8bd78a931878c8350693e1d6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00160_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00160_00002_U (
.fgallag_sel( I2ff66cdd7314276232715ef2361ad184[fgallag_SEL-1:0]),
.fgallag( fgallag_00160_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00160_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00160_00002 };

assign fgallag_final_00160_00002 = (I2ff66cdd7314276232715ef2361ad184[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00160_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00160_00003_U (
.fgallag_sel( Icf541c76bfaf37fe6111de037d205f15[fgallag_SEL-1:0]),
.fgallag( fgallag_00160_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00160_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00160_00003 };

assign fgallag_final_00160_00003 = (Icf541c76bfaf37fe6111de037d205f15[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00160_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00161_00000_U (
.fgallag_sel( I68319c8b9febef9f564832429c91b85a[fgallag_SEL-1:0]),
.fgallag( fgallag_00161_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00161_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00161_00000 };

assign fgallag_final_00161_00000 = (I68319c8b9febef9f564832429c91b85a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00161_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00161_00001_U (
.fgallag_sel( I127772614218dd7c50d3136b4f174d7a[fgallag_SEL-1:0]),
.fgallag( fgallag_00161_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00161_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00161_00001 };

assign fgallag_final_00161_00001 = (I127772614218dd7c50d3136b4f174d7a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00161_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00161_00002_U (
.fgallag_sel( Ib8d1aea4ad24c6ceb44f2cc672e1ff90[fgallag_SEL-1:0]),
.fgallag( fgallag_00161_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00161_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00161_00002 };

assign fgallag_final_00161_00002 = (Ib8d1aea4ad24c6ceb44f2cc672e1ff90[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00161_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00161_00003_U (
.fgallag_sel( I9ca26c8104bf15f48b19dc3256914544[fgallag_SEL-1:0]),
.fgallag( fgallag_00161_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00161_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00161_00003 };

assign fgallag_final_00161_00003 = (I9ca26c8104bf15f48b19dc3256914544[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00161_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00162_00000_U (
.fgallag_sel( Icc76d9ffc3f3d7b410205eeb8232a33b[fgallag_SEL-1:0]),
.fgallag( fgallag_00162_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00162_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00162_00000 };

assign fgallag_final_00162_00000 = (Icc76d9ffc3f3d7b410205eeb8232a33b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00162_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00162_00001_U (
.fgallag_sel( I7fc4551d8a0445f79b87b4ba5f2ffeaa[fgallag_SEL-1:0]),
.fgallag( fgallag_00162_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00162_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00162_00001 };

assign fgallag_final_00162_00001 = (I7fc4551d8a0445f79b87b4ba5f2ffeaa[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00162_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00162_00002_U (
.fgallag_sel( I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8[fgallag_SEL-1:0]),
.fgallag( fgallag_00162_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00162_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00162_00002 };

assign fgallag_final_00162_00002 = (I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00162_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00162_00003_U (
.fgallag_sel( Ie34c07af9f6adb9e4b636dce3d0682c0[fgallag_SEL-1:0]),
.fgallag( fgallag_00162_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00162_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00162_00003 };

assign fgallag_final_00162_00003 = (Ie34c07af9f6adb9e4b636dce3d0682c0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00162_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00163_00000_U (
.fgallag_sel( Ib869a349250a765d2f8660e0dbdcf312[fgallag_SEL-1:0]),
.fgallag( fgallag_00163_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00163_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00163_00000 };

assign fgallag_final_00163_00000 = (Ib869a349250a765d2f8660e0dbdcf312[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00163_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00163_00001_U (
.fgallag_sel( I1a4fb631fdc7b5454c266589962ff5f0[fgallag_SEL-1:0]),
.fgallag( fgallag_00163_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00163_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00163_00001 };

assign fgallag_final_00163_00001 = (I1a4fb631fdc7b5454c266589962ff5f0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00163_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00163_00002_U (
.fgallag_sel( I9de4e0e86e9edcf948d9eddf0401b94a[fgallag_SEL-1:0]),
.fgallag( fgallag_00163_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00163_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00163_00002 };

assign fgallag_final_00163_00002 = (I9de4e0e86e9edcf948d9eddf0401b94a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00163_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00163_00003_U (
.fgallag_sel( Iee7b4838986c962969c00a0bbe53ce0b[fgallag_SEL-1:0]),
.fgallag( fgallag_00163_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00163_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00163_00003 };

assign fgallag_final_00163_00003 = (Iee7b4838986c962969c00a0bbe53ce0b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00163_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00164_00000_U (
.fgallag_sel( Id81b11a8ca1dd8989e36cef637ae6aab[fgallag_SEL-1:0]),
.fgallag( fgallag_00164_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00164_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00164_00000 };

assign fgallag_final_00164_00000 = (Id81b11a8ca1dd8989e36cef637ae6aab[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00164_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00164_00001_U (
.fgallag_sel( Ibe96deab015b799fe7f69bae8432952c[fgallag_SEL-1:0]),
.fgallag( fgallag_00164_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00164_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00164_00001 };

assign fgallag_final_00164_00001 = (Ibe96deab015b799fe7f69bae8432952c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00164_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00164_00002_U (
.fgallag_sel( I986b52155cc1470299321a4933241ed7[fgallag_SEL-1:0]),
.fgallag( fgallag_00164_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00164_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00164_00002 };

assign fgallag_final_00164_00002 = (I986b52155cc1470299321a4933241ed7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00164_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00164_00003_U (
.fgallag_sel( I04be63a04f3942ce749cc9bd7540e055[fgallag_SEL-1:0]),
.fgallag( fgallag_00164_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00164_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00164_00003 };

assign fgallag_final_00164_00003 = (I04be63a04f3942ce749cc9bd7540e055[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00164_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00165_00000_U (
.fgallag_sel( Ia7adea5b0ec86e9fcd427a5468d72b64[fgallag_SEL-1:0]),
.fgallag( fgallag_00165_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00165_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00165_00000 };

assign fgallag_final_00165_00000 = (Ia7adea5b0ec86e9fcd427a5468d72b64[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00165_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00165_00001_U (
.fgallag_sel( Ie8990d8abd23f8f9f79d7fe38c57fa8c[fgallag_SEL-1:0]),
.fgallag( fgallag_00165_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00165_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00165_00001 };

assign fgallag_final_00165_00001 = (Ie8990d8abd23f8f9f79d7fe38c57fa8c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00165_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00165_00002_U (
.fgallag_sel( I9d2f90ddddbdbb525d5f070f32546b64[fgallag_SEL-1:0]),
.fgallag( fgallag_00165_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00165_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00165_00002 };

assign fgallag_final_00165_00002 = (I9d2f90ddddbdbb525d5f070f32546b64[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00165_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00165_00003_U (
.fgallag_sel( I905256d73bdb63bf860e15687350795f[fgallag_SEL-1:0]),
.fgallag( fgallag_00165_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00165_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00165_00003 };

assign fgallag_final_00165_00003 = (I905256d73bdb63bf860e15687350795f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00165_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00166_00000_U (
.fgallag_sel( I9adcfc18e4471209edbe9a379e996067[fgallag_SEL-1:0]),
.fgallag( fgallag_00166_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00166_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00166_00000 };

assign fgallag_final_00166_00000 = (I9adcfc18e4471209edbe9a379e996067[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00166_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00166_00001_U (
.fgallag_sel( I3d7d048348bf833f744a9f73889b7802[fgallag_SEL-1:0]),
.fgallag( fgallag_00166_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00166_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00166_00001 };

assign fgallag_final_00166_00001 = (I3d7d048348bf833f744a9f73889b7802[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00166_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00166_00002_U (
.fgallag_sel( Id619e8d4040014d0e415ff71c5e0591f[fgallag_SEL-1:0]),
.fgallag( fgallag_00166_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00166_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00166_00002 };

assign fgallag_final_00166_00002 = (Id619e8d4040014d0e415ff71c5e0591f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00166_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00166_00003_U (
.fgallag_sel( Iaf3de2ef283e03dd72002026e1299224[fgallag_SEL-1:0]),
.fgallag( fgallag_00166_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00166_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00166_00003 };

assign fgallag_final_00166_00003 = (Iaf3de2ef283e03dd72002026e1299224[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00166_00003 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00167_00000_U (
.fgallag_sel( I64551529c0028ec145407be7f5dfef71[fgallag_SEL-1:0]),
.fgallag( fgallag_00167_00000 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00167_00000 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00167_00000 };

assign fgallag_final_00167_00000 = (I64551529c0028ec145407be7f5dfef71[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00167_00000 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00167_00001_U (
.fgallag_sel( I5ebe580a943b65fb16ea722ba101fd05[fgallag_SEL-1:0]),
.fgallag( fgallag_00167_00001 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00167_00001 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00167_00001 };

assign fgallag_final_00167_00001 = (I5ebe580a943b65fb16ea722ba101fd05[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00167_00001 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00167_00002_U (
.fgallag_sel( I0921901599c43b27e701758026dd3ee1[fgallag_SEL-1:0]),
.fgallag( fgallag_00167_00002 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00167_00002 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00167_00002 };

assign fgallag_final_00167_00002 = (I0921901599c43b27e701758026dd3ee1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00167_00002 ;

Ic9c2f173881d25f8976d723957809f51 fgallag_00167_00003_U (
.fgallag_sel( I6033532f27c26b2d42bb3ea128f80dfa[fgallag_SEL-1:0]),
.fgallag( fgallag_00167_00003 ),
.start_in(start_d4 && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign fgallag_full_00167_00003 = { {(MAX_SUM_WDTH_L-fgallag_WDTH){1'b0}}, fgallag_00167_00003 };

assign fgallag_final_00167_00003 = (I6033532f27c26b2d42bb3ea128f80dfa[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : fgallag_full_00167_00003 ;







   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
               conv_qin_00000_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00000_00000  <=  0;
               conv_qin_00000_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00000_00001  <=  0;
               conv_qin_00000_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00000_00002  <=  0;
               conv_qin_00000_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00000_00003  <=  0;
               conv_qin_00000_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00000_00004  <=  0;
               conv_qin_00000_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00000_00005  <=  0;
               conv_qin_00000_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00000_00006  <=  0;
               conv_qin_00000_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00000_00007  <=  0;
               conv_qin_00001_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00001_00000  <=  0;
               conv_qin_00001_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00001_00001  <=  0;
               conv_qin_00001_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00001_00002  <=  0;
               conv_qin_00001_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00001_00003  <=  0;
               conv_qin_00001_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00001_00004  <=  0;
               conv_qin_00001_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00001_00005  <=  0;
               conv_qin_00001_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00001_00006  <=  0;
               conv_qin_00001_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00001_00007  <=  0;
               conv_qin_00002_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00002_00000  <=  0;
               conv_qin_00002_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00002_00001  <=  0;
               conv_qin_00002_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00002_00002  <=  0;
               conv_qin_00002_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00002_00003  <=  0;
               conv_qin_00002_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00002_00004  <=  0;
               conv_qin_00002_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00002_00005  <=  0;
               conv_qin_00002_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00002_00006  <=  0;
               conv_qin_00002_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00002_00007  <=  0;
               conv_qin_00003_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00003_00000  <=  0;
               conv_qin_00003_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00003_00001  <=  0;
               conv_qin_00003_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00003_00002  <=  0;
               conv_qin_00003_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00003_00003  <=  0;
               conv_qin_00003_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00003_00004  <=  0;
               conv_qin_00003_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00003_00005  <=  0;
               conv_qin_00003_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00003_00006  <=  0;
               conv_qin_00003_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00003_00007  <=  0;
               conv_qin_00004_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00004_00000  <=  0;
               conv_qin_00004_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00004_00001  <=  0;
               conv_qin_00004_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00004_00002  <=  0;
               conv_qin_00004_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00004_00003  <=  0;
               conv_qin_00004_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00004_00004  <=  0;
               conv_qin_00004_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00004_00005  <=  0;
               conv_qin_00004_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00004_00006  <=  0;
               conv_qin_00004_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00004_00007  <=  0;
               conv_qin_00004_00008  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00004_00008  <=  0;
               conv_qin_00004_00009  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00004_00009  <=  0;
               conv_qin_00005_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00005_00000  <=  0;
               conv_qin_00005_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00005_00001  <=  0;
               conv_qin_00005_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00005_00002  <=  0;
               conv_qin_00005_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00005_00003  <=  0;
               conv_qin_00005_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00005_00004  <=  0;
               conv_qin_00005_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00005_00005  <=  0;
               conv_qin_00005_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00005_00006  <=  0;
               conv_qin_00005_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00005_00007  <=  0;
               conv_qin_00005_00008  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00005_00008  <=  0;
               conv_qin_00005_00009  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00005_00009  <=  0;
               conv_qin_00006_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00006_00000  <=  0;
               conv_qin_00006_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00006_00001  <=  0;
               conv_qin_00006_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00006_00002  <=  0;
               conv_qin_00006_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00006_00003  <=  0;
               conv_qin_00006_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00006_00004  <=  0;
               conv_qin_00006_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00006_00005  <=  0;
               conv_qin_00006_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00006_00006  <=  0;
               conv_qin_00006_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00006_00007  <=  0;
               conv_qin_00006_00008  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00006_00008  <=  0;
               conv_qin_00006_00009  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00006_00009  <=  0;
               conv_qin_00007_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00007_00000  <=  0;
               conv_qin_00007_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00007_00001  <=  0;
               conv_qin_00007_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00007_00002  <=  0;
               conv_qin_00007_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00007_00003  <=  0;
               conv_qin_00007_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00007_00004  <=  0;
               conv_qin_00007_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00007_00005  <=  0;
               conv_qin_00007_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00007_00006  <=  0;
               conv_qin_00007_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00007_00007  <=  0;
               conv_qin_00007_00008  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00007_00008  <=  0;
               conv_qin_00007_00009  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00007_00009  <=  0;
               conv_qin_00008_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00008_00000  <=  0;
               conv_qin_00008_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00008_00001  <=  0;
               conv_qin_00008_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00008_00002  <=  0;
               conv_qin_00008_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00008_00003  <=  0;
               conv_qin_00008_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00008_00004  <=  0;
               conv_qin_00008_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00008_00005  <=  0;
               conv_qin_00008_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00008_00006  <=  0;
               conv_qin_00008_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00008_00007  <=  0;
               conv_qin_00009_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00009_00000  <=  0;
               conv_qin_00009_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00009_00001  <=  0;
               conv_qin_00009_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00009_00002  <=  0;
               conv_qin_00009_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00009_00003  <=  0;
               conv_qin_00009_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00009_00004  <=  0;
               conv_qin_00009_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00009_00005  <=  0;
               conv_qin_00009_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00009_00006  <=  0;
               conv_qin_00009_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00009_00007  <=  0;
               conv_qin_00010_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00010_00000  <=  0;
               conv_qin_00010_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00010_00001  <=  0;
               conv_qin_00010_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00010_00002  <=  0;
               conv_qin_00010_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00010_00003  <=  0;
               conv_qin_00010_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00010_00004  <=  0;
               conv_qin_00010_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00010_00005  <=  0;
               conv_qin_00010_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00010_00006  <=  0;
               conv_qin_00010_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00010_00007  <=  0;
               conv_qin_00011_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00011_00000  <=  0;
               conv_qin_00011_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00011_00001  <=  0;
               conv_qin_00011_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00011_00002  <=  0;
               conv_qin_00011_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00011_00003  <=  0;
               conv_qin_00011_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00011_00004  <=  0;
               conv_qin_00011_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00011_00005  <=  0;
               conv_qin_00011_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00011_00006  <=  0;
               conv_qin_00011_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00011_00007  <=  0;
               conv_qin_00012_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00012_00000  <=  0;
               conv_qin_00012_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00012_00001  <=  0;
               conv_qin_00012_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00012_00002  <=  0;
               conv_qin_00012_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00012_00003  <=  0;
               conv_qin_00012_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00012_00004  <=  0;
               conv_qin_00012_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00012_00005  <=  0;
               conv_qin_00012_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00012_00006  <=  0;
               conv_qin_00012_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00012_00007  <=  0;
               conv_qin_00012_00008  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00012_00008  <=  0;
               conv_qin_00012_00009  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00012_00009  <=  0;
               conv_qin_00013_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00013_00000  <=  0;
               conv_qin_00013_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00013_00001  <=  0;
               conv_qin_00013_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00013_00002  <=  0;
               conv_qin_00013_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00013_00003  <=  0;
               conv_qin_00013_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00013_00004  <=  0;
               conv_qin_00013_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00013_00005  <=  0;
               conv_qin_00013_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00013_00006  <=  0;
               conv_qin_00013_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00013_00007  <=  0;
               conv_qin_00013_00008  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00013_00008  <=  0;
               conv_qin_00013_00009  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00013_00009  <=  0;
               conv_qin_00014_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00014_00000  <=  0;
               conv_qin_00014_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00014_00001  <=  0;
               conv_qin_00014_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00014_00002  <=  0;
               conv_qin_00014_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00014_00003  <=  0;
               conv_qin_00014_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00014_00004  <=  0;
               conv_qin_00014_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00014_00005  <=  0;
               conv_qin_00014_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00014_00006  <=  0;
               conv_qin_00014_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00014_00007  <=  0;
               conv_qin_00014_00008  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00014_00008  <=  0;
               conv_qin_00014_00009  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00014_00009  <=  0;
               conv_qin_00015_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00015_00000  <=  0;
               conv_qin_00015_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00015_00001  <=  0;
               conv_qin_00015_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00015_00002  <=  0;
               conv_qin_00015_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00015_00003  <=  0;
               conv_qin_00015_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00015_00004  <=  0;
               conv_qin_00015_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00015_00005  <=  0;
               conv_qin_00015_00006  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00015_00006  <=  0;
               conv_qin_00015_00007  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00015_00007  <=  0;
               conv_qin_00015_00008  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00015_00008  <=  0;
               conv_qin_00015_00009  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00015_00009  <=  0;
               conv_qin_00016_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00016_00000  <=  0;
               conv_qin_00016_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00016_00001  <=  0;
               conv_qin_00016_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00016_00002  <=  0;
               conv_qin_00016_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00016_00003  <=  0;
               conv_qin_00017_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00017_00000  <=  0;
               conv_qin_00017_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00017_00001  <=  0;
               conv_qin_00017_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00017_00002  <=  0;
               conv_qin_00017_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00017_00003  <=  0;
               conv_qin_00018_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00018_00000  <=  0;
               conv_qin_00018_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00018_00001  <=  0;
               conv_qin_00018_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00018_00002  <=  0;
               conv_qin_00018_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00018_00003  <=  0;
               conv_qin_00019_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00019_00000  <=  0;
               conv_qin_00019_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00019_00001  <=  0;
               conv_qin_00019_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00019_00002  <=  0;
               conv_qin_00019_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00019_00003  <=  0;
               conv_qin_00020_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00020_00000  <=  0;
               conv_qin_00020_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00020_00001  <=  0;
               conv_qin_00020_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00020_00002  <=  0;
               conv_qin_00020_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00020_00003  <=  0;
               conv_qin_00020_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00020_00004  <=  0;
               conv_qin_00020_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00020_00005  <=  0;
               conv_qin_00021_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00021_00000  <=  0;
               conv_qin_00021_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00021_00001  <=  0;
               conv_qin_00021_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00021_00002  <=  0;
               conv_qin_00021_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00021_00003  <=  0;
               conv_qin_00021_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00021_00004  <=  0;
               conv_qin_00021_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00021_00005  <=  0;
               conv_qin_00022_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00022_00000  <=  0;
               conv_qin_00022_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00022_00001  <=  0;
               conv_qin_00022_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00022_00002  <=  0;
               conv_qin_00022_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00022_00003  <=  0;
               conv_qin_00022_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00022_00004  <=  0;
               conv_qin_00022_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00022_00005  <=  0;
               conv_qin_00023_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00023_00000  <=  0;
               conv_qin_00023_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00023_00001  <=  0;
               conv_qin_00023_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00023_00002  <=  0;
               conv_qin_00023_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00023_00003  <=  0;
               conv_qin_00023_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00023_00004  <=  0;
               conv_qin_00023_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00023_00005  <=  0;
               conv_qin_00024_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00024_00000  <=  0;
               conv_qin_00024_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00024_00001  <=  0;
               conv_qin_00024_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00024_00002  <=  0;
               conv_qin_00024_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00024_00003  <=  0;
               conv_qin_00024_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00024_00004  <=  0;
               conv_qin_00024_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00024_00005  <=  0;
               conv_qin_00025_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00025_00000  <=  0;
               conv_qin_00025_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00025_00001  <=  0;
               conv_qin_00025_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00025_00002  <=  0;
               conv_qin_00025_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00025_00003  <=  0;
               conv_qin_00025_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00025_00004  <=  0;
               conv_qin_00025_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00025_00005  <=  0;
               conv_qin_00026_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00026_00000  <=  0;
               conv_qin_00026_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00026_00001  <=  0;
               conv_qin_00026_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00026_00002  <=  0;
               conv_qin_00026_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00026_00003  <=  0;
               conv_qin_00026_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00026_00004  <=  0;
               conv_qin_00026_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00026_00005  <=  0;
               conv_qin_00027_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00027_00000  <=  0;
               conv_qin_00027_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00027_00001  <=  0;
               conv_qin_00027_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00027_00002  <=  0;
               conv_qin_00027_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00027_00003  <=  0;
               conv_qin_00027_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00027_00004  <=  0;
               conv_qin_00027_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00027_00005  <=  0;
               conv_qin_00028_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00028_00000  <=  0;
               conv_qin_00028_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00028_00001  <=  0;
               conv_qin_00028_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00028_00002  <=  0;
               conv_qin_00028_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00028_00003  <=  0;
               conv_qin_00028_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00028_00004  <=  0;
               conv_qin_00028_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00028_00005  <=  0;
               conv_qin_00029_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00029_00000  <=  0;
               conv_qin_00029_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00029_00001  <=  0;
               conv_qin_00029_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00029_00002  <=  0;
               conv_qin_00029_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00029_00003  <=  0;
               conv_qin_00029_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00029_00004  <=  0;
               conv_qin_00029_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00029_00005  <=  0;
               conv_qin_00030_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00030_00000  <=  0;
               conv_qin_00030_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00030_00001  <=  0;
               conv_qin_00030_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00030_00002  <=  0;
               conv_qin_00030_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00030_00003  <=  0;
               conv_qin_00030_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00030_00004  <=  0;
               conv_qin_00030_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00030_00005  <=  0;
               conv_qin_00031_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00031_00000  <=  0;
               conv_qin_00031_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00031_00001  <=  0;
               conv_qin_00031_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00031_00002  <=  0;
               conv_qin_00031_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00031_00003  <=  0;
               conv_qin_00031_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00031_00004  <=  0;
               conv_qin_00031_00005  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00031_00005  <=  0;
               conv_qin_00032_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00032_00000  <=  0;
               conv_qin_00032_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00032_00001  <=  0;
               conv_qin_00032_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00032_00002  <=  0;
               conv_qin_00032_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00032_00003  <=  0;
               conv_qin_00033_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00033_00000  <=  0;
               conv_qin_00033_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00033_00001  <=  0;
               conv_qin_00033_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00033_00002  <=  0;
               conv_qin_00033_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00033_00003  <=  0;
               conv_qin_00034_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00034_00000  <=  0;
               conv_qin_00034_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00034_00001  <=  0;
               conv_qin_00034_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00034_00002  <=  0;
               conv_qin_00034_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00034_00003  <=  0;
               conv_qin_00035_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00035_00000  <=  0;
               conv_qin_00035_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00035_00001  <=  0;
               conv_qin_00035_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00035_00002  <=  0;
               conv_qin_00035_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00035_00003  <=  0;
               conv_qin_00036_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00036_00000  <=  0;
               conv_qin_00036_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00036_00001  <=  0;
               conv_qin_00036_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00036_00002  <=  0;
               conv_qin_00036_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00036_00003  <=  0;
               conv_qin_00036_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00036_00004  <=  0;
               conv_qin_00037_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00037_00000  <=  0;
               conv_qin_00037_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00037_00001  <=  0;
               conv_qin_00037_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00037_00002  <=  0;
               conv_qin_00037_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00037_00003  <=  0;
               conv_qin_00037_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00037_00004  <=  0;
               conv_qin_00038_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00038_00000  <=  0;
               conv_qin_00038_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00038_00001  <=  0;
               conv_qin_00038_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00038_00002  <=  0;
               conv_qin_00038_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00038_00003  <=  0;
               conv_qin_00038_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00038_00004  <=  0;
               conv_qin_00039_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00039_00000  <=  0;
               conv_qin_00039_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00039_00001  <=  0;
               conv_qin_00039_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00039_00002  <=  0;
               conv_qin_00039_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00039_00003  <=  0;
               conv_qin_00039_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00039_00004  <=  0;
               conv_qin_00040_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00040_00000  <=  0;
               conv_qin_00040_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00040_00001  <=  0;
               conv_qin_00040_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00040_00002  <=  0;
               conv_qin_00040_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00040_00003  <=  0;
               conv_qin_00040_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00040_00004  <=  0;
               conv_qin_00041_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00041_00000  <=  0;
               conv_qin_00041_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00041_00001  <=  0;
               conv_qin_00041_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00041_00002  <=  0;
               conv_qin_00041_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00041_00003  <=  0;
               conv_qin_00041_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00041_00004  <=  0;
               conv_qin_00042_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00042_00000  <=  0;
               conv_qin_00042_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00042_00001  <=  0;
               conv_qin_00042_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00042_00002  <=  0;
               conv_qin_00042_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00042_00003  <=  0;
               conv_qin_00042_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00042_00004  <=  0;
               conv_qin_00043_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00043_00000  <=  0;
               conv_qin_00043_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00043_00001  <=  0;
               conv_qin_00043_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00043_00002  <=  0;
               conv_qin_00043_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00043_00003  <=  0;
               conv_qin_00043_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00043_00004  <=  0;
               conv_qin_00044_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00044_00000  <=  0;
               conv_qin_00044_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00044_00001  <=  0;
               conv_qin_00044_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00044_00002  <=  0;
               conv_qin_00044_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00044_00003  <=  0;
               conv_qin_00044_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00044_00004  <=  0;
               conv_qin_00045_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00045_00000  <=  0;
               conv_qin_00045_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00045_00001  <=  0;
               conv_qin_00045_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00045_00002  <=  0;
               conv_qin_00045_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00045_00003  <=  0;
               conv_qin_00045_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00045_00004  <=  0;
               conv_qin_00046_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00046_00000  <=  0;
               conv_qin_00046_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00046_00001  <=  0;
               conv_qin_00046_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00046_00002  <=  0;
               conv_qin_00046_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00046_00003  <=  0;
               conv_qin_00046_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00046_00004  <=  0;
               conv_qin_00047_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00047_00000  <=  0;
               conv_qin_00047_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00047_00001  <=  0;
               conv_qin_00047_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00047_00002  <=  0;
               conv_qin_00047_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00047_00003  <=  0;
               conv_qin_00047_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00047_00004  <=  0;
               conv_qin_00048_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00048_00000  <=  0;
               conv_qin_00048_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00048_00001  <=  0;
               conv_qin_00048_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00048_00002  <=  0;
               conv_qin_00048_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00048_00003  <=  0;
               conv_qin_00049_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00049_00000  <=  0;
               conv_qin_00049_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00049_00001  <=  0;
               conv_qin_00049_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00049_00002  <=  0;
               conv_qin_00049_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00049_00003  <=  0;
               conv_qin_00050_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00050_00000  <=  0;
               conv_qin_00050_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00050_00001  <=  0;
               conv_qin_00050_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00050_00002  <=  0;
               conv_qin_00050_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00050_00003  <=  0;
               conv_qin_00051_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00051_00000  <=  0;
               conv_qin_00051_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00051_00001  <=  0;
               conv_qin_00051_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00051_00002  <=  0;
               conv_qin_00051_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00051_00003  <=  0;
               conv_qin_00052_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00052_00000  <=  0;
               conv_qin_00052_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00052_00001  <=  0;
               conv_qin_00052_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00052_00002  <=  0;
               conv_qin_00052_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00052_00003  <=  0;
               conv_qin_00052_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00052_00004  <=  0;
               conv_qin_00053_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00053_00000  <=  0;
               conv_qin_00053_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00053_00001  <=  0;
               conv_qin_00053_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00053_00002  <=  0;
               conv_qin_00053_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00053_00003  <=  0;
               conv_qin_00053_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00053_00004  <=  0;
               conv_qin_00054_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00054_00000  <=  0;
               conv_qin_00054_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00054_00001  <=  0;
               conv_qin_00054_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00054_00002  <=  0;
               conv_qin_00054_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00054_00003  <=  0;
               conv_qin_00054_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00054_00004  <=  0;
               conv_qin_00055_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00055_00000  <=  0;
               conv_qin_00055_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00055_00001  <=  0;
               conv_qin_00055_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00055_00002  <=  0;
               conv_qin_00055_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00055_00003  <=  0;
               conv_qin_00055_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00055_00004  <=  0;
               conv_qin_00056_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00056_00000  <=  0;
               conv_qin_00056_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00056_00001  <=  0;
               conv_qin_00056_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00056_00002  <=  0;
               conv_qin_00056_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00056_00003  <=  0;
               conv_qin_00056_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00056_00004  <=  0;
               conv_qin_00057_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00057_00000  <=  0;
               conv_qin_00057_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00057_00001  <=  0;
               conv_qin_00057_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00057_00002  <=  0;
               conv_qin_00057_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00057_00003  <=  0;
               conv_qin_00057_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00057_00004  <=  0;
               conv_qin_00058_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00058_00000  <=  0;
               conv_qin_00058_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00058_00001  <=  0;
               conv_qin_00058_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00058_00002  <=  0;
               conv_qin_00058_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00058_00003  <=  0;
               conv_qin_00058_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00058_00004  <=  0;
               conv_qin_00059_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00059_00000  <=  0;
               conv_qin_00059_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00059_00001  <=  0;
               conv_qin_00059_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00059_00002  <=  0;
               conv_qin_00059_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00059_00003  <=  0;
               conv_qin_00059_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00059_00004  <=  0;
               conv_qin_00060_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00060_00000  <=  0;
               conv_qin_00060_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00060_00001  <=  0;
               conv_qin_00060_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00060_00002  <=  0;
               conv_qin_00060_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00060_00003  <=  0;
               conv_qin_00061_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00061_00000  <=  0;
               conv_qin_00061_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00061_00001  <=  0;
               conv_qin_00061_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00061_00002  <=  0;
               conv_qin_00061_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00061_00003  <=  0;
               conv_qin_00062_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00062_00000  <=  0;
               conv_qin_00062_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00062_00001  <=  0;
               conv_qin_00062_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00062_00002  <=  0;
               conv_qin_00062_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00062_00003  <=  0;
               conv_qin_00063_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00063_00000  <=  0;
               conv_qin_00063_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00063_00001  <=  0;
               conv_qin_00063_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00063_00002  <=  0;
               conv_qin_00063_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00063_00003  <=  0;
               conv_qin_00064_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00064_00000  <=  0;
               conv_qin_00064_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00064_00001  <=  0;
               conv_qin_00064_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00064_00002  <=  0;
               conv_qin_00064_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00064_00003  <=  0;
               conv_qin_00064_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00064_00004  <=  0;
               conv_qin_00065_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00065_00000  <=  0;
               conv_qin_00065_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00065_00001  <=  0;
               conv_qin_00065_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00065_00002  <=  0;
               conv_qin_00065_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00065_00003  <=  0;
               conv_qin_00065_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00065_00004  <=  0;
               conv_qin_00066_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00066_00000  <=  0;
               conv_qin_00066_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00066_00001  <=  0;
               conv_qin_00066_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00066_00002  <=  0;
               conv_qin_00066_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00066_00003  <=  0;
               conv_qin_00066_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00066_00004  <=  0;
               conv_qin_00067_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00067_00000  <=  0;
               conv_qin_00067_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00067_00001  <=  0;
               conv_qin_00067_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00067_00002  <=  0;
               conv_qin_00067_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00067_00003  <=  0;
               conv_qin_00067_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00067_00004  <=  0;
               conv_qin_00068_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00068_00000  <=  0;
               conv_qin_00068_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00068_00001  <=  0;
               conv_qin_00068_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00068_00002  <=  0;
               conv_qin_00068_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00068_00003  <=  0;
               conv_qin_00068_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00068_00004  <=  0;
               conv_qin_00069_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00069_00000  <=  0;
               conv_qin_00069_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00069_00001  <=  0;
               conv_qin_00069_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00069_00002  <=  0;
               conv_qin_00069_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00069_00003  <=  0;
               conv_qin_00069_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00069_00004  <=  0;
               conv_qin_00070_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00070_00000  <=  0;
               conv_qin_00070_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00070_00001  <=  0;
               conv_qin_00070_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00070_00002  <=  0;
               conv_qin_00070_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00070_00003  <=  0;
               conv_qin_00070_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00070_00004  <=  0;
               conv_qin_00071_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00071_00000  <=  0;
               conv_qin_00071_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00071_00001  <=  0;
               conv_qin_00071_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00071_00002  <=  0;
               conv_qin_00071_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00071_00003  <=  0;
               conv_qin_00071_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00071_00004  <=  0;
               conv_qin_00072_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00072_00000  <=  0;
               conv_qin_00072_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00072_00001  <=  0;
               conv_qin_00072_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00072_00002  <=  0;
               conv_qin_00072_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00072_00003  <=  0;
               conv_qin_00073_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00073_00000  <=  0;
               conv_qin_00073_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00073_00001  <=  0;
               conv_qin_00073_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00073_00002  <=  0;
               conv_qin_00073_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00073_00003  <=  0;
               conv_qin_00074_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00074_00000  <=  0;
               conv_qin_00074_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00074_00001  <=  0;
               conv_qin_00074_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00074_00002  <=  0;
               conv_qin_00074_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00074_00003  <=  0;
               conv_qin_00075_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00075_00000  <=  0;
               conv_qin_00075_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00075_00001  <=  0;
               conv_qin_00075_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00075_00002  <=  0;
               conv_qin_00075_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00075_00003  <=  0;
               conv_qin_00076_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00076_00000  <=  0;
               conv_qin_00076_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00076_00001  <=  0;
               conv_qin_00076_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00076_00002  <=  0;
               conv_qin_00076_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00076_00003  <=  0;
               conv_qin_00077_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00077_00000  <=  0;
               conv_qin_00077_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00077_00001  <=  0;
               conv_qin_00077_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00077_00002  <=  0;
               conv_qin_00077_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00077_00003  <=  0;
               conv_qin_00078_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00078_00000  <=  0;
               conv_qin_00078_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00078_00001  <=  0;
               conv_qin_00078_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00078_00002  <=  0;
               conv_qin_00078_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00078_00003  <=  0;
               conv_qin_00079_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00079_00000  <=  0;
               conv_qin_00079_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00079_00001  <=  0;
               conv_qin_00079_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00079_00002  <=  0;
               conv_qin_00079_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00079_00003  <=  0;
               conv_qin_00080_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00080_00000  <=  0;
               conv_qin_00080_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00080_00001  <=  0;
               conv_qin_00080_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00080_00002  <=  0;
               conv_qin_00080_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00080_00003  <=  0;
               conv_qin_00081_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00081_00000  <=  0;
               conv_qin_00081_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00081_00001  <=  0;
               conv_qin_00081_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00081_00002  <=  0;
               conv_qin_00081_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00081_00003  <=  0;
               conv_qin_00082_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00082_00000  <=  0;
               conv_qin_00082_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00082_00001  <=  0;
               conv_qin_00082_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00082_00002  <=  0;
               conv_qin_00082_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00082_00003  <=  0;
               conv_qin_00083_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00083_00000  <=  0;
               conv_qin_00083_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00083_00001  <=  0;
               conv_qin_00083_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00083_00002  <=  0;
               conv_qin_00083_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00083_00003  <=  0;
               conv_qin_00084_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00084_00000  <=  0;
               conv_qin_00084_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00084_00001  <=  0;
               conv_qin_00084_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00084_00002  <=  0;
               conv_qin_00084_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00084_00003  <=  0;
               conv_qin_00085_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00085_00000  <=  0;
               conv_qin_00085_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00085_00001  <=  0;
               conv_qin_00085_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00085_00002  <=  0;
               conv_qin_00085_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00085_00003  <=  0;
               conv_qin_00086_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00086_00000  <=  0;
               conv_qin_00086_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00086_00001  <=  0;
               conv_qin_00086_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00086_00002  <=  0;
               conv_qin_00086_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00086_00003  <=  0;
               conv_qin_00087_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00087_00000  <=  0;
               conv_qin_00087_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00087_00001  <=  0;
               conv_qin_00087_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00087_00002  <=  0;
               conv_qin_00087_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00087_00003  <=  0;
               conv_qin_00088_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00088_00000  <=  0;
               conv_qin_00088_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00088_00001  <=  0;
               conv_qin_00088_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00088_00002  <=  0;
               conv_qin_00089_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00089_00000  <=  0;
               conv_qin_00089_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00089_00001  <=  0;
               conv_qin_00089_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00089_00002  <=  0;
               conv_qin_00090_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00090_00000  <=  0;
               conv_qin_00090_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00090_00001  <=  0;
               conv_qin_00090_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00090_00002  <=  0;
               conv_qin_00091_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00091_00000  <=  0;
               conv_qin_00091_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00091_00001  <=  0;
               conv_qin_00091_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00091_00002  <=  0;
               conv_qin_00092_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00092_00000  <=  0;
               conv_qin_00092_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00092_00001  <=  0;
               conv_qin_00092_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00092_00002  <=  0;
               conv_qin_00092_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00092_00003  <=  0;
               conv_qin_00093_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00093_00000  <=  0;
               conv_qin_00093_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00093_00001  <=  0;
               conv_qin_00093_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00093_00002  <=  0;
               conv_qin_00093_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00093_00003  <=  0;
               conv_qin_00094_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00094_00000  <=  0;
               conv_qin_00094_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00094_00001  <=  0;
               conv_qin_00094_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00094_00002  <=  0;
               conv_qin_00094_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00094_00003  <=  0;
               conv_qin_00095_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00095_00000  <=  0;
               conv_qin_00095_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00095_00001  <=  0;
               conv_qin_00095_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00095_00002  <=  0;
               conv_qin_00095_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00095_00003  <=  0;
               conv_qin_00096_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00096_00000  <=  0;
               conv_qin_00096_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00096_00001  <=  0;
               conv_qin_00096_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00096_00002  <=  0;
               conv_qin_00096_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00096_00003  <=  0;
               conv_qin_00097_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00097_00000  <=  0;
               conv_qin_00097_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00097_00001  <=  0;
               conv_qin_00097_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00097_00002  <=  0;
               conv_qin_00097_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00097_00003  <=  0;
               conv_qin_00098_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00098_00000  <=  0;
               conv_qin_00098_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00098_00001  <=  0;
               conv_qin_00098_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00098_00002  <=  0;
               conv_qin_00098_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00098_00003  <=  0;
               conv_qin_00099_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00099_00000  <=  0;
               conv_qin_00099_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00099_00001  <=  0;
               conv_qin_00099_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00099_00002  <=  0;
               conv_qin_00099_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00099_00003  <=  0;
               conv_qin_00100_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00100_00000  <=  0;
               conv_qin_00100_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00100_00001  <=  0;
               conv_qin_00100_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00100_00002  <=  0;
               conv_qin_00101_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00101_00000  <=  0;
               conv_qin_00101_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00101_00001  <=  0;
               conv_qin_00101_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00101_00002  <=  0;
               conv_qin_00102_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00102_00000  <=  0;
               conv_qin_00102_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00102_00001  <=  0;
               conv_qin_00102_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00102_00002  <=  0;
               conv_qin_00103_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00103_00000  <=  0;
               conv_qin_00103_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00103_00001  <=  0;
               conv_qin_00103_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00103_00002  <=  0;
               conv_qin_00104_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00104_00000  <=  0;
               conv_qin_00104_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00104_00001  <=  0;
               conv_qin_00104_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00104_00002  <=  0;
               conv_qin_00104_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00104_00003  <=  0;
               conv_qin_00104_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00104_00004  <=  0;
               conv_qin_00105_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00105_00000  <=  0;
               conv_qin_00105_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00105_00001  <=  0;
               conv_qin_00105_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00105_00002  <=  0;
               conv_qin_00105_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00105_00003  <=  0;
               conv_qin_00105_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00105_00004  <=  0;
               conv_qin_00106_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00106_00000  <=  0;
               conv_qin_00106_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00106_00001  <=  0;
               conv_qin_00106_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00106_00002  <=  0;
               conv_qin_00106_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00106_00003  <=  0;
               conv_qin_00106_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00106_00004  <=  0;
               conv_qin_00107_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00107_00000  <=  0;
               conv_qin_00107_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00107_00001  <=  0;
               conv_qin_00107_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00107_00002  <=  0;
               conv_qin_00107_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00107_00003  <=  0;
               conv_qin_00107_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00107_00004  <=  0;
               conv_qin_00108_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00108_00000  <=  0;
               conv_qin_00108_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00108_00001  <=  0;
               conv_qin_00108_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00108_00002  <=  0;
               conv_qin_00109_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00109_00000  <=  0;
               conv_qin_00109_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00109_00001  <=  0;
               conv_qin_00109_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00109_00002  <=  0;
               conv_qin_00110_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00110_00000  <=  0;
               conv_qin_00110_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00110_00001  <=  0;
               conv_qin_00110_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00110_00002  <=  0;
               conv_qin_00111_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00111_00000  <=  0;
               conv_qin_00111_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00111_00001  <=  0;
               conv_qin_00111_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00111_00002  <=  0;
               conv_qin_00112_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00112_00000  <=  0;
               conv_qin_00112_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00112_00001  <=  0;
               conv_qin_00112_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00112_00002  <=  0;
               conv_qin_00112_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00112_00003  <=  0;
               conv_qin_00113_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00113_00000  <=  0;
               conv_qin_00113_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00113_00001  <=  0;
               conv_qin_00113_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00113_00002  <=  0;
               conv_qin_00113_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00113_00003  <=  0;
               conv_qin_00114_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00114_00000  <=  0;
               conv_qin_00114_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00114_00001  <=  0;
               conv_qin_00114_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00114_00002  <=  0;
               conv_qin_00114_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00114_00003  <=  0;
               conv_qin_00115_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00115_00000  <=  0;
               conv_qin_00115_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00115_00001  <=  0;
               conv_qin_00115_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00115_00002  <=  0;
               conv_qin_00115_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00115_00003  <=  0;
               conv_qin_00116_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00116_00000  <=  0;
               conv_qin_00116_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00116_00001  <=  0;
               conv_qin_00116_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00116_00002  <=  0;
               conv_qin_00117_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00117_00000  <=  0;
               conv_qin_00117_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00117_00001  <=  0;
               conv_qin_00117_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00117_00002  <=  0;
               conv_qin_00118_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00118_00000  <=  0;
               conv_qin_00118_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00118_00001  <=  0;
               conv_qin_00118_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00118_00002  <=  0;
               conv_qin_00119_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00119_00000  <=  0;
               conv_qin_00119_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00119_00001  <=  0;
               conv_qin_00119_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00119_00002  <=  0;
               conv_qin_00120_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00120_00000  <=  0;
               conv_qin_00120_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00120_00001  <=  0;
               conv_qin_00120_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00120_00002  <=  0;
               conv_qin_00120_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00120_00003  <=  0;
               conv_qin_00120_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00120_00004  <=  0;
               conv_qin_00121_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00121_00000  <=  0;
               conv_qin_00121_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00121_00001  <=  0;
               conv_qin_00121_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00121_00002  <=  0;
               conv_qin_00121_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00121_00003  <=  0;
               conv_qin_00121_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00121_00004  <=  0;
               conv_qin_00122_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00122_00000  <=  0;
               conv_qin_00122_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00122_00001  <=  0;
               conv_qin_00122_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00122_00002  <=  0;
               conv_qin_00122_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00122_00003  <=  0;
               conv_qin_00122_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00122_00004  <=  0;
               conv_qin_00123_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00123_00000  <=  0;
               conv_qin_00123_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00123_00001  <=  0;
               conv_qin_00123_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00123_00002  <=  0;
               conv_qin_00123_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00123_00003  <=  0;
               conv_qin_00123_00004  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00123_00004  <=  0;
               conv_qin_00124_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00124_00000  <=  0;
               conv_qin_00124_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00124_00001  <=  0;
               conv_qin_00124_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00124_00002  <=  0;
               conv_qin_00125_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00125_00000  <=  0;
               conv_qin_00125_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00125_00001  <=  0;
               conv_qin_00125_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00125_00002  <=  0;
               conv_qin_00126_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00126_00000  <=  0;
               conv_qin_00126_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00126_00001  <=  0;
               conv_qin_00126_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00126_00002  <=  0;
               conv_qin_00127_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00127_00000  <=  0;
               conv_qin_00127_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00127_00001  <=  0;
               conv_qin_00127_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00127_00002  <=  0;
               conv_qin_00128_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00128_00000  <=  0;
               conv_qin_00128_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00128_00001  <=  0;
               conv_qin_00128_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00128_00002  <=  0;
               conv_qin_00128_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00128_00003  <=  0;
               conv_qin_00129_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00129_00000  <=  0;
               conv_qin_00129_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00129_00001  <=  0;
               conv_qin_00129_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00129_00002  <=  0;
               conv_qin_00129_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00129_00003  <=  0;
               conv_qin_00130_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00130_00000  <=  0;
               conv_qin_00130_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00130_00001  <=  0;
               conv_qin_00130_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00130_00002  <=  0;
               conv_qin_00130_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00130_00003  <=  0;
               conv_qin_00131_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00131_00000  <=  0;
               conv_qin_00131_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00131_00001  <=  0;
               conv_qin_00131_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00131_00002  <=  0;
               conv_qin_00131_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00131_00003  <=  0;
               conv_qin_00132_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00132_00000  <=  0;
               conv_qin_00132_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00132_00001  <=  0;
               conv_qin_00132_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00132_00002  <=  0;
               conv_qin_00132_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00132_00003  <=  0;
               conv_qin_00133_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00133_00000  <=  0;
               conv_qin_00133_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00133_00001  <=  0;
               conv_qin_00133_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00133_00002  <=  0;
               conv_qin_00133_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00133_00003  <=  0;
               conv_qin_00134_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00134_00000  <=  0;
               conv_qin_00134_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00134_00001  <=  0;
               conv_qin_00134_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00134_00002  <=  0;
               conv_qin_00134_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00134_00003  <=  0;
               conv_qin_00135_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00135_00000  <=  0;
               conv_qin_00135_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00135_00001  <=  0;
               conv_qin_00135_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00135_00002  <=  0;
               conv_qin_00135_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00135_00003  <=  0;
               conv_qin_00136_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00136_00000  <=  0;
               conv_qin_00136_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00136_00001  <=  0;
               conv_qin_00136_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00136_00002  <=  0;
               conv_qin_00136_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00136_00003  <=  0;
               conv_qin_00137_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00137_00000  <=  0;
               conv_qin_00137_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00137_00001  <=  0;
               conv_qin_00137_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00137_00002  <=  0;
               conv_qin_00137_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00137_00003  <=  0;
               conv_qin_00138_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00138_00000  <=  0;
               conv_qin_00138_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00138_00001  <=  0;
               conv_qin_00138_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00138_00002  <=  0;
               conv_qin_00138_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00138_00003  <=  0;
               conv_qin_00139_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00139_00000  <=  0;
               conv_qin_00139_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00139_00001  <=  0;
               conv_qin_00139_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00139_00002  <=  0;
               conv_qin_00139_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00139_00003  <=  0;
               conv_qin_00140_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00140_00000  <=  0;
               conv_qin_00140_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00140_00001  <=  0;
               conv_qin_00140_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00140_00002  <=  0;
               conv_qin_00140_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00140_00003  <=  0;
               conv_qin_00141_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00141_00000  <=  0;
               conv_qin_00141_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00141_00001  <=  0;
               conv_qin_00141_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00141_00002  <=  0;
               conv_qin_00141_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00141_00003  <=  0;
               conv_qin_00142_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00142_00000  <=  0;
               conv_qin_00142_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00142_00001  <=  0;
               conv_qin_00142_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00142_00002  <=  0;
               conv_qin_00142_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00142_00003  <=  0;
               conv_qin_00143_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00143_00000  <=  0;
               conv_qin_00143_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00143_00001  <=  0;
               conv_qin_00143_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00143_00002  <=  0;
               conv_qin_00143_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00143_00003  <=  0;
               conv_qin_00144_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00144_00000  <=  0;
               conv_qin_00144_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00144_00001  <=  0;
               conv_qin_00144_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00144_00002  <=  0;
               conv_qin_00144_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00144_00003  <=  0;
               conv_qin_00145_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00145_00000  <=  0;
               conv_qin_00145_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00145_00001  <=  0;
               conv_qin_00145_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00145_00002  <=  0;
               conv_qin_00145_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00145_00003  <=  0;
               conv_qin_00146_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00146_00000  <=  0;
               conv_qin_00146_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00146_00001  <=  0;
               conv_qin_00146_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00146_00002  <=  0;
               conv_qin_00146_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00146_00003  <=  0;
               conv_qin_00147_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00147_00000  <=  0;
               conv_qin_00147_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00147_00001  <=  0;
               conv_qin_00147_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00147_00002  <=  0;
               conv_qin_00147_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00147_00003  <=  0;
               conv_qin_00148_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00148_00000  <=  0;
               conv_qin_00148_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00148_00001  <=  0;
               conv_qin_00148_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00148_00002  <=  0;
               conv_qin_00149_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00149_00000  <=  0;
               conv_qin_00149_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00149_00001  <=  0;
               conv_qin_00149_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00149_00002  <=  0;
               conv_qin_00150_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00150_00000  <=  0;
               conv_qin_00150_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00150_00001  <=  0;
               conv_qin_00150_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00150_00002  <=  0;
               conv_qin_00151_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00151_00000  <=  0;
               conv_qin_00151_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00151_00001  <=  0;
               conv_qin_00151_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00151_00002  <=  0;
               conv_qin_00152_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00152_00000  <=  0;
               conv_qin_00152_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00152_00001  <=  0;
               conv_qin_00152_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00152_00002  <=  0;
               conv_qin_00152_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00152_00003  <=  0;
               conv_qin_00153_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00153_00000  <=  0;
               conv_qin_00153_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00153_00001  <=  0;
               conv_qin_00153_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00153_00002  <=  0;
               conv_qin_00153_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00153_00003  <=  0;
               conv_qin_00154_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00154_00000  <=  0;
               conv_qin_00154_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00154_00001  <=  0;
               conv_qin_00154_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00154_00002  <=  0;
               conv_qin_00154_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00154_00003  <=  0;
               conv_qin_00155_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00155_00000  <=  0;
               conv_qin_00155_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00155_00001  <=  0;
               conv_qin_00155_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00155_00002  <=  0;
               conv_qin_00155_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00155_00003  <=  0;
               conv_qin_00156_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00156_00000  <=  0;
               conv_qin_00156_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00156_00001  <=  0;
               conv_qin_00156_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00156_00002  <=  0;
               conv_qin_00156_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00156_00003  <=  0;
               conv_qin_00157_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00157_00000  <=  0;
               conv_qin_00157_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00157_00001  <=  0;
               conv_qin_00157_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00157_00002  <=  0;
               conv_qin_00157_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00157_00003  <=  0;
               conv_qin_00158_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00158_00000  <=  0;
               conv_qin_00158_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00158_00001  <=  0;
               conv_qin_00158_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00158_00002  <=  0;
               conv_qin_00158_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00158_00003  <=  0;
               conv_qin_00159_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00159_00000  <=  0;
               conv_qin_00159_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00159_00001  <=  0;
               conv_qin_00159_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00159_00002  <=  0;
               conv_qin_00159_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00159_00003  <=  0;
               conv_qin_00160_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00160_00000  <=  0;
               conv_qin_00160_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00160_00001  <=  0;
               conv_qin_00160_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00160_00002  <=  0;
               conv_qin_00160_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00160_00003  <=  0;
               conv_qin_00161_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00161_00000  <=  0;
               conv_qin_00161_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00161_00001  <=  0;
               conv_qin_00161_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00161_00002  <=  0;
               conv_qin_00161_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00161_00003  <=  0;
               conv_qin_00162_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00162_00000  <=  0;
               conv_qin_00162_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00162_00001  <=  0;
               conv_qin_00162_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00162_00002  <=  0;
               conv_qin_00162_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00162_00003  <=  0;
               conv_qin_00163_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00163_00000  <=  0;
               conv_qin_00163_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00163_00001  <=  0;
               conv_qin_00163_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00163_00002  <=  0;
               conv_qin_00163_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00163_00003  <=  0;
               conv_qin_00164_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00164_00000  <=  0;
               conv_qin_00164_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00164_00001  <=  0;
               conv_qin_00164_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00164_00002  <=  0;
               conv_qin_00164_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00164_00003  <=  0;
               conv_qin_00165_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00165_00000  <=  0;
               conv_qin_00165_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00165_00001  <=  0;
               conv_qin_00165_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00165_00002  <=  0;
               conv_qin_00165_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00165_00003  <=  0;
               conv_qin_00166_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00166_00000  <=  0;
               conv_qin_00166_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00166_00001  <=  0;
               conv_qin_00166_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00166_00002  <=  0;
               conv_qin_00166_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00166_00003  <=  0;
               conv_qin_00167_00000  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00167_00000  <=  0;
               conv_qin_00167_00001  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00167_00001  <=  0;
               conv_qin_00167_00002  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00167_00002  <=  0;
               conv_qin_00167_00003  <= {(MAX_SUM_WDTH_L){1'b0}};
               sign_qin_00167_00003  <=  0;
       end else begin
            // Id66554a95b5375bec1ec7c8e6bbfea7d and tout should come Ied2b5c0139cec8ad2873829dc1117d50 same clock
             if (start_d5) begin
                if (sgnprod_00000 == conv_Sgntin_row_00000_00000 ) begin
                    conv_qin_00000_00000  <= tout_00000_00000;
                    sign_qin_00000_00000  <=  0;
                end else begin
                    conv_qin_00000_00000  <=  ~tout_00000_00000 + 1;
                    sign_qin_00000_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00000 == conv_Sgntin_row_00000_00001 ) begin
                    conv_qin_00000_00001  <= tout_00000_00001;
                    sign_qin_00000_00001  <=  0;
                end else begin
                    conv_qin_00000_00001  <=  ~tout_00000_00001 + 1;
                    sign_qin_00000_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00000 == conv_Sgntin_row_00000_00002 ) begin
                    conv_qin_00000_00002  <= tout_00000_00002;
                    sign_qin_00000_00002  <=  0;
                end else begin
                    conv_qin_00000_00002  <=  ~tout_00000_00002 + 1;
                    sign_qin_00000_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00000 == conv_Sgntin_row_00000_00003 ) begin
                    conv_qin_00000_00003  <= tout_00000_00003;
                    sign_qin_00000_00003  <=  0;
                end else begin
                    conv_qin_00000_00003  <=  ~tout_00000_00003 + 1;
                    sign_qin_00000_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00000 == conv_Sgntin_row_00000_00004 ) begin
                    conv_qin_00000_00004  <= tout_00000_00004;
                    sign_qin_00000_00004  <=  0;
                end else begin
                    conv_qin_00000_00004  <=  ~tout_00000_00004 + 1;
                    sign_qin_00000_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00000 == conv_Sgntin_row_00000_00005 ) begin
                    conv_qin_00000_00005  <= tout_00000_00005;
                    sign_qin_00000_00005  <=  0;
                end else begin
                    conv_qin_00000_00005  <=  ~tout_00000_00005 + 1;
                    sign_qin_00000_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00000 == conv_Sgntin_row_00000_00006 ) begin
                    conv_qin_00000_00006  <= tout_00000_00006;
                    sign_qin_00000_00006  <=  0;
                end else begin
                    conv_qin_00000_00006  <=  ~tout_00000_00006 + 1;
                    sign_qin_00000_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00000 == conv_Sgntin_row_00000_00007 ) begin
                    conv_qin_00000_00007  <= tout_00000_00007;
                    sign_qin_00000_00007  <=  0;
                end else begin
                    conv_qin_00000_00007  <=  ~tout_00000_00007 + 1;
                    sign_qin_00000_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00001 == conv_Sgntin_row_00001_00000 ) begin
                    conv_qin_00001_00000  <= tout_00001_00000;
                    sign_qin_00001_00000  <=  0;
                end else begin
                    conv_qin_00001_00000  <=  ~tout_00001_00000 + 1;
                    sign_qin_00001_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00001 == conv_Sgntin_row_00001_00001 ) begin
                    conv_qin_00001_00001  <= tout_00001_00001;
                    sign_qin_00001_00001  <=  0;
                end else begin
                    conv_qin_00001_00001  <=  ~tout_00001_00001 + 1;
                    sign_qin_00001_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00001 == conv_Sgntin_row_00001_00002 ) begin
                    conv_qin_00001_00002  <= tout_00001_00002;
                    sign_qin_00001_00002  <=  0;
                end else begin
                    conv_qin_00001_00002  <=  ~tout_00001_00002 + 1;
                    sign_qin_00001_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00001 == conv_Sgntin_row_00001_00003 ) begin
                    conv_qin_00001_00003  <= tout_00001_00003;
                    sign_qin_00001_00003  <=  0;
                end else begin
                    conv_qin_00001_00003  <=  ~tout_00001_00003 + 1;
                    sign_qin_00001_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00001 == conv_Sgntin_row_00001_00004 ) begin
                    conv_qin_00001_00004  <= tout_00001_00004;
                    sign_qin_00001_00004  <=  0;
                end else begin
                    conv_qin_00001_00004  <=  ~tout_00001_00004 + 1;
                    sign_qin_00001_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00001 == conv_Sgntin_row_00001_00005 ) begin
                    conv_qin_00001_00005  <= tout_00001_00005;
                    sign_qin_00001_00005  <=  0;
                end else begin
                    conv_qin_00001_00005  <=  ~tout_00001_00005 + 1;
                    sign_qin_00001_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00001 == conv_Sgntin_row_00001_00006 ) begin
                    conv_qin_00001_00006  <= tout_00001_00006;
                    sign_qin_00001_00006  <=  0;
                end else begin
                    conv_qin_00001_00006  <=  ~tout_00001_00006 + 1;
                    sign_qin_00001_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00001 == conv_Sgntin_row_00001_00007 ) begin
                    conv_qin_00001_00007  <= tout_00001_00007;
                    sign_qin_00001_00007  <=  0;
                end else begin
                    conv_qin_00001_00007  <=  ~tout_00001_00007 + 1;
                    sign_qin_00001_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00002 == conv_Sgntin_row_00002_00000 ) begin
                    conv_qin_00002_00000  <= tout_00002_00000;
                    sign_qin_00002_00000  <=  0;
                end else begin
                    conv_qin_00002_00000  <=  ~tout_00002_00000 + 1;
                    sign_qin_00002_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00002 == conv_Sgntin_row_00002_00001 ) begin
                    conv_qin_00002_00001  <= tout_00002_00001;
                    sign_qin_00002_00001  <=  0;
                end else begin
                    conv_qin_00002_00001  <=  ~tout_00002_00001 + 1;
                    sign_qin_00002_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00002 == conv_Sgntin_row_00002_00002 ) begin
                    conv_qin_00002_00002  <= tout_00002_00002;
                    sign_qin_00002_00002  <=  0;
                end else begin
                    conv_qin_00002_00002  <=  ~tout_00002_00002 + 1;
                    sign_qin_00002_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00002 == conv_Sgntin_row_00002_00003 ) begin
                    conv_qin_00002_00003  <= tout_00002_00003;
                    sign_qin_00002_00003  <=  0;
                end else begin
                    conv_qin_00002_00003  <=  ~tout_00002_00003 + 1;
                    sign_qin_00002_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00002 == conv_Sgntin_row_00002_00004 ) begin
                    conv_qin_00002_00004  <= tout_00002_00004;
                    sign_qin_00002_00004  <=  0;
                end else begin
                    conv_qin_00002_00004  <=  ~tout_00002_00004 + 1;
                    sign_qin_00002_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00002 == conv_Sgntin_row_00002_00005 ) begin
                    conv_qin_00002_00005  <= tout_00002_00005;
                    sign_qin_00002_00005  <=  0;
                end else begin
                    conv_qin_00002_00005  <=  ~tout_00002_00005 + 1;
                    sign_qin_00002_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00002 == conv_Sgntin_row_00002_00006 ) begin
                    conv_qin_00002_00006  <= tout_00002_00006;
                    sign_qin_00002_00006  <=  0;
                end else begin
                    conv_qin_00002_00006  <=  ~tout_00002_00006 + 1;
                    sign_qin_00002_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00002 == conv_Sgntin_row_00002_00007 ) begin
                    conv_qin_00002_00007  <= tout_00002_00007;
                    sign_qin_00002_00007  <=  0;
                end else begin
                    conv_qin_00002_00007  <=  ~tout_00002_00007 + 1;
                    sign_qin_00002_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00003 == conv_Sgntin_row_00003_00000 ) begin
                    conv_qin_00003_00000  <= tout_00003_00000;
                    sign_qin_00003_00000  <=  0;
                end else begin
                    conv_qin_00003_00000  <=  ~tout_00003_00000 + 1;
                    sign_qin_00003_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00003 == conv_Sgntin_row_00003_00001 ) begin
                    conv_qin_00003_00001  <= tout_00003_00001;
                    sign_qin_00003_00001  <=  0;
                end else begin
                    conv_qin_00003_00001  <=  ~tout_00003_00001 + 1;
                    sign_qin_00003_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00003 == conv_Sgntin_row_00003_00002 ) begin
                    conv_qin_00003_00002  <= tout_00003_00002;
                    sign_qin_00003_00002  <=  0;
                end else begin
                    conv_qin_00003_00002  <=  ~tout_00003_00002 + 1;
                    sign_qin_00003_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00003 == conv_Sgntin_row_00003_00003 ) begin
                    conv_qin_00003_00003  <= tout_00003_00003;
                    sign_qin_00003_00003  <=  0;
                end else begin
                    conv_qin_00003_00003  <=  ~tout_00003_00003 + 1;
                    sign_qin_00003_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00003 == conv_Sgntin_row_00003_00004 ) begin
                    conv_qin_00003_00004  <= tout_00003_00004;
                    sign_qin_00003_00004  <=  0;
                end else begin
                    conv_qin_00003_00004  <=  ~tout_00003_00004 + 1;
                    sign_qin_00003_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00003 == conv_Sgntin_row_00003_00005 ) begin
                    conv_qin_00003_00005  <= tout_00003_00005;
                    sign_qin_00003_00005  <=  0;
                end else begin
                    conv_qin_00003_00005  <=  ~tout_00003_00005 + 1;
                    sign_qin_00003_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00003 == conv_Sgntin_row_00003_00006 ) begin
                    conv_qin_00003_00006  <= tout_00003_00006;
                    sign_qin_00003_00006  <=  0;
                end else begin
                    conv_qin_00003_00006  <=  ~tout_00003_00006 + 1;
                    sign_qin_00003_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00003 == conv_Sgntin_row_00003_00007 ) begin
                    conv_qin_00003_00007  <= tout_00003_00007;
                    sign_qin_00003_00007  <=  0;
                end else begin
                    conv_qin_00003_00007  <=  ~tout_00003_00007 + 1;
                    sign_qin_00003_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00004 == conv_Sgntin_row_00004_00000 ) begin
                    conv_qin_00004_00000  <= tout_00004_00000;
                    sign_qin_00004_00000  <=  0;
                end else begin
                    conv_qin_00004_00000  <=  ~tout_00004_00000 + 1;
                    sign_qin_00004_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00004 == conv_Sgntin_row_00004_00001 ) begin
                    conv_qin_00004_00001  <= tout_00004_00001;
                    sign_qin_00004_00001  <=  0;
                end else begin
                    conv_qin_00004_00001  <=  ~tout_00004_00001 + 1;
                    sign_qin_00004_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00004 == conv_Sgntin_row_00004_00002 ) begin
                    conv_qin_00004_00002  <= tout_00004_00002;
                    sign_qin_00004_00002  <=  0;
                end else begin
                    conv_qin_00004_00002  <=  ~tout_00004_00002 + 1;
                    sign_qin_00004_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00004 == conv_Sgntin_row_00004_00003 ) begin
                    conv_qin_00004_00003  <= tout_00004_00003;
                    sign_qin_00004_00003  <=  0;
                end else begin
                    conv_qin_00004_00003  <=  ~tout_00004_00003 + 1;
                    sign_qin_00004_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00004 == conv_Sgntin_row_00004_00004 ) begin
                    conv_qin_00004_00004  <= tout_00004_00004;
                    sign_qin_00004_00004  <=  0;
                end else begin
                    conv_qin_00004_00004  <=  ~tout_00004_00004 + 1;
                    sign_qin_00004_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00004 == conv_Sgntin_row_00004_00005 ) begin
                    conv_qin_00004_00005  <= tout_00004_00005;
                    sign_qin_00004_00005  <=  0;
                end else begin
                    conv_qin_00004_00005  <=  ~tout_00004_00005 + 1;
                    sign_qin_00004_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00004 == conv_Sgntin_row_00004_00006 ) begin
                    conv_qin_00004_00006  <= tout_00004_00006;
                    sign_qin_00004_00006  <=  0;
                end else begin
                    conv_qin_00004_00006  <=  ~tout_00004_00006 + 1;
                    sign_qin_00004_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00004 == conv_Sgntin_row_00004_00007 ) begin
                    conv_qin_00004_00007  <= tout_00004_00007;
                    sign_qin_00004_00007  <=  0;
                end else begin
                    conv_qin_00004_00007  <=  ~tout_00004_00007 + 1;
                    sign_qin_00004_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00004 == conv_Sgntin_row_00004_00008 ) begin
                    conv_qin_00004_00008  <= tout_00004_00008;
                    sign_qin_00004_00008  <=  0;
                end else begin
                    conv_qin_00004_00008  <=  ~tout_00004_00008 + 1;
                    sign_qin_00004_00008  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00004 == conv_Sgntin_row_00004_00009 ) begin
                    conv_qin_00004_00009  <= tout_00004_00009;
                    sign_qin_00004_00009  <=  0;
                end else begin
                    conv_qin_00004_00009  <=  ~tout_00004_00009 + 1;
                    sign_qin_00004_00009  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00005 == conv_Sgntin_row_00005_00000 ) begin
                    conv_qin_00005_00000  <= tout_00005_00000;
                    sign_qin_00005_00000  <=  0;
                end else begin
                    conv_qin_00005_00000  <=  ~tout_00005_00000 + 1;
                    sign_qin_00005_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00005 == conv_Sgntin_row_00005_00001 ) begin
                    conv_qin_00005_00001  <= tout_00005_00001;
                    sign_qin_00005_00001  <=  0;
                end else begin
                    conv_qin_00005_00001  <=  ~tout_00005_00001 + 1;
                    sign_qin_00005_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00005 == conv_Sgntin_row_00005_00002 ) begin
                    conv_qin_00005_00002  <= tout_00005_00002;
                    sign_qin_00005_00002  <=  0;
                end else begin
                    conv_qin_00005_00002  <=  ~tout_00005_00002 + 1;
                    sign_qin_00005_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00005 == conv_Sgntin_row_00005_00003 ) begin
                    conv_qin_00005_00003  <= tout_00005_00003;
                    sign_qin_00005_00003  <=  0;
                end else begin
                    conv_qin_00005_00003  <=  ~tout_00005_00003 + 1;
                    sign_qin_00005_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00005 == conv_Sgntin_row_00005_00004 ) begin
                    conv_qin_00005_00004  <= tout_00005_00004;
                    sign_qin_00005_00004  <=  0;
                end else begin
                    conv_qin_00005_00004  <=  ~tout_00005_00004 + 1;
                    sign_qin_00005_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00005 == conv_Sgntin_row_00005_00005 ) begin
                    conv_qin_00005_00005  <= tout_00005_00005;
                    sign_qin_00005_00005  <=  0;
                end else begin
                    conv_qin_00005_00005  <=  ~tout_00005_00005 + 1;
                    sign_qin_00005_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00005 == conv_Sgntin_row_00005_00006 ) begin
                    conv_qin_00005_00006  <= tout_00005_00006;
                    sign_qin_00005_00006  <=  0;
                end else begin
                    conv_qin_00005_00006  <=  ~tout_00005_00006 + 1;
                    sign_qin_00005_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00005 == conv_Sgntin_row_00005_00007 ) begin
                    conv_qin_00005_00007  <= tout_00005_00007;
                    sign_qin_00005_00007  <=  0;
                end else begin
                    conv_qin_00005_00007  <=  ~tout_00005_00007 + 1;
                    sign_qin_00005_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00005 == conv_Sgntin_row_00005_00008 ) begin
                    conv_qin_00005_00008  <= tout_00005_00008;
                    sign_qin_00005_00008  <=  0;
                end else begin
                    conv_qin_00005_00008  <=  ~tout_00005_00008 + 1;
                    sign_qin_00005_00008  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00005 == conv_Sgntin_row_00005_00009 ) begin
                    conv_qin_00005_00009  <= tout_00005_00009;
                    sign_qin_00005_00009  <=  0;
                end else begin
                    conv_qin_00005_00009  <=  ~tout_00005_00009 + 1;
                    sign_qin_00005_00009  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00006 == conv_Sgntin_row_00006_00000 ) begin
                    conv_qin_00006_00000  <= tout_00006_00000;
                    sign_qin_00006_00000  <=  0;
                end else begin
                    conv_qin_00006_00000  <=  ~tout_00006_00000 + 1;
                    sign_qin_00006_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00006 == conv_Sgntin_row_00006_00001 ) begin
                    conv_qin_00006_00001  <= tout_00006_00001;
                    sign_qin_00006_00001  <=  0;
                end else begin
                    conv_qin_00006_00001  <=  ~tout_00006_00001 + 1;
                    sign_qin_00006_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00006 == conv_Sgntin_row_00006_00002 ) begin
                    conv_qin_00006_00002  <= tout_00006_00002;
                    sign_qin_00006_00002  <=  0;
                end else begin
                    conv_qin_00006_00002  <=  ~tout_00006_00002 + 1;
                    sign_qin_00006_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00006 == conv_Sgntin_row_00006_00003 ) begin
                    conv_qin_00006_00003  <= tout_00006_00003;
                    sign_qin_00006_00003  <=  0;
                end else begin
                    conv_qin_00006_00003  <=  ~tout_00006_00003 + 1;
                    sign_qin_00006_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00006 == conv_Sgntin_row_00006_00004 ) begin
                    conv_qin_00006_00004  <= tout_00006_00004;
                    sign_qin_00006_00004  <=  0;
                end else begin
                    conv_qin_00006_00004  <=  ~tout_00006_00004 + 1;
                    sign_qin_00006_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00006 == conv_Sgntin_row_00006_00005 ) begin
                    conv_qin_00006_00005  <= tout_00006_00005;
                    sign_qin_00006_00005  <=  0;
                end else begin
                    conv_qin_00006_00005  <=  ~tout_00006_00005 + 1;
                    sign_qin_00006_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00006 == conv_Sgntin_row_00006_00006 ) begin
                    conv_qin_00006_00006  <= tout_00006_00006;
                    sign_qin_00006_00006  <=  0;
                end else begin
                    conv_qin_00006_00006  <=  ~tout_00006_00006 + 1;
                    sign_qin_00006_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00006 == conv_Sgntin_row_00006_00007 ) begin
                    conv_qin_00006_00007  <= tout_00006_00007;
                    sign_qin_00006_00007  <=  0;
                end else begin
                    conv_qin_00006_00007  <=  ~tout_00006_00007 + 1;
                    sign_qin_00006_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00006 == conv_Sgntin_row_00006_00008 ) begin
                    conv_qin_00006_00008  <= tout_00006_00008;
                    sign_qin_00006_00008  <=  0;
                end else begin
                    conv_qin_00006_00008  <=  ~tout_00006_00008 + 1;
                    sign_qin_00006_00008  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00006 == conv_Sgntin_row_00006_00009 ) begin
                    conv_qin_00006_00009  <= tout_00006_00009;
                    sign_qin_00006_00009  <=  0;
                end else begin
                    conv_qin_00006_00009  <=  ~tout_00006_00009 + 1;
                    sign_qin_00006_00009  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00007 == conv_Sgntin_row_00007_00000 ) begin
                    conv_qin_00007_00000  <= tout_00007_00000;
                    sign_qin_00007_00000  <=  0;
                end else begin
                    conv_qin_00007_00000  <=  ~tout_00007_00000 + 1;
                    sign_qin_00007_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00007 == conv_Sgntin_row_00007_00001 ) begin
                    conv_qin_00007_00001  <= tout_00007_00001;
                    sign_qin_00007_00001  <=  0;
                end else begin
                    conv_qin_00007_00001  <=  ~tout_00007_00001 + 1;
                    sign_qin_00007_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00007 == conv_Sgntin_row_00007_00002 ) begin
                    conv_qin_00007_00002  <= tout_00007_00002;
                    sign_qin_00007_00002  <=  0;
                end else begin
                    conv_qin_00007_00002  <=  ~tout_00007_00002 + 1;
                    sign_qin_00007_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00007 == conv_Sgntin_row_00007_00003 ) begin
                    conv_qin_00007_00003  <= tout_00007_00003;
                    sign_qin_00007_00003  <=  0;
                end else begin
                    conv_qin_00007_00003  <=  ~tout_00007_00003 + 1;
                    sign_qin_00007_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00007 == conv_Sgntin_row_00007_00004 ) begin
                    conv_qin_00007_00004  <= tout_00007_00004;
                    sign_qin_00007_00004  <=  0;
                end else begin
                    conv_qin_00007_00004  <=  ~tout_00007_00004 + 1;
                    sign_qin_00007_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00007 == conv_Sgntin_row_00007_00005 ) begin
                    conv_qin_00007_00005  <= tout_00007_00005;
                    sign_qin_00007_00005  <=  0;
                end else begin
                    conv_qin_00007_00005  <=  ~tout_00007_00005 + 1;
                    sign_qin_00007_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00007 == conv_Sgntin_row_00007_00006 ) begin
                    conv_qin_00007_00006  <= tout_00007_00006;
                    sign_qin_00007_00006  <=  0;
                end else begin
                    conv_qin_00007_00006  <=  ~tout_00007_00006 + 1;
                    sign_qin_00007_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00007 == conv_Sgntin_row_00007_00007 ) begin
                    conv_qin_00007_00007  <= tout_00007_00007;
                    sign_qin_00007_00007  <=  0;
                end else begin
                    conv_qin_00007_00007  <=  ~tout_00007_00007 + 1;
                    sign_qin_00007_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00007 == conv_Sgntin_row_00007_00008 ) begin
                    conv_qin_00007_00008  <= tout_00007_00008;
                    sign_qin_00007_00008  <=  0;
                end else begin
                    conv_qin_00007_00008  <=  ~tout_00007_00008 + 1;
                    sign_qin_00007_00008  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00007 == conv_Sgntin_row_00007_00009 ) begin
                    conv_qin_00007_00009  <= tout_00007_00009;
                    sign_qin_00007_00009  <=  0;
                end else begin
                    conv_qin_00007_00009  <=  ~tout_00007_00009 + 1;
                    sign_qin_00007_00009  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00008 == conv_Sgntin_row_00008_00000 ) begin
                    conv_qin_00008_00000  <= tout_00008_00000;
                    sign_qin_00008_00000  <=  0;
                end else begin
                    conv_qin_00008_00000  <=  ~tout_00008_00000 + 1;
                    sign_qin_00008_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00008 == conv_Sgntin_row_00008_00001 ) begin
                    conv_qin_00008_00001  <= tout_00008_00001;
                    sign_qin_00008_00001  <=  0;
                end else begin
                    conv_qin_00008_00001  <=  ~tout_00008_00001 + 1;
                    sign_qin_00008_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00008 == conv_Sgntin_row_00008_00002 ) begin
                    conv_qin_00008_00002  <= tout_00008_00002;
                    sign_qin_00008_00002  <=  0;
                end else begin
                    conv_qin_00008_00002  <=  ~tout_00008_00002 + 1;
                    sign_qin_00008_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00008 == conv_Sgntin_row_00008_00003 ) begin
                    conv_qin_00008_00003  <= tout_00008_00003;
                    sign_qin_00008_00003  <=  0;
                end else begin
                    conv_qin_00008_00003  <=  ~tout_00008_00003 + 1;
                    sign_qin_00008_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00008 == conv_Sgntin_row_00008_00004 ) begin
                    conv_qin_00008_00004  <= tout_00008_00004;
                    sign_qin_00008_00004  <=  0;
                end else begin
                    conv_qin_00008_00004  <=  ~tout_00008_00004 + 1;
                    sign_qin_00008_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00008 == conv_Sgntin_row_00008_00005 ) begin
                    conv_qin_00008_00005  <= tout_00008_00005;
                    sign_qin_00008_00005  <=  0;
                end else begin
                    conv_qin_00008_00005  <=  ~tout_00008_00005 + 1;
                    sign_qin_00008_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00008 == conv_Sgntin_row_00008_00006 ) begin
                    conv_qin_00008_00006  <= tout_00008_00006;
                    sign_qin_00008_00006  <=  0;
                end else begin
                    conv_qin_00008_00006  <=  ~tout_00008_00006 + 1;
                    sign_qin_00008_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00008 == conv_Sgntin_row_00008_00007 ) begin
                    conv_qin_00008_00007  <= tout_00008_00007;
                    sign_qin_00008_00007  <=  0;
                end else begin
                    conv_qin_00008_00007  <=  ~tout_00008_00007 + 1;
                    sign_qin_00008_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00009 == conv_Sgntin_row_00009_00000 ) begin
                    conv_qin_00009_00000  <= tout_00009_00000;
                    sign_qin_00009_00000  <=  0;
                end else begin
                    conv_qin_00009_00000  <=  ~tout_00009_00000 + 1;
                    sign_qin_00009_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00009 == conv_Sgntin_row_00009_00001 ) begin
                    conv_qin_00009_00001  <= tout_00009_00001;
                    sign_qin_00009_00001  <=  0;
                end else begin
                    conv_qin_00009_00001  <=  ~tout_00009_00001 + 1;
                    sign_qin_00009_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00009 == conv_Sgntin_row_00009_00002 ) begin
                    conv_qin_00009_00002  <= tout_00009_00002;
                    sign_qin_00009_00002  <=  0;
                end else begin
                    conv_qin_00009_00002  <=  ~tout_00009_00002 + 1;
                    sign_qin_00009_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00009 == conv_Sgntin_row_00009_00003 ) begin
                    conv_qin_00009_00003  <= tout_00009_00003;
                    sign_qin_00009_00003  <=  0;
                end else begin
                    conv_qin_00009_00003  <=  ~tout_00009_00003 + 1;
                    sign_qin_00009_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00009 == conv_Sgntin_row_00009_00004 ) begin
                    conv_qin_00009_00004  <= tout_00009_00004;
                    sign_qin_00009_00004  <=  0;
                end else begin
                    conv_qin_00009_00004  <=  ~tout_00009_00004 + 1;
                    sign_qin_00009_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00009 == conv_Sgntin_row_00009_00005 ) begin
                    conv_qin_00009_00005  <= tout_00009_00005;
                    sign_qin_00009_00005  <=  0;
                end else begin
                    conv_qin_00009_00005  <=  ~tout_00009_00005 + 1;
                    sign_qin_00009_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00009 == conv_Sgntin_row_00009_00006 ) begin
                    conv_qin_00009_00006  <= tout_00009_00006;
                    sign_qin_00009_00006  <=  0;
                end else begin
                    conv_qin_00009_00006  <=  ~tout_00009_00006 + 1;
                    sign_qin_00009_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00009 == conv_Sgntin_row_00009_00007 ) begin
                    conv_qin_00009_00007  <= tout_00009_00007;
                    sign_qin_00009_00007  <=  0;
                end else begin
                    conv_qin_00009_00007  <=  ~tout_00009_00007 + 1;
                    sign_qin_00009_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00010 == conv_Sgntin_row_00010_00000 ) begin
                    conv_qin_00010_00000  <= tout_00010_00000;
                    sign_qin_00010_00000  <=  0;
                end else begin
                    conv_qin_00010_00000  <=  ~tout_00010_00000 + 1;
                    sign_qin_00010_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00010 == conv_Sgntin_row_00010_00001 ) begin
                    conv_qin_00010_00001  <= tout_00010_00001;
                    sign_qin_00010_00001  <=  0;
                end else begin
                    conv_qin_00010_00001  <=  ~tout_00010_00001 + 1;
                    sign_qin_00010_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00010 == conv_Sgntin_row_00010_00002 ) begin
                    conv_qin_00010_00002  <= tout_00010_00002;
                    sign_qin_00010_00002  <=  0;
                end else begin
                    conv_qin_00010_00002  <=  ~tout_00010_00002 + 1;
                    sign_qin_00010_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00010 == conv_Sgntin_row_00010_00003 ) begin
                    conv_qin_00010_00003  <= tout_00010_00003;
                    sign_qin_00010_00003  <=  0;
                end else begin
                    conv_qin_00010_00003  <=  ~tout_00010_00003 + 1;
                    sign_qin_00010_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00010 == conv_Sgntin_row_00010_00004 ) begin
                    conv_qin_00010_00004  <= tout_00010_00004;
                    sign_qin_00010_00004  <=  0;
                end else begin
                    conv_qin_00010_00004  <=  ~tout_00010_00004 + 1;
                    sign_qin_00010_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00010 == conv_Sgntin_row_00010_00005 ) begin
                    conv_qin_00010_00005  <= tout_00010_00005;
                    sign_qin_00010_00005  <=  0;
                end else begin
                    conv_qin_00010_00005  <=  ~tout_00010_00005 + 1;
                    sign_qin_00010_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00010 == conv_Sgntin_row_00010_00006 ) begin
                    conv_qin_00010_00006  <= tout_00010_00006;
                    sign_qin_00010_00006  <=  0;
                end else begin
                    conv_qin_00010_00006  <=  ~tout_00010_00006 + 1;
                    sign_qin_00010_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00010 == conv_Sgntin_row_00010_00007 ) begin
                    conv_qin_00010_00007  <= tout_00010_00007;
                    sign_qin_00010_00007  <=  0;
                end else begin
                    conv_qin_00010_00007  <=  ~tout_00010_00007 + 1;
                    sign_qin_00010_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00011 == conv_Sgntin_row_00011_00000 ) begin
                    conv_qin_00011_00000  <= tout_00011_00000;
                    sign_qin_00011_00000  <=  0;
                end else begin
                    conv_qin_00011_00000  <=  ~tout_00011_00000 + 1;
                    sign_qin_00011_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00011 == conv_Sgntin_row_00011_00001 ) begin
                    conv_qin_00011_00001  <= tout_00011_00001;
                    sign_qin_00011_00001  <=  0;
                end else begin
                    conv_qin_00011_00001  <=  ~tout_00011_00001 + 1;
                    sign_qin_00011_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00011 == conv_Sgntin_row_00011_00002 ) begin
                    conv_qin_00011_00002  <= tout_00011_00002;
                    sign_qin_00011_00002  <=  0;
                end else begin
                    conv_qin_00011_00002  <=  ~tout_00011_00002 + 1;
                    sign_qin_00011_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00011 == conv_Sgntin_row_00011_00003 ) begin
                    conv_qin_00011_00003  <= tout_00011_00003;
                    sign_qin_00011_00003  <=  0;
                end else begin
                    conv_qin_00011_00003  <=  ~tout_00011_00003 + 1;
                    sign_qin_00011_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00011 == conv_Sgntin_row_00011_00004 ) begin
                    conv_qin_00011_00004  <= tout_00011_00004;
                    sign_qin_00011_00004  <=  0;
                end else begin
                    conv_qin_00011_00004  <=  ~tout_00011_00004 + 1;
                    sign_qin_00011_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00011 == conv_Sgntin_row_00011_00005 ) begin
                    conv_qin_00011_00005  <= tout_00011_00005;
                    sign_qin_00011_00005  <=  0;
                end else begin
                    conv_qin_00011_00005  <=  ~tout_00011_00005 + 1;
                    sign_qin_00011_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00011 == conv_Sgntin_row_00011_00006 ) begin
                    conv_qin_00011_00006  <= tout_00011_00006;
                    sign_qin_00011_00006  <=  0;
                end else begin
                    conv_qin_00011_00006  <=  ~tout_00011_00006 + 1;
                    sign_qin_00011_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00011 == conv_Sgntin_row_00011_00007 ) begin
                    conv_qin_00011_00007  <= tout_00011_00007;
                    sign_qin_00011_00007  <=  0;
                end else begin
                    conv_qin_00011_00007  <=  ~tout_00011_00007 + 1;
                    sign_qin_00011_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00012 == conv_Sgntin_row_00012_00000 ) begin
                    conv_qin_00012_00000  <= tout_00012_00000;
                    sign_qin_00012_00000  <=  0;
                end else begin
                    conv_qin_00012_00000  <=  ~tout_00012_00000 + 1;
                    sign_qin_00012_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00012 == conv_Sgntin_row_00012_00001 ) begin
                    conv_qin_00012_00001  <= tout_00012_00001;
                    sign_qin_00012_00001  <=  0;
                end else begin
                    conv_qin_00012_00001  <=  ~tout_00012_00001 + 1;
                    sign_qin_00012_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00012 == conv_Sgntin_row_00012_00002 ) begin
                    conv_qin_00012_00002  <= tout_00012_00002;
                    sign_qin_00012_00002  <=  0;
                end else begin
                    conv_qin_00012_00002  <=  ~tout_00012_00002 + 1;
                    sign_qin_00012_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00012 == conv_Sgntin_row_00012_00003 ) begin
                    conv_qin_00012_00003  <= tout_00012_00003;
                    sign_qin_00012_00003  <=  0;
                end else begin
                    conv_qin_00012_00003  <=  ~tout_00012_00003 + 1;
                    sign_qin_00012_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00012 == conv_Sgntin_row_00012_00004 ) begin
                    conv_qin_00012_00004  <= tout_00012_00004;
                    sign_qin_00012_00004  <=  0;
                end else begin
                    conv_qin_00012_00004  <=  ~tout_00012_00004 + 1;
                    sign_qin_00012_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00012 == conv_Sgntin_row_00012_00005 ) begin
                    conv_qin_00012_00005  <= tout_00012_00005;
                    sign_qin_00012_00005  <=  0;
                end else begin
                    conv_qin_00012_00005  <=  ~tout_00012_00005 + 1;
                    sign_qin_00012_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00012 == conv_Sgntin_row_00012_00006 ) begin
                    conv_qin_00012_00006  <= tout_00012_00006;
                    sign_qin_00012_00006  <=  0;
                end else begin
                    conv_qin_00012_00006  <=  ~tout_00012_00006 + 1;
                    sign_qin_00012_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00012 == conv_Sgntin_row_00012_00007 ) begin
                    conv_qin_00012_00007  <= tout_00012_00007;
                    sign_qin_00012_00007  <=  0;
                end else begin
                    conv_qin_00012_00007  <=  ~tout_00012_00007 + 1;
                    sign_qin_00012_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00012 == conv_Sgntin_row_00012_00008 ) begin
                    conv_qin_00012_00008  <= tout_00012_00008;
                    sign_qin_00012_00008  <=  0;
                end else begin
                    conv_qin_00012_00008  <=  ~tout_00012_00008 + 1;
                    sign_qin_00012_00008  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00012 == conv_Sgntin_row_00012_00009 ) begin
                    conv_qin_00012_00009  <= tout_00012_00009;
                    sign_qin_00012_00009  <=  0;
                end else begin
                    conv_qin_00012_00009  <=  ~tout_00012_00009 + 1;
                    sign_qin_00012_00009  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00013 == conv_Sgntin_row_00013_00000 ) begin
                    conv_qin_00013_00000  <= tout_00013_00000;
                    sign_qin_00013_00000  <=  0;
                end else begin
                    conv_qin_00013_00000  <=  ~tout_00013_00000 + 1;
                    sign_qin_00013_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00013 == conv_Sgntin_row_00013_00001 ) begin
                    conv_qin_00013_00001  <= tout_00013_00001;
                    sign_qin_00013_00001  <=  0;
                end else begin
                    conv_qin_00013_00001  <=  ~tout_00013_00001 + 1;
                    sign_qin_00013_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00013 == conv_Sgntin_row_00013_00002 ) begin
                    conv_qin_00013_00002  <= tout_00013_00002;
                    sign_qin_00013_00002  <=  0;
                end else begin
                    conv_qin_00013_00002  <=  ~tout_00013_00002 + 1;
                    sign_qin_00013_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00013 == conv_Sgntin_row_00013_00003 ) begin
                    conv_qin_00013_00003  <= tout_00013_00003;
                    sign_qin_00013_00003  <=  0;
                end else begin
                    conv_qin_00013_00003  <=  ~tout_00013_00003 + 1;
                    sign_qin_00013_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00013 == conv_Sgntin_row_00013_00004 ) begin
                    conv_qin_00013_00004  <= tout_00013_00004;
                    sign_qin_00013_00004  <=  0;
                end else begin
                    conv_qin_00013_00004  <=  ~tout_00013_00004 + 1;
                    sign_qin_00013_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00013 == conv_Sgntin_row_00013_00005 ) begin
                    conv_qin_00013_00005  <= tout_00013_00005;
                    sign_qin_00013_00005  <=  0;
                end else begin
                    conv_qin_00013_00005  <=  ~tout_00013_00005 + 1;
                    sign_qin_00013_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00013 == conv_Sgntin_row_00013_00006 ) begin
                    conv_qin_00013_00006  <= tout_00013_00006;
                    sign_qin_00013_00006  <=  0;
                end else begin
                    conv_qin_00013_00006  <=  ~tout_00013_00006 + 1;
                    sign_qin_00013_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00013 == conv_Sgntin_row_00013_00007 ) begin
                    conv_qin_00013_00007  <= tout_00013_00007;
                    sign_qin_00013_00007  <=  0;
                end else begin
                    conv_qin_00013_00007  <=  ~tout_00013_00007 + 1;
                    sign_qin_00013_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00013 == conv_Sgntin_row_00013_00008 ) begin
                    conv_qin_00013_00008  <= tout_00013_00008;
                    sign_qin_00013_00008  <=  0;
                end else begin
                    conv_qin_00013_00008  <=  ~tout_00013_00008 + 1;
                    sign_qin_00013_00008  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00013 == conv_Sgntin_row_00013_00009 ) begin
                    conv_qin_00013_00009  <= tout_00013_00009;
                    sign_qin_00013_00009  <=  0;
                end else begin
                    conv_qin_00013_00009  <=  ~tout_00013_00009 + 1;
                    sign_qin_00013_00009  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00014 == conv_Sgntin_row_00014_00000 ) begin
                    conv_qin_00014_00000  <= tout_00014_00000;
                    sign_qin_00014_00000  <=  0;
                end else begin
                    conv_qin_00014_00000  <=  ~tout_00014_00000 + 1;
                    sign_qin_00014_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00014 == conv_Sgntin_row_00014_00001 ) begin
                    conv_qin_00014_00001  <= tout_00014_00001;
                    sign_qin_00014_00001  <=  0;
                end else begin
                    conv_qin_00014_00001  <=  ~tout_00014_00001 + 1;
                    sign_qin_00014_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00014 == conv_Sgntin_row_00014_00002 ) begin
                    conv_qin_00014_00002  <= tout_00014_00002;
                    sign_qin_00014_00002  <=  0;
                end else begin
                    conv_qin_00014_00002  <=  ~tout_00014_00002 + 1;
                    sign_qin_00014_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00014 == conv_Sgntin_row_00014_00003 ) begin
                    conv_qin_00014_00003  <= tout_00014_00003;
                    sign_qin_00014_00003  <=  0;
                end else begin
                    conv_qin_00014_00003  <=  ~tout_00014_00003 + 1;
                    sign_qin_00014_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00014 == conv_Sgntin_row_00014_00004 ) begin
                    conv_qin_00014_00004  <= tout_00014_00004;
                    sign_qin_00014_00004  <=  0;
                end else begin
                    conv_qin_00014_00004  <=  ~tout_00014_00004 + 1;
                    sign_qin_00014_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00014 == conv_Sgntin_row_00014_00005 ) begin
                    conv_qin_00014_00005  <= tout_00014_00005;
                    sign_qin_00014_00005  <=  0;
                end else begin
                    conv_qin_00014_00005  <=  ~tout_00014_00005 + 1;
                    sign_qin_00014_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00014 == conv_Sgntin_row_00014_00006 ) begin
                    conv_qin_00014_00006  <= tout_00014_00006;
                    sign_qin_00014_00006  <=  0;
                end else begin
                    conv_qin_00014_00006  <=  ~tout_00014_00006 + 1;
                    sign_qin_00014_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00014 == conv_Sgntin_row_00014_00007 ) begin
                    conv_qin_00014_00007  <= tout_00014_00007;
                    sign_qin_00014_00007  <=  0;
                end else begin
                    conv_qin_00014_00007  <=  ~tout_00014_00007 + 1;
                    sign_qin_00014_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00014 == conv_Sgntin_row_00014_00008 ) begin
                    conv_qin_00014_00008  <= tout_00014_00008;
                    sign_qin_00014_00008  <=  0;
                end else begin
                    conv_qin_00014_00008  <=  ~tout_00014_00008 + 1;
                    sign_qin_00014_00008  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00014 == conv_Sgntin_row_00014_00009 ) begin
                    conv_qin_00014_00009  <= tout_00014_00009;
                    sign_qin_00014_00009  <=  0;
                end else begin
                    conv_qin_00014_00009  <=  ~tout_00014_00009 + 1;
                    sign_qin_00014_00009  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00015 == conv_Sgntin_row_00015_00000 ) begin
                    conv_qin_00015_00000  <= tout_00015_00000;
                    sign_qin_00015_00000  <=  0;
                end else begin
                    conv_qin_00015_00000  <=  ~tout_00015_00000 + 1;
                    sign_qin_00015_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00015 == conv_Sgntin_row_00015_00001 ) begin
                    conv_qin_00015_00001  <= tout_00015_00001;
                    sign_qin_00015_00001  <=  0;
                end else begin
                    conv_qin_00015_00001  <=  ~tout_00015_00001 + 1;
                    sign_qin_00015_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00015 == conv_Sgntin_row_00015_00002 ) begin
                    conv_qin_00015_00002  <= tout_00015_00002;
                    sign_qin_00015_00002  <=  0;
                end else begin
                    conv_qin_00015_00002  <=  ~tout_00015_00002 + 1;
                    sign_qin_00015_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00015 == conv_Sgntin_row_00015_00003 ) begin
                    conv_qin_00015_00003  <= tout_00015_00003;
                    sign_qin_00015_00003  <=  0;
                end else begin
                    conv_qin_00015_00003  <=  ~tout_00015_00003 + 1;
                    sign_qin_00015_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00015 == conv_Sgntin_row_00015_00004 ) begin
                    conv_qin_00015_00004  <= tout_00015_00004;
                    sign_qin_00015_00004  <=  0;
                end else begin
                    conv_qin_00015_00004  <=  ~tout_00015_00004 + 1;
                    sign_qin_00015_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00015 == conv_Sgntin_row_00015_00005 ) begin
                    conv_qin_00015_00005  <= tout_00015_00005;
                    sign_qin_00015_00005  <=  0;
                end else begin
                    conv_qin_00015_00005  <=  ~tout_00015_00005 + 1;
                    sign_qin_00015_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00015 == conv_Sgntin_row_00015_00006 ) begin
                    conv_qin_00015_00006  <= tout_00015_00006;
                    sign_qin_00015_00006  <=  0;
                end else begin
                    conv_qin_00015_00006  <=  ~tout_00015_00006 + 1;
                    sign_qin_00015_00006  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00015 == conv_Sgntin_row_00015_00007 ) begin
                    conv_qin_00015_00007  <= tout_00015_00007;
                    sign_qin_00015_00007  <=  0;
                end else begin
                    conv_qin_00015_00007  <=  ~tout_00015_00007 + 1;
                    sign_qin_00015_00007  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00015 == conv_Sgntin_row_00015_00008 ) begin
                    conv_qin_00015_00008  <= tout_00015_00008;
                    sign_qin_00015_00008  <=  0;
                end else begin
                    conv_qin_00015_00008  <=  ~tout_00015_00008 + 1;
                    sign_qin_00015_00008  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00015 == conv_Sgntin_row_00015_00009 ) begin
                    conv_qin_00015_00009  <= tout_00015_00009;
                    sign_qin_00015_00009  <=  0;
                end else begin
                    conv_qin_00015_00009  <=  ~tout_00015_00009 + 1;
                    sign_qin_00015_00009  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00016 == conv_Sgntin_row_00016_00000 ) begin
                    conv_qin_00016_00000  <= tout_00016_00000;
                    sign_qin_00016_00000  <=  0;
                end else begin
                    conv_qin_00016_00000  <=  ~tout_00016_00000 + 1;
                    sign_qin_00016_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00016 == conv_Sgntin_row_00016_00001 ) begin
                    conv_qin_00016_00001  <= tout_00016_00001;
                    sign_qin_00016_00001  <=  0;
                end else begin
                    conv_qin_00016_00001  <=  ~tout_00016_00001 + 1;
                    sign_qin_00016_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00016 == conv_Sgntin_row_00016_00002 ) begin
                    conv_qin_00016_00002  <= tout_00016_00002;
                    sign_qin_00016_00002  <=  0;
                end else begin
                    conv_qin_00016_00002  <=  ~tout_00016_00002 + 1;
                    sign_qin_00016_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00016 == conv_Sgntin_row_00016_00003 ) begin
                    conv_qin_00016_00003  <= tout_00016_00003;
                    sign_qin_00016_00003  <=  0;
                end else begin
                    conv_qin_00016_00003  <=  ~tout_00016_00003 + 1;
                    sign_qin_00016_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00017 == conv_Sgntin_row_00017_00000 ) begin
                    conv_qin_00017_00000  <= tout_00017_00000;
                    sign_qin_00017_00000  <=  0;
                end else begin
                    conv_qin_00017_00000  <=  ~tout_00017_00000 + 1;
                    sign_qin_00017_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00017 == conv_Sgntin_row_00017_00001 ) begin
                    conv_qin_00017_00001  <= tout_00017_00001;
                    sign_qin_00017_00001  <=  0;
                end else begin
                    conv_qin_00017_00001  <=  ~tout_00017_00001 + 1;
                    sign_qin_00017_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00017 == conv_Sgntin_row_00017_00002 ) begin
                    conv_qin_00017_00002  <= tout_00017_00002;
                    sign_qin_00017_00002  <=  0;
                end else begin
                    conv_qin_00017_00002  <=  ~tout_00017_00002 + 1;
                    sign_qin_00017_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00017 == conv_Sgntin_row_00017_00003 ) begin
                    conv_qin_00017_00003  <= tout_00017_00003;
                    sign_qin_00017_00003  <=  0;
                end else begin
                    conv_qin_00017_00003  <=  ~tout_00017_00003 + 1;
                    sign_qin_00017_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00018 == conv_Sgntin_row_00018_00000 ) begin
                    conv_qin_00018_00000  <= tout_00018_00000;
                    sign_qin_00018_00000  <=  0;
                end else begin
                    conv_qin_00018_00000  <=  ~tout_00018_00000 + 1;
                    sign_qin_00018_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00018 == conv_Sgntin_row_00018_00001 ) begin
                    conv_qin_00018_00001  <= tout_00018_00001;
                    sign_qin_00018_00001  <=  0;
                end else begin
                    conv_qin_00018_00001  <=  ~tout_00018_00001 + 1;
                    sign_qin_00018_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00018 == conv_Sgntin_row_00018_00002 ) begin
                    conv_qin_00018_00002  <= tout_00018_00002;
                    sign_qin_00018_00002  <=  0;
                end else begin
                    conv_qin_00018_00002  <=  ~tout_00018_00002 + 1;
                    sign_qin_00018_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00018 == conv_Sgntin_row_00018_00003 ) begin
                    conv_qin_00018_00003  <= tout_00018_00003;
                    sign_qin_00018_00003  <=  0;
                end else begin
                    conv_qin_00018_00003  <=  ~tout_00018_00003 + 1;
                    sign_qin_00018_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00019 == conv_Sgntin_row_00019_00000 ) begin
                    conv_qin_00019_00000  <= tout_00019_00000;
                    sign_qin_00019_00000  <=  0;
                end else begin
                    conv_qin_00019_00000  <=  ~tout_00019_00000 + 1;
                    sign_qin_00019_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00019 == conv_Sgntin_row_00019_00001 ) begin
                    conv_qin_00019_00001  <= tout_00019_00001;
                    sign_qin_00019_00001  <=  0;
                end else begin
                    conv_qin_00019_00001  <=  ~tout_00019_00001 + 1;
                    sign_qin_00019_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00019 == conv_Sgntin_row_00019_00002 ) begin
                    conv_qin_00019_00002  <= tout_00019_00002;
                    sign_qin_00019_00002  <=  0;
                end else begin
                    conv_qin_00019_00002  <=  ~tout_00019_00002 + 1;
                    sign_qin_00019_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00019 == conv_Sgntin_row_00019_00003 ) begin
                    conv_qin_00019_00003  <= tout_00019_00003;
                    sign_qin_00019_00003  <=  0;
                end else begin
                    conv_qin_00019_00003  <=  ~tout_00019_00003 + 1;
                    sign_qin_00019_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00020 == conv_Sgntin_row_00020_00000 ) begin
                    conv_qin_00020_00000  <= tout_00020_00000;
                    sign_qin_00020_00000  <=  0;
                end else begin
                    conv_qin_00020_00000  <=  ~tout_00020_00000 + 1;
                    sign_qin_00020_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00020 == conv_Sgntin_row_00020_00001 ) begin
                    conv_qin_00020_00001  <= tout_00020_00001;
                    sign_qin_00020_00001  <=  0;
                end else begin
                    conv_qin_00020_00001  <=  ~tout_00020_00001 + 1;
                    sign_qin_00020_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00020 == conv_Sgntin_row_00020_00002 ) begin
                    conv_qin_00020_00002  <= tout_00020_00002;
                    sign_qin_00020_00002  <=  0;
                end else begin
                    conv_qin_00020_00002  <=  ~tout_00020_00002 + 1;
                    sign_qin_00020_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00020 == conv_Sgntin_row_00020_00003 ) begin
                    conv_qin_00020_00003  <= tout_00020_00003;
                    sign_qin_00020_00003  <=  0;
                end else begin
                    conv_qin_00020_00003  <=  ~tout_00020_00003 + 1;
                    sign_qin_00020_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00020 == conv_Sgntin_row_00020_00004 ) begin
                    conv_qin_00020_00004  <= tout_00020_00004;
                    sign_qin_00020_00004  <=  0;
                end else begin
                    conv_qin_00020_00004  <=  ~tout_00020_00004 + 1;
                    sign_qin_00020_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00020 == conv_Sgntin_row_00020_00005 ) begin
                    conv_qin_00020_00005  <= tout_00020_00005;
                    sign_qin_00020_00005  <=  0;
                end else begin
                    conv_qin_00020_00005  <=  ~tout_00020_00005 + 1;
                    sign_qin_00020_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00021 == conv_Sgntin_row_00021_00000 ) begin
                    conv_qin_00021_00000  <= tout_00021_00000;
                    sign_qin_00021_00000  <=  0;
                end else begin
                    conv_qin_00021_00000  <=  ~tout_00021_00000 + 1;
                    sign_qin_00021_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00021 == conv_Sgntin_row_00021_00001 ) begin
                    conv_qin_00021_00001  <= tout_00021_00001;
                    sign_qin_00021_00001  <=  0;
                end else begin
                    conv_qin_00021_00001  <=  ~tout_00021_00001 + 1;
                    sign_qin_00021_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00021 == conv_Sgntin_row_00021_00002 ) begin
                    conv_qin_00021_00002  <= tout_00021_00002;
                    sign_qin_00021_00002  <=  0;
                end else begin
                    conv_qin_00021_00002  <=  ~tout_00021_00002 + 1;
                    sign_qin_00021_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00021 == conv_Sgntin_row_00021_00003 ) begin
                    conv_qin_00021_00003  <= tout_00021_00003;
                    sign_qin_00021_00003  <=  0;
                end else begin
                    conv_qin_00021_00003  <=  ~tout_00021_00003 + 1;
                    sign_qin_00021_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00021 == conv_Sgntin_row_00021_00004 ) begin
                    conv_qin_00021_00004  <= tout_00021_00004;
                    sign_qin_00021_00004  <=  0;
                end else begin
                    conv_qin_00021_00004  <=  ~tout_00021_00004 + 1;
                    sign_qin_00021_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00021 == conv_Sgntin_row_00021_00005 ) begin
                    conv_qin_00021_00005  <= tout_00021_00005;
                    sign_qin_00021_00005  <=  0;
                end else begin
                    conv_qin_00021_00005  <=  ~tout_00021_00005 + 1;
                    sign_qin_00021_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00022 == conv_Sgntin_row_00022_00000 ) begin
                    conv_qin_00022_00000  <= tout_00022_00000;
                    sign_qin_00022_00000  <=  0;
                end else begin
                    conv_qin_00022_00000  <=  ~tout_00022_00000 + 1;
                    sign_qin_00022_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00022 == conv_Sgntin_row_00022_00001 ) begin
                    conv_qin_00022_00001  <= tout_00022_00001;
                    sign_qin_00022_00001  <=  0;
                end else begin
                    conv_qin_00022_00001  <=  ~tout_00022_00001 + 1;
                    sign_qin_00022_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00022 == conv_Sgntin_row_00022_00002 ) begin
                    conv_qin_00022_00002  <= tout_00022_00002;
                    sign_qin_00022_00002  <=  0;
                end else begin
                    conv_qin_00022_00002  <=  ~tout_00022_00002 + 1;
                    sign_qin_00022_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00022 == conv_Sgntin_row_00022_00003 ) begin
                    conv_qin_00022_00003  <= tout_00022_00003;
                    sign_qin_00022_00003  <=  0;
                end else begin
                    conv_qin_00022_00003  <=  ~tout_00022_00003 + 1;
                    sign_qin_00022_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00022 == conv_Sgntin_row_00022_00004 ) begin
                    conv_qin_00022_00004  <= tout_00022_00004;
                    sign_qin_00022_00004  <=  0;
                end else begin
                    conv_qin_00022_00004  <=  ~tout_00022_00004 + 1;
                    sign_qin_00022_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00022 == conv_Sgntin_row_00022_00005 ) begin
                    conv_qin_00022_00005  <= tout_00022_00005;
                    sign_qin_00022_00005  <=  0;
                end else begin
                    conv_qin_00022_00005  <=  ~tout_00022_00005 + 1;
                    sign_qin_00022_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00023 == conv_Sgntin_row_00023_00000 ) begin
                    conv_qin_00023_00000  <= tout_00023_00000;
                    sign_qin_00023_00000  <=  0;
                end else begin
                    conv_qin_00023_00000  <=  ~tout_00023_00000 + 1;
                    sign_qin_00023_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00023 == conv_Sgntin_row_00023_00001 ) begin
                    conv_qin_00023_00001  <= tout_00023_00001;
                    sign_qin_00023_00001  <=  0;
                end else begin
                    conv_qin_00023_00001  <=  ~tout_00023_00001 + 1;
                    sign_qin_00023_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00023 == conv_Sgntin_row_00023_00002 ) begin
                    conv_qin_00023_00002  <= tout_00023_00002;
                    sign_qin_00023_00002  <=  0;
                end else begin
                    conv_qin_00023_00002  <=  ~tout_00023_00002 + 1;
                    sign_qin_00023_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00023 == conv_Sgntin_row_00023_00003 ) begin
                    conv_qin_00023_00003  <= tout_00023_00003;
                    sign_qin_00023_00003  <=  0;
                end else begin
                    conv_qin_00023_00003  <=  ~tout_00023_00003 + 1;
                    sign_qin_00023_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00023 == conv_Sgntin_row_00023_00004 ) begin
                    conv_qin_00023_00004  <= tout_00023_00004;
                    sign_qin_00023_00004  <=  0;
                end else begin
                    conv_qin_00023_00004  <=  ~tout_00023_00004 + 1;
                    sign_qin_00023_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00023 == conv_Sgntin_row_00023_00005 ) begin
                    conv_qin_00023_00005  <= tout_00023_00005;
                    sign_qin_00023_00005  <=  0;
                end else begin
                    conv_qin_00023_00005  <=  ~tout_00023_00005 + 1;
                    sign_qin_00023_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00024 == conv_Sgntin_row_00024_00000 ) begin
                    conv_qin_00024_00000  <= tout_00024_00000;
                    sign_qin_00024_00000  <=  0;
                end else begin
                    conv_qin_00024_00000  <=  ~tout_00024_00000 + 1;
                    sign_qin_00024_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00024 == conv_Sgntin_row_00024_00001 ) begin
                    conv_qin_00024_00001  <= tout_00024_00001;
                    sign_qin_00024_00001  <=  0;
                end else begin
                    conv_qin_00024_00001  <=  ~tout_00024_00001 + 1;
                    sign_qin_00024_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00024 == conv_Sgntin_row_00024_00002 ) begin
                    conv_qin_00024_00002  <= tout_00024_00002;
                    sign_qin_00024_00002  <=  0;
                end else begin
                    conv_qin_00024_00002  <=  ~tout_00024_00002 + 1;
                    sign_qin_00024_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00024 == conv_Sgntin_row_00024_00003 ) begin
                    conv_qin_00024_00003  <= tout_00024_00003;
                    sign_qin_00024_00003  <=  0;
                end else begin
                    conv_qin_00024_00003  <=  ~tout_00024_00003 + 1;
                    sign_qin_00024_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00024 == conv_Sgntin_row_00024_00004 ) begin
                    conv_qin_00024_00004  <= tout_00024_00004;
                    sign_qin_00024_00004  <=  0;
                end else begin
                    conv_qin_00024_00004  <=  ~tout_00024_00004 + 1;
                    sign_qin_00024_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00024 == conv_Sgntin_row_00024_00005 ) begin
                    conv_qin_00024_00005  <= tout_00024_00005;
                    sign_qin_00024_00005  <=  0;
                end else begin
                    conv_qin_00024_00005  <=  ~tout_00024_00005 + 1;
                    sign_qin_00024_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00025 == conv_Sgntin_row_00025_00000 ) begin
                    conv_qin_00025_00000  <= tout_00025_00000;
                    sign_qin_00025_00000  <=  0;
                end else begin
                    conv_qin_00025_00000  <=  ~tout_00025_00000 + 1;
                    sign_qin_00025_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00025 == conv_Sgntin_row_00025_00001 ) begin
                    conv_qin_00025_00001  <= tout_00025_00001;
                    sign_qin_00025_00001  <=  0;
                end else begin
                    conv_qin_00025_00001  <=  ~tout_00025_00001 + 1;
                    sign_qin_00025_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00025 == conv_Sgntin_row_00025_00002 ) begin
                    conv_qin_00025_00002  <= tout_00025_00002;
                    sign_qin_00025_00002  <=  0;
                end else begin
                    conv_qin_00025_00002  <=  ~tout_00025_00002 + 1;
                    sign_qin_00025_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00025 == conv_Sgntin_row_00025_00003 ) begin
                    conv_qin_00025_00003  <= tout_00025_00003;
                    sign_qin_00025_00003  <=  0;
                end else begin
                    conv_qin_00025_00003  <=  ~tout_00025_00003 + 1;
                    sign_qin_00025_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00025 == conv_Sgntin_row_00025_00004 ) begin
                    conv_qin_00025_00004  <= tout_00025_00004;
                    sign_qin_00025_00004  <=  0;
                end else begin
                    conv_qin_00025_00004  <=  ~tout_00025_00004 + 1;
                    sign_qin_00025_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00025 == conv_Sgntin_row_00025_00005 ) begin
                    conv_qin_00025_00005  <= tout_00025_00005;
                    sign_qin_00025_00005  <=  0;
                end else begin
                    conv_qin_00025_00005  <=  ~tout_00025_00005 + 1;
                    sign_qin_00025_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00026 == conv_Sgntin_row_00026_00000 ) begin
                    conv_qin_00026_00000  <= tout_00026_00000;
                    sign_qin_00026_00000  <=  0;
                end else begin
                    conv_qin_00026_00000  <=  ~tout_00026_00000 + 1;
                    sign_qin_00026_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00026 == conv_Sgntin_row_00026_00001 ) begin
                    conv_qin_00026_00001  <= tout_00026_00001;
                    sign_qin_00026_00001  <=  0;
                end else begin
                    conv_qin_00026_00001  <=  ~tout_00026_00001 + 1;
                    sign_qin_00026_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00026 == conv_Sgntin_row_00026_00002 ) begin
                    conv_qin_00026_00002  <= tout_00026_00002;
                    sign_qin_00026_00002  <=  0;
                end else begin
                    conv_qin_00026_00002  <=  ~tout_00026_00002 + 1;
                    sign_qin_00026_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00026 == conv_Sgntin_row_00026_00003 ) begin
                    conv_qin_00026_00003  <= tout_00026_00003;
                    sign_qin_00026_00003  <=  0;
                end else begin
                    conv_qin_00026_00003  <=  ~tout_00026_00003 + 1;
                    sign_qin_00026_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00026 == conv_Sgntin_row_00026_00004 ) begin
                    conv_qin_00026_00004  <= tout_00026_00004;
                    sign_qin_00026_00004  <=  0;
                end else begin
                    conv_qin_00026_00004  <=  ~tout_00026_00004 + 1;
                    sign_qin_00026_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00026 == conv_Sgntin_row_00026_00005 ) begin
                    conv_qin_00026_00005  <= tout_00026_00005;
                    sign_qin_00026_00005  <=  0;
                end else begin
                    conv_qin_00026_00005  <=  ~tout_00026_00005 + 1;
                    sign_qin_00026_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00027 == conv_Sgntin_row_00027_00000 ) begin
                    conv_qin_00027_00000  <= tout_00027_00000;
                    sign_qin_00027_00000  <=  0;
                end else begin
                    conv_qin_00027_00000  <=  ~tout_00027_00000 + 1;
                    sign_qin_00027_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00027 == conv_Sgntin_row_00027_00001 ) begin
                    conv_qin_00027_00001  <= tout_00027_00001;
                    sign_qin_00027_00001  <=  0;
                end else begin
                    conv_qin_00027_00001  <=  ~tout_00027_00001 + 1;
                    sign_qin_00027_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00027 == conv_Sgntin_row_00027_00002 ) begin
                    conv_qin_00027_00002  <= tout_00027_00002;
                    sign_qin_00027_00002  <=  0;
                end else begin
                    conv_qin_00027_00002  <=  ~tout_00027_00002 + 1;
                    sign_qin_00027_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00027 == conv_Sgntin_row_00027_00003 ) begin
                    conv_qin_00027_00003  <= tout_00027_00003;
                    sign_qin_00027_00003  <=  0;
                end else begin
                    conv_qin_00027_00003  <=  ~tout_00027_00003 + 1;
                    sign_qin_00027_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00027 == conv_Sgntin_row_00027_00004 ) begin
                    conv_qin_00027_00004  <= tout_00027_00004;
                    sign_qin_00027_00004  <=  0;
                end else begin
                    conv_qin_00027_00004  <=  ~tout_00027_00004 + 1;
                    sign_qin_00027_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00027 == conv_Sgntin_row_00027_00005 ) begin
                    conv_qin_00027_00005  <= tout_00027_00005;
                    sign_qin_00027_00005  <=  0;
                end else begin
                    conv_qin_00027_00005  <=  ~tout_00027_00005 + 1;
                    sign_qin_00027_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00028 == conv_Sgntin_row_00028_00000 ) begin
                    conv_qin_00028_00000  <= tout_00028_00000;
                    sign_qin_00028_00000  <=  0;
                end else begin
                    conv_qin_00028_00000  <=  ~tout_00028_00000 + 1;
                    sign_qin_00028_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00028 == conv_Sgntin_row_00028_00001 ) begin
                    conv_qin_00028_00001  <= tout_00028_00001;
                    sign_qin_00028_00001  <=  0;
                end else begin
                    conv_qin_00028_00001  <=  ~tout_00028_00001 + 1;
                    sign_qin_00028_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00028 == conv_Sgntin_row_00028_00002 ) begin
                    conv_qin_00028_00002  <= tout_00028_00002;
                    sign_qin_00028_00002  <=  0;
                end else begin
                    conv_qin_00028_00002  <=  ~tout_00028_00002 + 1;
                    sign_qin_00028_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00028 == conv_Sgntin_row_00028_00003 ) begin
                    conv_qin_00028_00003  <= tout_00028_00003;
                    sign_qin_00028_00003  <=  0;
                end else begin
                    conv_qin_00028_00003  <=  ~tout_00028_00003 + 1;
                    sign_qin_00028_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00028 == conv_Sgntin_row_00028_00004 ) begin
                    conv_qin_00028_00004  <= tout_00028_00004;
                    sign_qin_00028_00004  <=  0;
                end else begin
                    conv_qin_00028_00004  <=  ~tout_00028_00004 + 1;
                    sign_qin_00028_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00028 == conv_Sgntin_row_00028_00005 ) begin
                    conv_qin_00028_00005  <= tout_00028_00005;
                    sign_qin_00028_00005  <=  0;
                end else begin
                    conv_qin_00028_00005  <=  ~tout_00028_00005 + 1;
                    sign_qin_00028_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00029 == conv_Sgntin_row_00029_00000 ) begin
                    conv_qin_00029_00000  <= tout_00029_00000;
                    sign_qin_00029_00000  <=  0;
                end else begin
                    conv_qin_00029_00000  <=  ~tout_00029_00000 + 1;
                    sign_qin_00029_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00029 == conv_Sgntin_row_00029_00001 ) begin
                    conv_qin_00029_00001  <= tout_00029_00001;
                    sign_qin_00029_00001  <=  0;
                end else begin
                    conv_qin_00029_00001  <=  ~tout_00029_00001 + 1;
                    sign_qin_00029_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00029 == conv_Sgntin_row_00029_00002 ) begin
                    conv_qin_00029_00002  <= tout_00029_00002;
                    sign_qin_00029_00002  <=  0;
                end else begin
                    conv_qin_00029_00002  <=  ~tout_00029_00002 + 1;
                    sign_qin_00029_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00029 == conv_Sgntin_row_00029_00003 ) begin
                    conv_qin_00029_00003  <= tout_00029_00003;
                    sign_qin_00029_00003  <=  0;
                end else begin
                    conv_qin_00029_00003  <=  ~tout_00029_00003 + 1;
                    sign_qin_00029_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00029 == conv_Sgntin_row_00029_00004 ) begin
                    conv_qin_00029_00004  <= tout_00029_00004;
                    sign_qin_00029_00004  <=  0;
                end else begin
                    conv_qin_00029_00004  <=  ~tout_00029_00004 + 1;
                    sign_qin_00029_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00029 == conv_Sgntin_row_00029_00005 ) begin
                    conv_qin_00029_00005  <= tout_00029_00005;
                    sign_qin_00029_00005  <=  0;
                end else begin
                    conv_qin_00029_00005  <=  ~tout_00029_00005 + 1;
                    sign_qin_00029_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00030 == conv_Sgntin_row_00030_00000 ) begin
                    conv_qin_00030_00000  <= tout_00030_00000;
                    sign_qin_00030_00000  <=  0;
                end else begin
                    conv_qin_00030_00000  <=  ~tout_00030_00000 + 1;
                    sign_qin_00030_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00030 == conv_Sgntin_row_00030_00001 ) begin
                    conv_qin_00030_00001  <= tout_00030_00001;
                    sign_qin_00030_00001  <=  0;
                end else begin
                    conv_qin_00030_00001  <=  ~tout_00030_00001 + 1;
                    sign_qin_00030_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00030 == conv_Sgntin_row_00030_00002 ) begin
                    conv_qin_00030_00002  <= tout_00030_00002;
                    sign_qin_00030_00002  <=  0;
                end else begin
                    conv_qin_00030_00002  <=  ~tout_00030_00002 + 1;
                    sign_qin_00030_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00030 == conv_Sgntin_row_00030_00003 ) begin
                    conv_qin_00030_00003  <= tout_00030_00003;
                    sign_qin_00030_00003  <=  0;
                end else begin
                    conv_qin_00030_00003  <=  ~tout_00030_00003 + 1;
                    sign_qin_00030_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00030 == conv_Sgntin_row_00030_00004 ) begin
                    conv_qin_00030_00004  <= tout_00030_00004;
                    sign_qin_00030_00004  <=  0;
                end else begin
                    conv_qin_00030_00004  <=  ~tout_00030_00004 + 1;
                    sign_qin_00030_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00030 == conv_Sgntin_row_00030_00005 ) begin
                    conv_qin_00030_00005  <= tout_00030_00005;
                    sign_qin_00030_00005  <=  0;
                end else begin
                    conv_qin_00030_00005  <=  ~tout_00030_00005 + 1;
                    sign_qin_00030_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00031 == conv_Sgntin_row_00031_00000 ) begin
                    conv_qin_00031_00000  <= tout_00031_00000;
                    sign_qin_00031_00000  <=  0;
                end else begin
                    conv_qin_00031_00000  <=  ~tout_00031_00000 + 1;
                    sign_qin_00031_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00031 == conv_Sgntin_row_00031_00001 ) begin
                    conv_qin_00031_00001  <= tout_00031_00001;
                    sign_qin_00031_00001  <=  0;
                end else begin
                    conv_qin_00031_00001  <=  ~tout_00031_00001 + 1;
                    sign_qin_00031_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00031 == conv_Sgntin_row_00031_00002 ) begin
                    conv_qin_00031_00002  <= tout_00031_00002;
                    sign_qin_00031_00002  <=  0;
                end else begin
                    conv_qin_00031_00002  <=  ~tout_00031_00002 + 1;
                    sign_qin_00031_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00031 == conv_Sgntin_row_00031_00003 ) begin
                    conv_qin_00031_00003  <= tout_00031_00003;
                    sign_qin_00031_00003  <=  0;
                end else begin
                    conv_qin_00031_00003  <=  ~tout_00031_00003 + 1;
                    sign_qin_00031_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00031 == conv_Sgntin_row_00031_00004 ) begin
                    conv_qin_00031_00004  <= tout_00031_00004;
                    sign_qin_00031_00004  <=  0;
                end else begin
                    conv_qin_00031_00004  <=  ~tout_00031_00004 + 1;
                    sign_qin_00031_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00031 == conv_Sgntin_row_00031_00005 ) begin
                    conv_qin_00031_00005  <= tout_00031_00005;
                    sign_qin_00031_00005  <=  0;
                end else begin
                    conv_qin_00031_00005  <=  ~tout_00031_00005 + 1;
                    sign_qin_00031_00005  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00032 == conv_Sgntin_row_00032_00000 ) begin
                    conv_qin_00032_00000  <= tout_00032_00000;
                    sign_qin_00032_00000  <=  0;
                end else begin
                    conv_qin_00032_00000  <=  ~tout_00032_00000 + 1;
                    sign_qin_00032_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00032 == conv_Sgntin_row_00032_00001 ) begin
                    conv_qin_00032_00001  <= tout_00032_00001;
                    sign_qin_00032_00001  <=  0;
                end else begin
                    conv_qin_00032_00001  <=  ~tout_00032_00001 + 1;
                    sign_qin_00032_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00032 == conv_Sgntin_row_00032_00002 ) begin
                    conv_qin_00032_00002  <= tout_00032_00002;
                    sign_qin_00032_00002  <=  0;
                end else begin
                    conv_qin_00032_00002  <=  ~tout_00032_00002 + 1;
                    sign_qin_00032_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00032 == conv_Sgntin_row_00032_00003 ) begin
                    conv_qin_00032_00003  <= tout_00032_00003;
                    sign_qin_00032_00003  <=  0;
                end else begin
                    conv_qin_00032_00003  <=  ~tout_00032_00003 + 1;
                    sign_qin_00032_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00033 == conv_Sgntin_row_00033_00000 ) begin
                    conv_qin_00033_00000  <= tout_00033_00000;
                    sign_qin_00033_00000  <=  0;
                end else begin
                    conv_qin_00033_00000  <=  ~tout_00033_00000 + 1;
                    sign_qin_00033_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00033 == conv_Sgntin_row_00033_00001 ) begin
                    conv_qin_00033_00001  <= tout_00033_00001;
                    sign_qin_00033_00001  <=  0;
                end else begin
                    conv_qin_00033_00001  <=  ~tout_00033_00001 + 1;
                    sign_qin_00033_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00033 == conv_Sgntin_row_00033_00002 ) begin
                    conv_qin_00033_00002  <= tout_00033_00002;
                    sign_qin_00033_00002  <=  0;
                end else begin
                    conv_qin_00033_00002  <=  ~tout_00033_00002 + 1;
                    sign_qin_00033_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00033 == conv_Sgntin_row_00033_00003 ) begin
                    conv_qin_00033_00003  <= tout_00033_00003;
                    sign_qin_00033_00003  <=  0;
                end else begin
                    conv_qin_00033_00003  <=  ~tout_00033_00003 + 1;
                    sign_qin_00033_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00034 == conv_Sgntin_row_00034_00000 ) begin
                    conv_qin_00034_00000  <= tout_00034_00000;
                    sign_qin_00034_00000  <=  0;
                end else begin
                    conv_qin_00034_00000  <=  ~tout_00034_00000 + 1;
                    sign_qin_00034_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00034 == conv_Sgntin_row_00034_00001 ) begin
                    conv_qin_00034_00001  <= tout_00034_00001;
                    sign_qin_00034_00001  <=  0;
                end else begin
                    conv_qin_00034_00001  <=  ~tout_00034_00001 + 1;
                    sign_qin_00034_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00034 == conv_Sgntin_row_00034_00002 ) begin
                    conv_qin_00034_00002  <= tout_00034_00002;
                    sign_qin_00034_00002  <=  0;
                end else begin
                    conv_qin_00034_00002  <=  ~tout_00034_00002 + 1;
                    sign_qin_00034_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00034 == conv_Sgntin_row_00034_00003 ) begin
                    conv_qin_00034_00003  <= tout_00034_00003;
                    sign_qin_00034_00003  <=  0;
                end else begin
                    conv_qin_00034_00003  <=  ~tout_00034_00003 + 1;
                    sign_qin_00034_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00035 == conv_Sgntin_row_00035_00000 ) begin
                    conv_qin_00035_00000  <= tout_00035_00000;
                    sign_qin_00035_00000  <=  0;
                end else begin
                    conv_qin_00035_00000  <=  ~tout_00035_00000 + 1;
                    sign_qin_00035_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00035 == conv_Sgntin_row_00035_00001 ) begin
                    conv_qin_00035_00001  <= tout_00035_00001;
                    sign_qin_00035_00001  <=  0;
                end else begin
                    conv_qin_00035_00001  <=  ~tout_00035_00001 + 1;
                    sign_qin_00035_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00035 == conv_Sgntin_row_00035_00002 ) begin
                    conv_qin_00035_00002  <= tout_00035_00002;
                    sign_qin_00035_00002  <=  0;
                end else begin
                    conv_qin_00035_00002  <=  ~tout_00035_00002 + 1;
                    sign_qin_00035_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00035 == conv_Sgntin_row_00035_00003 ) begin
                    conv_qin_00035_00003  <= tout_00035_00003;
                    sign_qin_00035_00003  <=  0;
                end else begin
                    conv_qin_00035_00003  <=  ~tout_00035_00003 + 1;
                    sign_qin_00035_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00036 == conv_Sgntin_row_00036_00000 ) begin
                    conv_qin_00036_00000  <= tout_00036_00000;
                    sign_qin_00036_00000  <=  0;
                end else begin
                    conv_qin_00036_00000  <=  ~tout_00036_00000 + 1;
                    sign_qin_00036_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00036 == conv_Sgntin_row_00036_00001 ) begin
                    conv_qin_00036_00001  <= tout_00036_00001;
                    sign_qin_00036_00001  <=  0;
                end else begin
                    conv_qin_00036_00001  <=  ~tout_00036_00001 + 1;
                    sign_qin_00036_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00036 == conv_Sgntin_row_00036_00002 ) begin
                    conv_qin_00036_00002  <= tout_00036_00002;
                    sign_qin_00036_00002  <=  0;
                end else begin
                    conv_qin_00036_00002  <=  ~tout_00036_00002 + 1;
                    sign_qin_00036_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00036 == conv_Sgntin_row_00036_00003 ) begin
                    conv_qin_00036_00003  <= tout_00036_00003;
                    sign_qin_00036_00003  <=  0;
                end else begin
                    conv_qin_00036_00003  <=  ~tout_00036_00003 + 1;
                    sign_qin_00036_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00036 == conv_Sgntin_row_00036_00004 ) begin
                    conv_qin_00036_00004  <= tout_00036_00004;
                    sign_qin_00036_00004  <=  0;
                end else begin
                    conv_qin_00036_00004  <=  ~tout_00036_00004 + 1;
                    sign_qin_00036_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00037 == conv_Sgntin_row_00037_00000 ) begin
                    conv_qin_00037_00000  <= tout_00037_00000;
                    sign_qin_00037_00000  <=  0;
                end else begin
                    conv_qin_00037_00000  <=  ~tout_00037_00000 + 1;
                    sign_qin_00037_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00037 == conv_Sgntin_row_00037_00001 ) begin
                    conv_qin_00037_00001  <= tout_00037_00001;
                    sign_qin_00037_00001  <=  0;
                end else begin
                    conv_qin_00037_00001  <=  ~tout_00037_00001 + 1;
                    sign_qin_00037_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00037 == conv_Sgntin_row_00037_00002 ) begin
                    conv_qin_00037_00002  <= tout_00037_00002;
                    sign_qin_00037_00002  <=  0;
                end else begin
                    conv_qin_00037_00002  <=  ~tout_00037_00002 + 1;
                    sign_qin_00037_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00037 == conv_Sgntin_row_00037_00003 ) begin
                    conv_qin_00037_00003  <= tout_00037_00003;
                    sign_qin_00037_00003  <=  0;
                end else begin
                    conv_qin_00037_00003  <=  ~tout_00037_00003 + 1;
                    sign_qin_00037_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00037 == conv_Sgntin_row_00037_00004 ) begin
                    conv_qin_00037_00004  <= tout_00037_00004;
                    sign_qin_00037_00004  <=  0;
                end else begin
                    conv_qin_00037_00004  <=  ~tout_00037_00004 + 1;
                    sign_qin_00037_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00038 == conv_Sgntin_row_00038_00000 ) begin
                    conv_qin_00038_00000  <= tout_00038_00000;
                    sign_qin_00038_00000  <=  0;
                end else begin
                    conv_qin_00038_00000  <=  ~tout_00038_00000 + 1;
                    sign_qin_00038_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00038 == conv_Sgntin_row_00038_00001 ) begin
                    conv_qin_00038_00001  <= tout_00038_00001;
                    sign_qin_00038_00001  <=  0;
                end else begin
                    conv_qin_00038_00001  <=  ~tout_00038_00001 + 1;
                    sign_qin_00038_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00038 == conv_Sgntin_row_00038_00002 ) begin
                    conv_qin_00038_00002  <= tout_00038_00002;
                    sign_qin_00038_00002  <=  0;
                end else begin
                    conv_qin_00038_00002  <=  ~tout_00038_00002 + 1;
                    sign_qin_00038_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00038 == conv_Sgntin_row_00038_00003 ) begin
                    conv_qin_00038_00003  <= tout_00038_00003;
                    sign_qin_00038_00003  <=  0;
                end else begin
                    conv_qin_00038_00003  <=  ~tout_00038_00003 + 1;
                    sign_qin_00038_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00038 == conv_Sgntin_row_00038_00004 ) begin
                    conv_qin_00038_00004  <= tout_00038_00004;
                    sign_qin_00038_00004  <=  0;
                end else begin
                    conv_qin_00038_00004  <=  ~tout_00038_00004 + 1;
                    sign_qin_00038_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00039 == conv_Sgntin_row_00039_00000 ) begin
                    conv_qin_00039_00000  <= tout_00039_00000;
                    sign_qin_00039_00000  <=  0;
                end else begin
                    conv_qin_00039_00000  <=  ~tout_00039_00000 + 1;
                    sign_qin_00039_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00039 == conv_Sgntin_row_00039_00001 ) begin
                    conv_qin_00039_00001  <= tout_00039_00001;
                    sign_qin_00039_00001  <=  0;
                end else begin
                    conv_qin_00039_00001  <=  ~tout_00039_00001 + 1;
                    sign_qin_00039_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00039 == conv_Sgntin_row_00039_00002 ) begin
                    conv_qin_00039_00002  <= tout_00039_00002;
                    sign_qin_00039_00002  <=  0;
                end else begin
                    conv_qin_00039_00002  <=  ~tout_00039_00002 + 1;
                    sign_qin_00039_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00039 == conv_Sgntin_row_00039_00003 ) begin
                    conv_qin_00039_00003  <= tout_00039_00003;
                    sign_qin_00039_00003  <=  0;
                end else begin
                    conv_qin_00039_00003  <=  ~tout_00039_00003 + 1;
                    sign_qin_00039_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00039 == conv_Sgntin_row_00039_00004 ) begin
                    conv_qin_00039_00004  <= tout_00039_00004;
                    sign_qin_00039_00004  <=  0;
                end else begin
                    conv_qin_00039_00004  <=  ~tout_00039_00004 + 1;
                    sign_qin_00039_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00040 == conv_Sgntin_row_00040_00000 ) begin
                    conv_qin_00040_00000  <= tout_00040_00000;
                    sign_qin_00040_00000  <=  0;
                end else begin
                    conv_qin_00040_00000  <=  ~tout_00040_00000 + 1;
                    sign_qin_00040_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00040 == conv_Sgntin_row_00040_00001 ) begin
                    conv_qin_00040_00001  <= tout_00040_00001;
                    sign_qin_00040_00001  <=  0;
                end else begin
                    conv_qin_00040_00001  <=  ~tout_00040_00001 + 1;
                    sign_qin_00040_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00040 == conv_Sgntin_row_00040_00002 ) begin
                    conv_qin_00040_00002  <= tout_00040_00002;
                    sign_qin_00040_00002  <=  0;
                end else begin
                    conv_qin_00040_00002  <=  ~tout_00040_00002 + 1;
                    sign_qin_00040_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00040 == conv_Sgntin_row_00040_00003 ) begin
                    conv_qin_00040_00003  <= tout_00040_00003;
                    sign_qin_00040_00003  <=  0;
                end else begin
                    conv_qin_00040_00003  <=  ~tout_00040_00003 + 1;
                    sign_qin_00040_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00040 == conv_Sgntin_row_00040_00004 ) begin
                    conv_qin_00040_00004  <= tout_00040_00004;
                    sign_qin_00040_00004  <=  0;
                end else begin
                    conv_qin_00040_00004  <=  ~tout_00040_00004 + 1;
                    sign_qin_00040_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00041 == conv_Sgntin_row_00041_00000 ) begin
                    conv_qin_00041_00000  <= tout_00041_00000;
                    sign_qin_00041_00000  <=  0;
                end else begin
                    conv_qin_00041_00000  <=  ~tout_00041_00000 + 1;
                    sign_qin_00041_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00041 == conv_Sgntin_row_00041_00001 ) begin
                    conv_qin_00041_00001  <= tout_00041_00001;
                    sign_qin_00041_00001  <=  0;
                end else begin
                    conv_qin_00041_00001  <=  ~tout_00041_00001 + 1;
                    sign_qin_00041_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00041 == conv_Sgntin_row_00041_00002 ) begin
                    conv_qin_00041_00002  <= tout_00041_00002;
                    sign_qin_00041_00002  <=  0;
                end else begin
                    conv_qin_00041_00002  <=  ~tout_00041_00002 + 1;
                    sign_qin_00041_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00041 == conv_Sgntin_row_00041_00003 ) begin
                    conv_qin_00041_00003  <= tout_00041_00003;
                    sign_qin_00041_00003  <=  0;
                end else begin
                    conv_qin_00041_00003  <=  ~tout_00041_00003 + 1;
                    sign_qin_00041_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00041 == conv_Sgntin_row_00041_00004 ) begin
                    conv_qin_00041_00004  <= tout_00041_00004;
                    sign_qin_00041_00004  <=  0;
                end else begin
                    conv_qin_00041_00004  <=  ~tout_00041_00004 + 1;
                    sign_qin_00041_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00042 == conv_Sgntin_row_00042_00000 ) begin
                    conv_qin_00042_00000  <= tout_00042_00000;
                    sign_qin_00042_00000  <=  0;
                end else begin
                    conv_qin_00042_00000  <=  ~tout_00042_00000 + 1;
                    sign_qin_00042_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00042 == conv_Sgntin_row_00042_00001 ) begin
                    conv_qin_00042_00001  <= tout_00042_00001;
                    sign_qin_00042_00001  <=  0;
                end else begin
                    conv_qin_00042_00001  <=  ~tout_00042_00001 + 1;
                    sign_qin_00042_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00042 == conv_Sgntin_row_00042_00002 ) begin
                    conv_qin_00042_00002  <= tout_00042_00002;
                    sign_qin_00042_00002  <=  0;
                end else begin
                    conv_qin_00042_00002  <=  ~tout_00042_00002 + 1;
                    sign_qin_00042_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00042 == conv_Sgntin_row_00042_00003 ) begin
                    conv_qin_00042_00003  <= tout_00042_00003;
                    sign_qin_00042_00003  <=  0;
                end else begin
                    conv_qin_00042_00003  <=  ~tout_00042_00003 + 1;
                    sign_qin_00042_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00042 == conv_Sgntin_row_00042_00004 ) begin
                    conv_qin_00042_00004  <= tout_00042_00004;
                    sign_qin_00042_00004  <=  0;
                end else begin
                    conv_qin_00042_00004  <=  ~tout_00042_00004 + 1;
                    sign_qin_00042_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00043 == conv_Sgntin_row_00043_00000 ) begin
                    conv_qin_00043_00000  <= tout_00043_00000;
                    sign_qin_00043_00000  <=  0;
                end else begin
                    conv_qin_00043_00000  <=  ~tout_00043_00000 + 1;
                    sign_qin_00043_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00043 == conv_Sgntin_row_00043_00001 ) begin
                    conv_qin_00043_00001  <= tout_00043_00001;
                    sign_qin_00043_00001  <=  0;
                end else begin
                    conv_qin_00043_00001  <=  ~tout_00043_00001 + 1;
                    sign_qin_00043_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00043 == conv_Sgntin_row_00043_00002 ) begin
                    conv_qin_00043_00002  <= tout_00043_00002;
                    sign_qin_00043_00002  <=  0;
                end else begin
                    conv_qin_00043_00002  <=  ~tout_00043_00002 + 1;
                    sign_qin_00043_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00043 == conv_Sgntin_row_00043_00003 ) begin
                    conv_qin_00043_00003  <= tout_00043_00003;
                    sign_qin_00043_00003  <=  0;
                end else begin
                    conv_qin_00043_00003  <=  ~tout_00043_00003 + 1;
                    sign_qin_00043_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00043 == conv_Sgntin_row_00043_00004 ) begin
                    conv_qin_00043_00004  <= tout_00043_00004;
                    sign_qin_00043_00004  <=  0;
                end else begin
                    conv_qin_00043_00004  <=  ~tout_00043_00004 + 1;
                    sign_qin_00043_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00044 == conv_Sgntin_row_00044_00000 ) begin
                    conv_qin_00044_00000  <= tout_00044_00000;
                    sign_qin_00044_00000  <=  0;
                end else begin
                    conv_qin_00044_00000  <=  ~tout_00044_00000 + 1;
                    sign_qin_00044_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00044 == conv_Sgntin_row_00044_00001 ) begin
                    conv_qin_00044_00001  <= tout_00044_00001;
                    sign_qin_00044_00001  <=  0;
                end else begin
                    conv_qin_00044_00001  <=  ~tout_00044_00001 + 1;
                    sign_qin_00044_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00044 == conv_Sgntin_row_00044_00002 ) begin
                    conv_qin_00044_00002  <= tout_00044_00002;
                    sign_qin_00044_00002  <=  0;
                end else begin
                    conv_qin_00044_00002  <=  ~tout_00044_00002 + 1;
                    sign_qin_00044_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00044 == conv_Sgntin_row_00044_00003 ) begin
                    conv_qin_00044_00003  <= tout_00044_00003;
                    sign_qin_00044_00003  <=  0;
                end else begin
                    conv_qin_00044_00003  <=  ~tout_00044_00003 + 1;
                    sign_qin_00044_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00044 == conv_Sgntin_row_00044_00004 ) begin
                    conv_qin_00044_00004  <= tout_00044_00004;
                    sign_qin_00044_00004  <=  0;
                end else begin
                    conv_qin_00044_00004  <=  ~tout_00044_00004 + 1;
                    sign_qin_00044_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00045 == conv_Sgntin_row_00045_00000 ) begin
                    conv_qin_00045_00000  <= tout_00045_00000;
                    sign_qin_00045_00000  <=  0;
                end else begin
                    conv_qin_00045_00000  <=  ~tout_00045_00000 + 1;
                    sign_qin_00045_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00045 == conv_Sgntin_row_00045_00001 ) begin
                    conv_qin_00045_00001  <= tout_00045_00001;
                    sign_qin_00045_00001  <=  0;
                end else begin
                    conv_qin_00045_00001  <=  ~tout_00045_00001 + 1;
                    sign_qin_00045_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00045 == conv_Sgntin_row_00045_00002 ) begin
                    conv_qin_00045_00002  <= tout_00045_00002;
                    sign_qin_00045_00002  <=  0;
                end else begin
                    conv_qin_00045_00002  <=  ~tout_00045_00002 + 1;
                    sign_qin_00045_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00045 == conv_Sgntin_row_00045_00003 ) begin
                    conv_qin_00045_00003  <= tout_00045_00003;
                    sign_qin_00045_00003  <=  0;
                end else begin
                    conv_qin_00045_00003  <=  ~tout_00045_00003 + 1;
                    sign_qin_00045_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00045 == conv_Sgntin_row_00045_00004 ) begin
                    conv_qin_00045_00004  <= tout_00045_00004;
                    sign_qin_00045_00004  <=  0;
                end else begin
                    conv_qin_00045_00004  <=  ~tout_00045_00004 + 1;
                    sign_qin_00045_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00046 == conv_Sgntin_row_00046_00000 ) begin
                    conv_qin_00046_00000  <= tout_00046_00000;
                    sign_qin_00046_00000  <=  0;
                end else begin
                    conv_qin_00046_00000  <=  ~tout_00046_00000 + 1;
                    sign_qin_00046_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00046 == conv_Sgntin_row_00046_00001 ) begin
                    conv_qin_00046_00001  <= tout_00046_00001;
                    sign_qin_00046_00001  <=  0;
                end else begin
                    conv_qin_00046_00001  <=  ~tout_00046_00001 + 1;
                    sign_qin_00046_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00046 == conv_Sgntin_row_00046_00002 ) begin
                    conv_qin_00046_00002  <= tout_00046_00002;
                    sign_qin_00046_00002  <=  0;
                end else begin
                    conv_qin_00046_00002  <=  ~tout_00046_00002 + 1;
                    sign_qin_00046_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00046 == conv_Sgntin_row_00046_00003 ) begin
                    conv_qin_00046_00003  <= tout_00046_00003;
                    sign_qin_00046_00003  <=  0;
                end else begin
                    conv_qin_00046_00003  <=  ~tout_00046_00003 + 1;
                    sign_qin_00046_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00046 == conv_Sgntin_row_00046_00004 ) begin
                    conv_qin_00046_00004  <= tout_00046_00004;
                    sign_qin_00046_00004  <=  0;
                end else begin
                    conv_qin_00046_00004  <=  ~tout_00046_00004 + 1;
                    sign_qin_00046_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00047 == conv_Sgntin_row_00047_00000 ) begin
                    conv_qin_00047_00000  <= tout_00047_00000;
                    sign_qin_00047_00000  <=  0;
                end else begin
                    conv_qin_00047_00000  <=  ~tout_00047_00000 + 1;
                    sign_qin_00047_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00047 == conv_Sgntin_row_00047_00001 ) begin
                    conv_qin_00047_00001  <= tout_00047_00001;
                    sign_qin_00047_00001  <=  0;
                end else begin
                    conv_qin_00047_00001  <=  ~tout_00047_00001 + 1;
                    sign_qin_00047_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00047 == conv_Sgntin_row_00047_00002 ) begin
                    conv_qin_00047_00002  <= tout_00047_00002;
                    sign_qin_00047_00002  <=  0;
                end else begin
                    conv_qin_00047_00002  <=  ~tout_00047_00002 + 1;
                    sign_qin_00047_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00047 == conv_Sgntin_row_00047_00003 ) begin
                    conv_qin_00047_00003  <= tout_00047_00003;
                    sign_qin_00047_00003  <=  0;
                end else begin
                    conv_qin_00047_00003  <=  ~tout_00047_00003 + 1;
                    sign_qin_00047_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00047 == conv_Sgntin_row_00047_00004 ) begin
                    conv_qin_00047_00004  <= tout_00047_00004;
                    sign_qin_00047_00004  <=  0;
                end else begin
                    conv_qin_00047_00004  <=  ~tout_00047_00004 + 1;
                    sign_qin_00047_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00048 == conv_Sgntin_row_00048_00000 ) begin
                    conv_qin_00048_00000  <= tout_00048_00000;
                    sign_qin_00048_00000  <=  0;
                end else begin
                    conv_qin_00048_00000  <=  ~tout_00048_00000 + 1;
                    sign_qin_00048_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00048 == conv_Sgntin_row_00048_00001 ) begin
                    conv_qin_00048_00001  <= tout_00048_00001;
                    sign_qin_00048_00001  <=  0;
                end else begin
                    conv_qin_00048_00001  <=  ~tout_00048_00001 + 1;
                    sign_qin_00048_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00048 == conv_Sgntin_row_00048_00002 ) begin
                    conv_qin_00048_00002  <= tout_00048_00002;
                    sign_qin_00048_00002  <=  0;
                end else begin
                    conv_qin_00048_00002  <=  ~tout_00048_00002 + 1;
                    sign_qin_00048_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00048 == conv_Sgntin_row_00048_00003 ) begin
                    conv_qin_00048_00003  <= tout_00048_00003;
                    sign_qin_00048_00003  <=  0;
                end else begin
                    conv_qin_00048_00003  <=  ~tout_00048_00003 + 1;
                    sign_qin_00048_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00049 == conv_Sgntin_row_00049_00000 ) begin
                    conv_qin_00049_00000  <= tout_00049_00000;
                    sign_qin_00049_00000  <=  0;
                end else begin
                    conv_qin_00049_00000  <=  ~tout_00049_00000 + 1;
                    sign_qin_00049_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00049 == conv_Sgntin_row_00049_00001 ) begin
                    conv_qin_00049_00001  <= tout_00049_00001;
                    sign_qin_00049_00001  <=  0;
                end else begin
                    conv_qin_00049_00001  <=  ~tout_00049_00001 + 1;
                    sign_qin_00049_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00049 == conv_Sgntin_row_00049_00002 ) begin
                    conv_qin_00049_00002  <= tout_00049_00002;
                    sign_qin_00049_00002  <=  0;
                end else begin
                    conv_qin_00049_00002  <=  ~tout_00049_00002 + 1;
                    sign_qin_00049_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00049 == conv_Sgntin_row_00049_00003 ) begin
                    conv_qin_00049_00003  <= tout_00049_00003;
                    sign_qin_00049_00003  <=  0;
                end else begin
                    conv_qin_00049_00003  <=  ~tout_00049_00003 + 1;
                    sign_qin_00049_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00050 == conv_Sgntin_row_00050_00000 ) begin
                    conv_qin_00050_00000  <= tout_00050_00000;
                    sign_qin_00050_00000  <=  0;
                end else begin
                    conv_qin_00050_00000  <=  ~tout_00050_00000 + 1;
                    sign_qin_00050_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00050 == conv_Sgntin_row_00050_00001 ) begin
                    conv_qin_00050_00001  <= tout_00050_00001;
                    sign_qin_00050_00001  <=  0;
                end else begin
                    conv_qin_00050_00001  <=  ~tout_00050_00001 + 1;
                    sign_qin_00050_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00050 == conv_Sgntin_row_00050_00002 ) begin
                    conv_qin_00050_00002  <= tout_00050_00002;
                    sign_qin_00050_00002  <=  0;
                end else begin
                    conv_qin_00050_00002  <=  ~tout_00050_00002 + 1;
                    sign_qin_00050_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00050 == conv_Sgntin_row_00050_00003 ) begin
                    conv_qin_00050_00003  <= tout_00050_00003;
                    sign_qin_00050_00003  <=  0;
                end else begin
                    conv_qin_00050_00003  <=  ~tout_00050_00003 + 1;
                    sign_qin_00050_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00051 == conv_Sgntin_row_00051_00000 ) begin
                    conv_qin_00051_00000  <= tout_00051_00000;
                    sign_qin_00051_00000  <=  0;
                end else begin
                    conv_qin_00051_00000  <=  ~tout_00051_00000 + 1;
                    sign_qin_00051_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00051 == conv_Sgntin_row_00051_00001 ) begin
                    conv_qin_00051_00001  <= tout_00051_00001;
                    sign_qin_00051_00001  <=  0;
                end else begin
                    conv_qin_00051_00001  <=  ~tout_00051_00001 + 1;
                    sign_qin_00051_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00051 == conv_Sgntin_row_00051_00002 ) begin
                    conv_qin_00051_00002  <= tout_00051_00002;
                    sign_qin_00051_00002  <=  0;
                end else begin
                    conv_qin_00051_00002  <=  ~tout_00051_00002 + 1;
                    sign_qin_00051_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00051 == conv_Sgntin_row_00051_00003 ) begin
                    conv_qin_00051_00003  <= tout_00051_00003;
                    sign_qin_00051_00003  <=  0;
                end else begin
                    conv_qin_00051_00003  <=  ~tout_00051_00003 + 1;
                    sign_qin_00051_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00052 == conv_Sgntin_row_00052_00000 ) begin
                    conv_qin_00052_00000  <= tout_00052_00000;
                    sign_qin_00052_00000  <=  0;
                end else begin
                    conv_qin_00052_00000  <=  ~tout_00052_00000 + 1;
                    sign_qin_00052_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00052 == conv_Sgntin_row_00052_00001 ) begin
                    conv_qin_00052_00001  <= tout_00052_00001;
                    sign_qin_00052_00001  <=  0;
                end else begin
                    conv_qin_00052_00001  <=  ~tout_00052_00001 + 1;
                    sign_qin_00052_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00052 == conv_Sgntin_row_00052_00002 ) begin
                    conv_qin_00052_00002  <= tout_00052_00002;
                    sign_qin_00052_00002  <=  0;
                end else begin
                    conv_qin_00052_00002  <=  ~tout_00052_00002 + 1;
                    sign_qin_00052_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00052 == conv_Sgntin_row_00052_00003 ) begin
                    conv_qin_00052_00003  <= tout_00052_00003;
                    sign_qin_00052_00003  <=  0;
                end else begin
                    conv_qin_00052_00003  <=  ~tout_00052_00003 + 1;
                    sign_qin_00052_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00052 == conv_Sgntin_row_00052_00004 ) begin
                    conv_qin_00052_00004  <= tout_00052_00004;
                    sign_qin_00052_00004  <=  0;
                end else begin
                    conv_qin_00052_00004  <=  ~tout_00052_00004 + 1;
                    sign_qin_00052_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00053 == conv_Sgntin_row_00053_00000 ) begin
                    conv_qin_00053_00000  <= tout_00053_00000;
                    sign_qin_00053_00000  <=  0;
                end else begin
                    conv_qin_00053_00000  <=  ~tout_00053_00000 + 1;
                    sign_qin_00053_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00053 == conv_Sgntin_row_00053_00001 ) begin
                    conv_qin_00053_00001  <= tout_00053_00001;
                    sign_qin_00053_00001  <=  0;
                end else begin
                    conv_qin_00053_00001  <=  ~tout_00053_00001 + 1;
                    sign_qin_00053_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00053 == conv_Sgntin_row_00053_00002 ) begin
                    conv_qin_00053_00002  <= tout_00053_00002;
                    sign_qin_00053_00002  <=  0;
                end else begin
                    conv_qin_00053_00002  <=  ~tout_00053_00002 + 1;
                    sign_qin_00053_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00053 == conv_Sgntin_row_00053_00003 ) begin
                    conv_qin_00053_00003  <= tout_00053_00003;
                    sign_qin_00053_00003  <=  0;
                end else begin
                    conv_qin_00053_00003  <=  ~tout_00053_00003 + 1;
                    sign_qin_00053_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00053 == conv_Sgntin_row_00053_00004 ) begin
                    conv_qin_00053_00004  <= tout_00053_00004;
                    sign_qin_00053_00004  <=  0;
                end else begin
                    conv_qin_00053_00004  <=  ~tout_00053_00004 + 1;
                    sign_qin_00053_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00054 == conv_Sgntin_row_00054_00000 ) begin
                    conv_qin_00054_00000  <= tout_00054_00000;
                    sign_qin_00054_00000  <=  0;
                end else begin
                    conv_qin_00054_00000  <=  ~tout_00054_00000 + 1;
                    sign_qin_00054_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00054 == conv_Sgntin_row_00054_00001 ) begin
                    conv_qin_00054_00001  <= tout_00054_00001;
                    sign_qin_00054_00001  <=  0;
                end else begin
                    conv_qin_00054_00001  <=  ~tout_00054_00001 + 1;
                    sign_qin_00054_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00054 == conv_Sgntin_row_00054_00002 ) begin
                    conv_qin_00054_00002  <= tout_00054_00002;
                    sign_qin_00054_00002  <=  0;
                end else begin
                    conv_qin_00054_00002  <=  ~tout_00054_00002 + 1;
                    sign_qin_00054_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00054 == conv_Sgntin_row_00054_00003 ) begin
                    conv_qin_00054_00003  <= tout_00054_00003;
                    sign_qin_00054_00003  <=  0;
                end else begin
                    conv_qin_00054_00003  <=  ~tout_00054_00003 + 1;
                    sign_qin_00054_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00054 == conv_Sgntin_row_00054_00004 ) begin
                    conv_qin_00054_00004  <= tout_00054_00004;
                    sign_qin_00054_00004  <=  0;
                end else begin
                    conv_qin_00054_00004  <=  ~tout_00054_00004 + 1;
                    sign_qin_00054_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00055 == conv_Sgntin_row_00055_00000 ) begin
                    conv_qin_00055_00000  <= tout_00055_00000;
                    sign_qin_00055_00000  <=  0;
                end else begin
                    conv_qin_00055_00000  <=  ~tout_00055_00000 + 1;
                    sign_qin_00055_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00055 == conv_Sgntin_row_00055_00001 ) begin
                    conv_qin_00055_00001  <= tout_00055_00001;
                    sign_qin_00055_00001  <=  0;
                end else begin
                    conv_qin_00055_00001  <=  ~tout_00055_00001 + 1;
                    sign_qin_00055_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00055 == conv_Sgntin_row_00055_00002 ) begin
                    conv_qin_00055_00002  <= tout_00055_00002;
                    sign_qin_00055_00002  <=  0;
                end else begin
                    conv_qin_00055_00002  <=  ~tout_00055_00002 + 1;
                    sign_qin_00055_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00055 == conv_Sgntin_row_00055_00003 ) begin
                    conv_qin_00055_00003  <= tout_00055_00003;
                    sign_qin_00055_00003  <=  0;
                end else begin
                    conv_qin_00055_00003  <=  ~tout_00055_00003 + 1;
                    sign_qin_00055_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00055 == conv_Sgntin_row_00055_00004 ) begin
                    conv_qin_00055_00004  <= tout_00055_00004;
                    sign_qin_00055_00004  <=  0;
                end else begin
                    conv_qin_00055_00004  <=  ~tout_00055_00004 + 1;
                    sign_qin_00055_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00056 == conv_Sgntin_row_00056_00000 ) begin
                    conv_qin_00056_00000  <= tout_00056_00000;
                    sign_qin_00056_00000  <=  0;
                end else begin
                    conv_qin_00056_00000  <=  ~tout_00056_00000 + 1;
                    sign_qin_00056_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00056 == conv_Sgntin_row_00056_00001 ) begin
                    conv_qin_00056_00001  <= tout_00056_00001;
                    sign_qin_00056_00001  <=  0;
                end else begin
                    conv_qin_00056_00001  <=  ~tout_00056_00001 + 1;
                    sign_qin_00056_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00056 == conv_Sgntin_row_00056_00002 ) begin
                    conv_qin_00056_00002  <= tout_00056_00002;
                    sign_qin_00056_00002  <=  0;
                end else begin
                    conv_qin_00056_00002  <=  ~tout_00056_00002 + 1;
                    sign_qin_00056_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00056 == conv_Sgntin_row_00056_00003 ) begin
                    conv_qin_00056_00003  <= tout_00056_00003;
                    sign_qin_00056_00003  <=  0;
                end else begin
                    conv_qin_00056_00003  <=  ~tout_00056_00003 + 1;
                    sign_qin_00056_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00056 == conv_Sgntin_row_00056_00004 ) begin
                    conv_qin_00056_00004  <= tout_00056_00004;
                    sign_qin_00056_00004  <=  0;
                end else begin
                    conv_qin_00056_00004  <=  ~tout_00056_00004 + 1;
                    sign_qin_00056_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00057 == conv_Sgntin_row_00057_00000 ) begin
                    conv_qin_00057_00000  <= tout_00057_00000;
                    sign_qin_00057_00000  <=  0;
                end else begin
                    conv_qin_00057_00000  <=  ~tout_00057_00000 + 1;
                    sign_qin_00057_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00057 == conv_Sgntin_row_00057_00001 ) begin
                    conv_qin_00057_00001  <= tout_00057_00001;
                    sign_qin_00057_00001  <=  0;
                end else begin
                    conv_qin_00057_00001  <=  ~tout_00057_00001 + 1;
                    sign_qin_00057_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00057 == conv_Sgntin_row_00057_00002 ) begin
                    conv_qin_00057_00002  <= tout_00057_00002;
                    sign_qin_00057_00002  <=  0;
                end else begin
                    conv_qin_00057_00002  <=  ~tout_00057_00002 + 1;
                    sign_qin_00057_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00057 == conv_Sgntin_row_00057_00003 ) begin
                    conv_qin_00057_00003  <= tout_00057_00003;
                    sign_qin_00057_00003  <=  0;
                end else begin
                    conv_qin_00057_00003  <=  ~tout_00057_00003 + 1;
                    sign_qin_00057_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00057 == conv_Sgntin_row_00057_00004 ) begin
                    conv_qin_00057_00004  <= tout_00057_00004;
                    sign_qin_00057_00004  <=  0;
                end else begin
                    conv_qin_00057_00004  <=  ~tout_00057_00004 + 1;
                    sign_qin_00057_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00058 == conv_Sgntin_row_00058_00000 ) begin
                    conv_qin_00058_00000  <= tout_00058_00000;
                    sign_qin_00058_00000  <=  0;
                end else begin
                    conv_qin_00058_00000  <=  ~tout_00058_00000 + 1;
                    sign_qin_00058_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00058 == conv_Sgntin_row_00058_00001 ) begin
                    conv_qin_00058_00001  <= tout_00058_00001;
                    sign_qin_00058_00001  <=  0;
                end else begin
                    conv_qin_00058_00001  <=  ~tout_00058_00001 + 1;
                    sign_qin_00058_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00058 == conv_Sgntin_row_00058_00002 ) begin
                    conv_qin_00058_00002  <= tout_00058_00002;
                    sign_qin_00058_00002  <=  0;
                end else begin
                    conv_qin_00058_00002  <=  ~tout_00058_00002 + 1;
                    sign_qin_00058_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00058 == conv_Sgntin_row_00058_00003 ) begin
                    conv_qin_00058_00003  <= tout_00058_00003;
                    sign_qin_00058_00003  <=  0;
                end else begin
                    conv_qin_00058_00003  <=  ~tout_00058_00003 + 1;
                    sign_qin_00058_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00058 == conv_Sgntin_row_00058_00004 ) begin
                    conv_qin_00058_00004  <= tout_00058_00004;
                    sign_qin_00058_00004  <=  0;
                end else begin
                    conv_qin_00058_00004  <=  ~tout_00058_00004 + 1;
                    sign_qin_00058_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00059 == conv_Sgntin_row_00059_00000 ) begin
                    conv_qin_00059_00000  <= tout_00059_00000;
                    sign_qin_00059_00000  <=  0;
                end else begin
                    conv_qin_00059_00000  <=  ~tout_00059_00000 + 1;
                    sign_qin_00059_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00059 == conv_Sgntin_row_00059_00001 ) begin
                    conv_qin_00059_00001  <= tout_00059_00001;
                    sign_qin_00059_00001  <=  0;
                end else begin
                    conv_qin_00059_00001  <=  ~tout_00059_00001 + 1;
                    sign_qin_00059_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00059 == conv_Sgntin_row_00059_00002 ) begin
                    conv_qin_00059_00002  <= tout_00059_00002;
                    sign_qin_00059_00002  <=  0;
                end else begin
                    conv_qin_00059_00002  <=  ~tout_00059_00002 + 1;
                    sign_qin_00059_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00059 == conv_Sgntin_row_00059_00003 ) begin
                    conv_qin_00059_00003  <= tout_00059_00003;
                    sign_qin_00059_00003  <=  0;
                end else begin
                    conv_qin_00059_00003  <=  ~tout_00059_00003 + 1;
                    sign_qin_00059_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00059 == conv_Sgntin_row_00059_00004 ) begin
                    conv_qin_00059_00004  <= tout_00059_00004;
                    sign_qin_00059_00004  <=  0;
                end else begin
                    conv_qin_00059_00004  <=  ~tout_00059_00004 + 1;
                    sign_qin_00059_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00060 == conv_Sgntin_row_00060_00000 ) begin
                    conv_qin_00060_00000  <= tout_00060_00000;
                    sign_qin_00060_00000  <=  0;
                end else begin
                    conv_qin_00060_00000  <=  ~tout_00060_00000 + 1;
                    sign_qin_00060_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00060 == conv_Sgntin_row_00060_00001 ) begin
                    conv_qin_00060_00001  <= tout_00060_00001;
                    sign_qin_00060_00001  <=  0;
                end else begin
                    conv_qin_00060_00001  <=  ~tout_00060_00001 + 1;
                    sign_qin_00060_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00060 == conv_Sgntin_row_00060_00002 ) begin
                    conv_qin_00060_00002  <= tout_00060_00002;
                    sign_qin_00060_00002  <=  0;
                end else begin
                    conv_qin_00060_00002  <=  ~tout_00060_00002 + 1;
                    sign_qin_00060_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00060 == conv_Sgntin_row_00060_00003 ) begin
                    conv_qin_00060_00003  <= tout_00060_00003;
                    sign_qin_00060_00003  <=  0;
                end else begin
                    conv_qin_00060_00003  <=  ~tout_00060_00003 + 1;
                    sign_qin_00060_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00061 == conv_Sgntin_row_00061_00000 ) begin
                    conv_qin_00061_00000  <= tout_00061_00000;
                    sign_qin_00061_00000  <=  0;
                end else begin
                    conv_qin_00061_00000  <=  ~tout_00061_00000 + 1;
                    sign_qin_00061_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00061 == conv_Sgntin_row_00061_00001 ) begin
                    conv_qin_00061_00001  <= tout_00061_00001;
                    sign_qin_00061_00001  <=  0;
                end else begin
                    conv_qin_00061_00001  <=  ~tout_00061_00001 + 1;
                    sign_qin_00061_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00061 == conv_Sgntin_row_00061_00002 ) begin
                    conv_qin_00061_00002  <= tout_00061_00002;
                    sign_qin_00061_00002  <=  0;
                end else begin
                    conv_qin_00061_00002  <=  ~tout_00061_00002 + 1;
                    sign_qin_00061_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00061 == conv_Sgntin_row_00061_00003 ) begin
                    conv_qin_00061_00003  <= tout_00061_00003;
                    sign_qin_00061_00003  <=  0;
                end else begin
                    conv_qin_00061_00003  <=  ~tout_00061_00003 + 1;
                    sign_qin_00061_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00062 == conv_Sgntin_row_00062_00000 ) begin
                    conv_qin_00062_00000  <= tout_00062_00000;
                    sign_qin_00062_00000  <=  0;
                end else begin
                    conv_qin_00062_00000  <=  ~tout_00062_00000 + 1;
                    sign_qin_00062_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00062 == conv_Sgntin_row_00062_00001 ) begin
                    conv_qin_00062_00001  <= tout_00062_00001;
                    sign_qin_00062_00001  <=  0;
                end else begin
                    conv_qin_00062_00001  <=  ~tout_00062_00001 + 1;
                    sign_qin_00062_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00062 == conv_Sgntin_row_00062_00002 ) begin
                    conv_qin_00062_00002  <= tout_00062_00002;
                    sign_qin_00062_00002  <=  0;
                end else begin
                    conv_qin_00062_00002  <=  ~tout_00062_00002 + 1;
                    sign_qin_00062_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00062 == conv_Sgntin_row_00062_00003 ) begin
                    conv_qin_00062_00003  <= tout_00062_00003;
                    sign_qin_00062_00003  <=  0;
                end else begin
                    conv_qin_00062_00003  <=  ~tout_00062_00003 + 1;
                    sign_qin_00062_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00063 == conv_Sgntin_row_00063_00000 ) begin
                    conv_qin_00063_00000  <= tout_00063_00000;
                    sign_qin_00063_00000  <=  0;
                end else begin
                    conv_qin_00063_00000  <=  ~tout_00063_00000 + 1;
                    sign_qin_00063_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00063 == conv_Sgntin_row_00063_00001 ) begin
                    conv_qin_00063_00001  <= tout_00063_00001;
                    sign_qin_00063_00001  <=  0;
                end else begin
                    conv_qin_00063_00001  <=  ~tout_00063_00001 + 1;
                    sign_qin_00063_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00063 == conv_Sgntin_row_00063_00002 ) begin
                    conv_qin_00063_00002  <= tout_00063_00002;
                    sign_qin_00063_00002  <=  0;
                end else begin
                    conv_qin_00063_00002  <=  ~tout_00063_00002 + 1;
                    sign_qin_00063_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00063 == conv_Sgntin_row_00063_00003 ) begin
                    conv_qin_00063_00003  <= tout_00063_00003;
                    sign_qin_00063_00003  <=  0;
                end else begin
                    conv_qin_00063_00003  <=  ~tout_00063_00003 + 1;
                    sign_qin_00063_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00064 == conv_Sgntin_row_00064_00000 ) begin
                    conv_qin_00064_00000  <= tout_00064_00000;
                    sign_qin_00064_00000  <=  0;
                end else begin
                    conv_qin_00064_00000  <=  ~tout_00064_00000 + 1;
                    sign_qin_00064_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00064 == conv_Sgntin_row_00064_00001 ) begin
                    conv_qin_00064_00001  <= tout_00064_00001;
                    sign_qin_00064_00001  <=  0;
                end else begin
                    conv_qin_00064_00001  <=  ~tout_00064_00001 + 1;
                    sign_qin_00064_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00064 == conv_Sgntin_row_00064_00002 ) begin
                    conv_qin_00064_00002  <= tout_00064_00002;
                    sign_qin_00064_00002  <=  0;
                end else begin
                    conv_qin_00064_00002  <=  ~tout_00064_00002 + 1;
                    sign_qin_00064_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00064 == conv_Sgntin_row_00064_00003 ) begin
                    conv_qin_00064_00003  <= tout_00064_00003;
                    sign_qin_00064_00003  <=  0;
                end else begin
                    conv_qin_00064_00003  <=  ~tout_00064_00003 + 1;
                    sign_qin_00064_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00064 == conv_Sgntin_row_00064_00004 ) begin
                    conv_qin_00064_00004  <= tout_00064_00004;
                    sign_qin_00064_00004  <=  0;
                end else begin
                    conv_qin_00064_00004  <=  ~tout_00064_00004 + 1;
                    sign_qin_00064_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00065 == conv_Sgntin_row_00065_00000 ) begin
                    conv_qin_00065_00000  <= tout_00065_00000;
                    sign_qin_00065_00000  <=  0;
                end else begin
                    conv_qin_00065_00000  <=  ~tout_00065_00000 + 1;
                    sign_qin_00065_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00065 == conv_Sgntin_row_00065_00001 ) begin
                    conv_qin_00065_00001  <= tout_00065_00001;
                    sign_qin_00065_00001  <=  0;
                end else begin
                    conv_qin_00065_00001  <=  ~tout_00065_00001 + 1;
                    sign_qin_00065_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00065 == conv_Sgntin_row_00065_00002 ) begin
                    conv_qin_00065_00002  <= tout_00065_00002;
                    sign_qin_00065_00002  <=  0;
                end else begin
                    conv_qin_00065_00002  <=  ~tout_00065_00002 + 1;
                    sign_qin_00065_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00065 == conv_Sgntin_row_00065_00003 ) begin
                    conv_qin_00065_00003  <= tout_00065_00003;
                    sign_qin_00065_00003  <=  0;
                end else begin
                    conv_qin_00065_00003  <=  ~tout_00065_00003 + 1;
                    sign_qin_00065_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00065 == conv_Sgntin_row_00065_00004 ) begin
                    conv_qin_00065_00004  <= tout_00065_00004;
                    sign_qin_00065_00004  <=  0;
                end else begin
                    conv_qin_00065_00004  <=  ~tout_00065_00004 + 1;
                    sign_qin_00065_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00066 == conv_Sgntin_row_00066_00000 ) begin
                    conv_qin_00066_00000  <= tout_00066_00000;
                    sign_qin_00066_00000  <=  0;
                end else begin
                    conv_qin_00066_00000  <=  ~tout_00066_00000 + 1;
                    sign_qin_00066_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00066 == conv_Sgntin_row_00066_00001 ) begin
                    conv_qin_00066_00001  <= tout_00066_00001;
                    sign_qin_00066_00001  <=  0;
                end else begin
                    conv_qin_00066_00001  <=  ~tout_00066_00001 + 1;
                    sign_qin_00066_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00066 == conv_Sgntin_row_00066_00002 ) begin
                    conv_qin_00066_00002  <= tout_00066_00002;
                    sign_qin_00066_00002  <=  0;
                end else begin
                    conv_qin_00066_00002  <=  ~tout_00066_00002 + 1;
                    sign_qin_00066_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00066 == conv_Sgntin_row_00066_00003 ) begin
                    conv_qin_00066_00003  <= tout_00066_00003;
                    sign_qin_00066_00003  <=  0;
                end else begin
                    conv_qin_00066_00003  <=  ~tout_00066_00003 + 1;
                    sign_qin_00066_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00066 == conv_Sgntin_row_00066_00004 ) begin
                    conv_qin_00066_00004  <= tout_00066_00004;
                    sign_qin_00066_00004  <=  0;
                end else begin
                    conv_qin_00066_00004  <=  ~tout_00066_00004 + 1;
                    sign_qin_00066_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00067 == conv_Sgntin_row_00067_00000 ) begin
                    conv_qin_00067_00000  <= tout_00067_00000;
                    sign_qin_00067_00000  <=  0;
                end else begin
                    conv_qin_00067_00000  <=  ~tout_00067_00000 + 1;
                    sign_qin_00067_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00067 == conv_Sgntin_row_00067_00001 ) begin
                    conv_qin_00067_00001  <= tout_00067_00001;
                    sign_qin_00067_00001  <=  0;
                end else begin
                    conv_qin_00067_00001  <=  ~tout_00067_00001 + 1;
                    sign_qin_00067_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00067 == conv_Sgntin_row_00067_00002 ) begin
                    conv_qin_00067_00002  <= tout_00067_00002;
                    sign_qin_00067_00002  <=  0;
                end else begin
                    conv_qin_00067_00002  <=  ~tout_00067_00002 + 1;
                    sign_qin_00067_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00067 == conv_Sgntin_row_00067_00003 ) begin
                    conv_qin_00067_00003  <= tout_00067_00003;
                    sign_qin_00067_00003  <=  0;
                end else begin
                    conv_qin_00067_00003  <=  ~tout_00067_00003 + 1;
                    sign_qin_00067_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00067 == conv_Sgntin_row_00067_00004 ) begin
                    conv_qin_00067_00004  <= tout_00067_00004;
                    sign_qin_00067_00004  <=  0;
                end else begin
                    conv_qin_00067_00004  <=  ~tout_00067_00004 + 1;
                    sign_qin_00067_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00068 == conv_Sgntin_row_00068_00000 ) begin
                    conv_qin_00068_00000  <= tout_00068_00000;
                    sign_qin_00068_00000  <=  0;
                end else begin
                    conv_qin_00068_00000  <=  ~tout_00068_00000 + 1;
                    sign_qin_00068_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00068 == conv_Sgntin_row_00068_00001 ) begin
                    conv_qin_00068_00001  <= tout_00068_00001;
                    sign_qin_00068_00001  <=  0;
                end else begin
                    conv_qin_00068_00001  <=  ~tout_00068_00001 + 1;
                    sign_qin_00068_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00068 == conv_Sgntin_row_00068_00002 ) begin
                    conv_qin_00068_00002  <= tout_00068_00002;
                    sign_qin_00068_00002  <=  0;
                end else begin
                    conv_qin_00068_00002  <=  ~tout_00068_00002 + 1;
                    sign_qin_00068_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00068 == conv_Sgntin_row_00068_00003 ) begin
                    conv_qin_00068_00003  <= tout_00068_00003;
                    sign_qin_00068_00003  <=  0;
                end else begin
                    conv_qin_00068_00003  <=  ~tout_00068_00003 + 1;
                    sign_qin_00068_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00068 == conv_Sgntin_row_00068_00004 ) begin
                    conv_qin_00068_00004  <= tout_00068_00004;
                    sign_qin_00068_00004  <=  0;
                end else begin
                    conv_qin_00068_00004  <=  ~tout_00068_00004 + 1;
                    sign_qin_00068_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00069 == conv_Sgntin_row_00069_00000 ) begin
                    conv_qin_00069_00000  <= tout_00069_00000;
                    sign_qin_00069_00000  <=  0;
                end else begin
                    conv_qin_00069_00000  <=  ~tout_00069_00000 + 1;
                    sign_qin_00069_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00069 == conv_Sgntin_row_00069_00001 ) begin
                    conv_qin_00069_00001  <= tout_00069_00001;
                    sign_qin_00069_00001  <=  0;
                end else begin
                    conv_qin_00069_00001  <=  ~tout_00069_00001 + 1;
                    sign_qin_00069_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00069 == conv_Sgntin_row_00069_00002 ) begin
                    conv_qin_00069_00002  <= tout_00069_00002;
                    sign_qin_00069_00002  <=  0;
                end else begin
                    conv_qin_00069_00002  <=  ~tout_00069_00002 + 1;
                    sign_qin_00069_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00069 == conv_Sgntin_row_00069_00003 ) begin
                    conv_qin_00069_00003  <= tout_00069_00003;
                    sign_qin_00069_00003  <=  0;
                end else begin
                    conv_qin_00069_00003  <=  ~tout_00069_00003 + 1;
                    sign_qin_00069_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00069 == conv_Sgntin_row_00069_00004 ) begin
                    conv_qin_00069_00004  <= tout_00069_00004;
                    sign_qin_00069_00004  <=  0;
                end else begin
                    conv_qin_00069_00004  <=  ~tout_00069_00004 + 1;
                    sign_qin_00069_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00070 == conv_Sgntin_row_00070_00000 ) begin
                    conv_qin_00070_00000  <= tout_00070_00000;
                    sign_qin_00070_00000  <=  0;
                end else begin
                    conv_qin_00070_00000  <=  ~tout_00070_00000 + 1;
                    sign_qin_00070_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00070 == conv_Sgntin_row_00070_00001 ) begin
                    conv_qin_00070_00001  <= tout_00070_00001;
                    sign_qin_00070_00001  <=  0;
                end else begin
                    conv_qin_00070_00001  <=  ~tout_00070_00001 + 1;
                    sign_qin_00070_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00070 == conv_Sgntin_row_00070_00002 ) begin
                    conv_qin_00070_00002  <= tout_00070_00002;
                    sign_qin_00070_00002  <=  0;
                end else begin
                    conv_qin_00070_00002  <=  ~tout_00070_00002 + 1;
                    sign_qin_00070_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00070 == conv_Sgntin_row_00070_00003 ) begin
                    conv_qin_00070_00003  <= tout_00070_00003;
                    sign_qin_00070_00003  <=  0;
                end else begin
                    conv_qin_00070_00003  <=  ~tout_00070_00003 + 1;
                    sign_qin_00070_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00070 == conv_Sgntin_row_00070_00004 ) begin
                    conv_qin_00070_00004  <= tout_00070_00004;
                    sign_qin_00070_00004  <=  0;
                end else begin
                    conv_qin_00070_00004  <=  ~tout_00070_00004 + 1;
                    sign_qin_00070_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00071 == conv_Sgntin_row_00071_00000 ) begin
                    conv_qin_00071_00000  <= tout_00071_00000;
                    sign_qin_00071_00000  <=  0;
                end else begin
                    conv_qin_00071_00000  <=  ~tout_00071_00000 + 1;
                    sign_qin_00071_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00071 == conv_Sgntin_row_00071_00001 ) begin
                    conv_qin_00071_00001  <= tout_00071_00001;
                    sign_qin_00071_00001  <=  0;
                end else begin
                    conv_qin_00071_00001  <=  ~tout_00071_00001 + 1;
                    sign_qin_00071_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00071 == conv_Sgntin_row_00071_00002 ) begin
                    conv_qin_00071_00002  <= tout_00071_00002;
                    sign_qin_00071_00002  <=  0;
                end else begin
                    conv_qin_00071_00002  <=  ~tout_00071_00002 + 1;
                    sign_qin_00071_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00071 == conv_Sgntin_row_00071_00003 ) begin
                    conv_qin_00071_00003  <= tout_00071_00003;
                    sign_qin_00071_00003  <=  0;
                end else begin
                    conv_qin_00071_00003  <=  ~tout_00071_00003 + 1;
                    sign_qin_00071_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00071 == conv_Sgntin_row_00071_00004 ) begin
                    conv_qin_00071_00004  <= tout_00071_00004;
                    sign_qin_00071_00004  <=  0;
                end else begin
                    conv_qin_00071_00004  <=  ~tout_00071_00004 + 1;
                    sign_qin_00071_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00072 == conv_Sgntin_row_00072_00000 ) begin
                    conv_qin_00072_00000  <= tout_00072_00000;
                    sign_qin_00072_00000  <=  0;
                end else begin
                    conv_qin_00072_00000  <=  ~tout_00072_00000 + 1;
                    sign_qin_00072_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00072 == conv_Sgntin_row_00072_00001 ) begin
                    conv_qin_00072_00001  <= tout_00072_00001;
                    sign_qin_00072_00001  <=  0;
                end else begin
                    conv_qin_00072_00001  <=  ~tout_00072_00001 + 1;
                    sign_qin_00072_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00072 == conv_Sgntin_row_00072_00002 ) begin
                    conv_qin_00072_00002  <= tout_00072_00002;
                    sign_qin_00072_00002  <=  0;
                end else begin
                    conv_qin_00072_00002  <=  ~tout_00072_00002 + 1;
                    sign_qin_00072_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00072 == conv_Sgntin_row_00072_00003 ) begin
                    conv_qin_00072_00003  <= tout_00072_00003;
                    sign_qin_00072_00003  <=  0;
                end else begin
                    conv_qin_00072_00003  <=  ~tout_00072_00003 + 1;
                    sign_qin_00072_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00073 == conv_Sgntin_row_00073_00000 ) begin
                    conv_qin_00073_00000  <= tout_00073_00000;
                    sign_qin_00073_00000  <=  0;
                end else begin
                    conv_qin_00073_00000  <=  ~tout_00073_00000 + 1;
                    sign_qin_00073_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00073 == conv_Sgntin_row_00073_00001 ) begin
                    conv_qin_00073_00001  <= tout_00073_00001;
                    sign_qin_00073_00001  <=  0;
                end else begin
                    conv_qin_00073_00001  <=  ~tout_00073_00001 + 1;
                    sign_qin_00073_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00073 == conv_Sgntin_row_00073_00002 ) begin
                    conv_qin_00073_00002  <= tout_00073_00002;
                    sign_qin_00073_00002  <=  0;
                end else begin
                    conv_qin_00073_00002  <=  ~tout_00073_00002 + 1;
                    sign_qin_00073_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00073 == conv_Sgntin_row_00073_00003 ) begin
                    conv_qin_00073_00003  <= tout_00073_00003;
                    sign_qin_00073_00003  <=  0;
                end else begin
                    conv_qin_00073_00003  <=  ~tout_00073_00003 + 1;
                    sign_qin_00073_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00074 == conv_Sgntin_row_00074_00000 ) begin
                    conv_qin_00074_00000  <= tout_00074_00000;
                    sign_qin_00074_00000  <=  0;
                end else begin
                    conv_qin_00074_00000  <=  ~tout_00074_00000 + 1;
                    sign_qin_00074_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00074 == conv_Sgntin_row_00074_00001 ) begin
                    conv_qin_00074_00001  <= tout_00074_00001;
                    sign_qin_00074_00001  <=  0;
                end else begin
                    conv_qin_00074_00001  <=  ~tout_00074_00001 + 1;
                    sign_qin_00074_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00074 == conv_Sgntin_row_00074_00002 ) begin
                    conv_qin_00074_00002  <= tout_00074_00002;
                    sign_qin_00074_00002  <=  0;
                end else begin
                    conv_qin_00074_00002  <=  ~tout_00074_00002 + 1;
                    sign_qin_00074_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00074 == conv_Sgntin_row_00074_00003 ) begin
                    conv_qin_00074_00003  <= tout_00074_00003;
                    sign_qin_00074_00003  <=  0;
                end else begin
                    conv_qin_00074_00003  <=  ~tout_00074_00003 + 1;
                    sign_qin_00074_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00075 == conv_Sgntin_row_00075_00000 ) begin
                    conv_qin_00075_00000  <= tout_00075_00000;
                    sign_qin_00075_00000  <=  0;
                end else begin
                    conv_qin_00075_00000  <=  ~tout_00075_00000 + 1;
                    sign_qin_00075_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00075 == conv_Sgntin_row_00075_00001 ) begin
                    conv_qin_00075_00001  <= tout_00075_00001;
                    sign_qin_00075_00001  <=  0;
                end else begin
                    conv_qin_00075_00001  <=  ~tout_00075_00001 + 1;
                    sign_qin_00075_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00075 == conv_Sgntin_row_00075_00002 ) begin
                    conv_qin_00075_00002  <= tout_00075_00002;
                    sign_qin_00075_00002  <=  0;
                end else begin
                    conv_qin_00075_00002  <=  ~tout_00075_00002 + 1;
                    sign_qin_00075_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00075 == conv_Sgntin_row_00075_00003 ) begin
                    conv_qin_00075_00003  <= tout_00075_00003;
                    sign_qin_00075_00003  <=  0;
                end else begin
                    conv_qin_00075_00003  <=  ~tout_00075_00003 + 1;
                    sign_qin_00075_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00076 == conv_Sgntin_row_00076_00000 ) begin
                    conv_qin_00076_00000  <= tout_00076_00000;
                    sign_qin_00076_00000  <=  0;
                end else begin
                    conv_qin_00076_00000  <=  ~tout_00076_00000 + 1;
                    sign_qin_00076_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00076 == conv_Sgntin_row_00076_00001 ) begin
                    conv_qin_00076_00001  <= tout_00076_00001;
                    sign_qin_00076_00001  <=  0;
                end else begin
                    conv_qin_00076_00001  <=  ~tout_00076_00001 + 1;
                    sign_qin_00076_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00076 == conv_Sgntin_row_00076_00002 ) begin
                    conv_qin_00076_00002  <= tout_00076_00002;
                    sign_qin_00076_00002  <=  0;
                end else begin
                    conv_qin_00076_00002  <=  ~tout_00076_00002 + 1;
                    sign_qin_00076_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00076 == conv_Sgntin_row_00076_00003 ) begin
                    conv_qin_00076_00003  <= tout_00076_00003;
                    sign_qin_00076_00003  <=  0;
                end else begin
                    conv_qin_00076_00003  <=  ~tout_00076_00003 + 1;
                    sign_qin_00076_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00077 == conv_Sgntin_row_00077_00000 ) begin
                    conv_qin_00077_00000  <= tout_00077_00000;
                    sign_qin_00077_00000  <=  0;
                end else begin
                    conv_qin_00077_00000  <=  ~tout_00077_00000 + 1;
                    sign_qin_00077_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00077 == conv_Sgntin_row_00077_00001 ) begin
                    conv_qin_00077_00001  <= tout_00077_00001;
                    sign_qin_00077_00001  <=  0;
                end else begin
                    conv_qin_00077_00001  <=  ~tout_00077_00001 + 1;
                    sign_qin_00077_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00077 == conv_Sgntin_row_00077_00002 ) begin
                    conv_qin_00077_00002  <= tout_00077_00002;
                    sign_qin_00077_00002  <=  0;
                end else begin
                    conv_qin_00077_00002  <=  ~tout_00077_00002 + 1;
                    sign_qin_00077_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00077 == conv_Sgntin_row_00077_00003 ) begin
                    conv_qin_00077_00003  <= tout_00077_00003;
                    sign_qin_00077_00003  <=  0;
                end else begin
                    conv_qin_00077_00003  <=  ~tout_00077_00003 + 1;
                    sign_qin_00077_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00078 == conv_Sgntin_row_00078_00000 ) begin
                    conv_qin_00078_00000  <= tout_00078_00000;
                    sign_qin_00078_00000  <=  0;
                end else begin
                    conv_qin_00078_00000  <=  ~tout_00078_00000 + 1;
                    sign_qin_00078_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00078 == conv_Sgntin_row_00078_00001 ) begin
                    conv_qin_00078_00001  <= tout_00078_00001;
                    sign_qin_00078_00001  <=  0;
                end else begin
                    conv_qin_00078_00001  <=  ~tout_00078_00001 + 1;
                    sign_qin_00078_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00078 == conv_Sgntin_row_00078_00002 ) begin
                    conv_qin_00078_00002  <= tout_00078_00002;
                    sign_qin_00078_00002  <=  0;
                end else begin
                    conv_qin_00078_00002  <=  ~tout_00078_00002 + 1;
                    sign_qin_00078_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00078 == conv_Sgntin_row_00078_00003 ) begin
                    conv_qin_00078_00003  <= tout_00078_00003;
                    sign_qin_00078_00003  <=  0;
                end else begin
                    conv_qin_00078_00003  <=  ~tout_00078_00003 + 1;
                    sign_qin_00078_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00079 == conv_Sgntin_row_00079_00000 ) begin
                    conv_qin_00079_00000  <= tout_00079_00000;
                    sign_qin_00079_00000  <=  0;
                end else begin
                    conv_qin_00079_00000  <=  ~tout_00079_00000 + 1;
                    sign_qin_00079_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00079 == conv_Sgntin_row_00079_00001 ) begin
                    conv_qin_00079_00001  <= tout_00079_00001;
                    sign_qin_00079_00001  <=  0;
                end else begin
                    conv_qin_00079_00001  <=  ~tout_00079_00001 + 1;
                    sign_qin_00079_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00079 == conv_Sgntin_row_00079_00002 ) begin
                    conv_qin_00079_00002  <= tout_00079_00002;
                    sign_qin_00079_00002  <=  0;
                end else begin
                    conv_qin_00079_00002  <=  ~tout_00079_00002 + 1;
                    sign_qin_00079_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00079 == conv_Sgntin_row_00079_00003 ) begin
                    conv_qin_00079_00003  <= tout_00079_00003;
                    sign_qin_00079_00003  <=  0;
                end else begin
                    conv_qin_00079_00003  <=  ~tout_00079_00003 + 1;
                    sign_qin_00079_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00080 == conv_Sgntin_row_00080_00000 ) begin
                    conv_qin_00080_00000  <= tout_00080_00000;
                    sign_qin_00080_00000  <=  0;
                end else begin
                    conv_qin_00080_00000  <=  ~tout_00080_00000 + 1;
                    sign_qin_00080_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00080 == conv_Sgntin_row_00080_00001 ) begin
                    conv_qin_00080_00001  <= tout_00080_00001;
                    sign_qin_00080_00001  <=  0;
                end else begin
                    conv_qin_00080_00001  <=  ~tout_00080_00001 + 1;
                    sign_qin_00080_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00080 == conv_Sgntin_row_00080_00002 ) begin
                    conv_qin_00080_00002  <= tout_00080_00002;
                    sign_qin_00080_00002  <=  0;
                end else begin
                    conv_qin_00080_00002  <=  ~tout_00080_00002 + 1;
                    sign_qin_00080_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00080 == conv_Sgntin_row_00080_00003 ) begin
                    conv_qin_00080_00003  <= tout_00080_00003;
                    sign_qin_00080_00003  <=  0;
                end else begin
                    conv_qin_00080_00003  <=  ~tout_00080_00003 + 1;
                    sign_qin_00080_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00081 == conv_Sgntin_row_00081_00000 ) begin
                    conv_qin_00081_00000  <= tout_00081_00000;
                    sign_qin_00081_00000  <=  0;
                end else begin
                    conv_qin_00081_00000  <=  ~tout_00081_00000 + 1;
                    sign_qin_00081_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00081 == conv_Sgntin_row_00081_00001 ) begin
                    conv_qin_00081_00001  <= tout_00081_00001;
                    sign_qin_00081_00001  <=  0;
                end else begin
                    conv_qin_00081_00001  <=  ~tout_00081_00001 + 1;
                    sign_qin_00081_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00081 == conv_Sgntin_row_00081_00002 ) begin
                    conv_qin_00081_00002  <= tout_00081_00002;
                    sign_qin_00081_00002  <=  0;
                end else begin
                    conv_qin_00081_00002  <=  ~tout_00081_00002 + 1;
                    sign_qin_00081_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00081 == conv_Sgntin_row_00081_00003 ) begin
                    conv_qin_00081_00003  <= tout_00081_00003;
                    sign_qin_00081_00003  <=  0;
                end else begin
                    conv_qin_00081_00003  <=  ~tout_00081_00003 + 1;
                    sign_qin_00081_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00082 == conv_Sgntin_row_00082_00000 ) begin
                    conv_qin_00082_00000  <= tout_00082_00000;
                    sign_qin_00082_00000  <=  0;
                end else begin
                    conv_qin_00082_00000  <=  ~tout_00082_00000 + 1;
                    sign_qin_00082_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00082 == conv_Sgntin_row_00082_00001 ) begin
                    conv_qin_00082_00001  <= tout_00082_00001;
                    sign_qin_00082_00001  <=  0;
                end else begin
                    conv_qin_00082_00001  <=  ~tout_00082_00001 + 1;
                    sign_qin_00082_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00082 == conv_Sgntin_row_00082_00002 ) begin
                    conv_qin_00082_00002  <= tout_00082_00002;
                    sign_qin_00082_00002  <=  0;
                end else begin
                    conv_qin_00082_00002  <=  ~tout_00082_00002 + 1;
                    sign_qin_00082_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00082 == conv_Sgntin_row_00082_00003 ) begin
                    conv_qin_00082_00003  <= tout_00082_00003;
                    sign_qin_00082_00003  <=  0;
                end else begin
                    conv_qin_00082_00003  <=  ~tout_00082_00003 + 1;
                    sign_qin_00082_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00083 == conv_Sgntin_row_00083_00000 ) begin
                    conv_qin_00083_00000  <= tout_00083_00000;
                    sign_qin_00083_00000  <=  0;
                end else begin
                    conv_qin_00083_00000  <=  ~tout_00083_00000 + 1;
                    sign_qin_00083_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00083 == conv_Sgntin_row_00083_00001 ) begin
                    conv_qin_00083_00001  <= tout_00083_00001;
                    sign_qin_00083_00001  <=  0;
                end else begin
                    conv_qin_00083_00001  <=  ~tout_00083_00001 + 1;
                    sign_qin_00083_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00083 == conv_Sgntin_row_00083_00002 ) begin
                    conv_qin_00083_00002  <= tout_00083_00002;
                    sign_qin_00083_00002  <=  0;
                end else begin
                    conv_qin_00083_00002  <=  ~tout_00083_00002 + 1;
                    sign_qin_00083_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00083 == conv_Sgntin_row_00083_00003 ) begin
                    conv_qin_00083_00003  <= tout_00083_00003;
                    sign_qin_00083_00003  <=  0;
                end else begin
                    conv_qin_00083_00003  <=  ~tout_00083_00003 + 1;
                    sign_qin_00083_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00084 == conv_Sgntin_row_00084_00000 ) begin
                    conv_qin_00084_00000  <= tout_00084_00000;
                    sign_qin_00084_00000  <=  0;
                end else begin
                    conv_qin_00084_00000  <=  ~tout_00084_00000 + 1;
                    sign_qin_00084_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00084 == conv_Sgntin_row_00084_00001 ) begin
                    conv_qin_00084_00001  <= tout_00084_00001;
                    sign_qin_00084_00001  <=  0;
                end else begin
                    conv_qin_00084_00001  <=  ~tout_00084_00001 + 1;
                    sign_qin_00084_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00084 == conv_Sgntin_row_00084_00002 ) begin
                    conv_qin_00084_00002  <= tout_00084_00002;
                    sign_qin_00084_00002  <=  0;
                end else begin
                    conv_qin_00084_00002  <=  ~tout_00084_00002 + 1;
                    sign_qin_00084_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00084 == conv_Sgntin_row_00084_00003 ) begin
                    conv_qin_00084_00003  <= tout_00084_00003;
                    sign_qin_00084_00003  <=  0;
                end else begin
                    conv_qin_00084_00003  <=  ~tout_00084_00003 + 1;
                    sign_qin_00084_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00085 == conv_Sgntin_row_00085_00000 ) begin
                    conv_qin_00085_00000  <= tout_00085_00000;
                    sign_qin_00085_00000  <=  0;
                end else begin
                    conv_qin_00085_00000  <=  ~tout_00085_00000 + 1;
                    sign_qin_00085_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00085 == conv_Sgntin_row_00085_00001 ) begin
                    conv_qin_00085_00001  <= tout_00085_00001;
                    sign_qin_00085_00001  <=  0;
                end else begin
                    conv_qin_00085_00001  <=  ~tout_00085_00001 + 1;
                    sign_qin_00085_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00085 == conv_Sgntin_row_00085_00002 ) begin
                    conv_qin_00085_00002  <= tout_00085_00002;
                    sign_qin_00085_00002  <=  0;
                end else begin
                    conv_qin_00085_00002  <=  ~tout_00085_00002 + 1;
                    sign_qin_00085_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00085 == conv_Sgntin_row_00085_00003 ) begin
                    conv_qin_00085_00003  <= tout_00085_00003;
                    sign_qin_00085_00003  <=  0;
                end else begin
                    conv_qin_00085_00003  <=  ~tout_00085_00003 + 1;
                    sign_qin_00085_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00086 == conv_Sgntin_row_00086_00000 ) begin
                    conv_qin_00086_00000  <= tout_00086_00000;
                    sign_qin_00086_00000  <=  0;
                end else begin
                    conv_qin_00086_00000  <=  ~tout_00086_00000 + 1;
                    sign_qin_00086_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00086 == conv_Sgntin_row_00086_00001 ) begin
                    conv_qin_00086_00001  <= tout_00086_00001;
                    sign_qin_00086_00001  <=  0;
                end else begin
                    conv_qin_00086_00001  <=  ~tout_00086_00001 + 1;
                    sign_qin_00086_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00086 == conv_Sgntin_row_00086_00002 ) begin
                    conv_qin_00086_00002  <= tout_00086_00002;
                    sign_qin_00086_00002  <=  0;
                end else begin
                    conv_qin_00086_00002  <=  ~tout_00086_00002 + 1;
                    sign_qin_00086_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00086 == conv_Sgntin_row_00086_00003 ) begin
                    conv_qin_00086_00003  <= tout_00086_00003;
                    sign_qin_00086_00003  <=  0;
                end else begin
                    conv_qin_00086_00003  <=  ~tout_00086_00003 + 1;
                    sign_qin_00086_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00087 == conv_Sgntin_row_00087_00000 ) begin
                    conv_qin_00087_00000  <= tout_00087_00000;
                    sign_qin_00087_00000  <=  0;
                end else begin
                    conv_qin_00087_00000  <=  ~tout_00087_00000 + 1;
                    sign_qin_00087_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00087 == conv_Sgntin_row_00087_00001 ) begin
                    conv_qin_00087_00001  <= tout_00087_00001;
                    sign_qin_00087_00001  <=  0;
                end else begin
                    conv_qin_00087_00001  <=  ~tout_00087_00001 + 1;
                    sign_qin_00087_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00087 == conv_Sgntin_row_00087_00002 ) begin
                    conv_qin_00087_00002  <= tout_00087_00002;
                    sign_qin_00087_00002  <=  0;
                end else begin
                    conv_qin_00087_00002  <=  ~tout_00087_00002 + 1;
                    sign_qin_00087_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00087 == conv_Sgntin_row_00087_00003 ) begin
                    conv_qin_00087_00003  <= tout_00087_00003;
                    sign_qin_00087_00003  <=  0;
                end else begin
                    conv_qin_00087_00003  <=  ~tout_00087_00003 + 1;
                    sign_qin_00087_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00088 == conv_Sgntin_row_00088_00000 ) begin
                    conv_qin_00088_00000  <= tout_00088_00000;
                    sign_qin_00088_00000  <=  0;
                end else begin
                    conv_qin_00088_00000  <=  ~tout_00088_00000 + 1;
                    sign_qin_00088_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00088 == conv_Sgntin_row_00088_00001 ) begin
                    conv_qin_00088_00001  <= tout_00088_00001;
                    sign_qin_00088_00001  <=  0;
                end else begin
                    conv_qin_00088_00001  <=  ~tout_00088_00001 + 1;
                    sign_qin_00088_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00088 == conv_Sgntin_row_00088_00002 ) begin
                    conv_qin_00088_00002  <= tout_00088_00002;
                    sign_qin_00088_00002  <=  0;
                end else begin
                    conv_qin_00088_00002  <=  ~tout_00088_00002 + 1;
                    sign_qin_00088_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00089 == conv_Sgntin_row_00089_00000 ) begin
                    conv_qin_00089_00000  <= tout_00089_00000;
                    sign_qin_00089_00000  <=  0;
                end else begin
                    conv_qin_00089_00000  <=  ~tout_00089_00000 + 1;
                    sign_qin_00089_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00089 == conv_Sgntin_row_00089_00001 ) begin
                    conv_qin_00089_00001  <= tout_00089_00001;
                    sign_qin_00089_00001  <=  0;
                end else begin
                    conv_qin_00089_00001  <=  ~tout_00089_00001 + 1;
                    sign_qin_00089_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00089 == conv_Sgntin_row_00089_00002 ) begin
                    conv_qin_00089_00002  <= tout_00089_00002;
                    sign_qin_00089_00002  <=  0;
                end else begin
                    conv_qin_00089_00002  <=  ~tout_00089_00002 + 1;
                    sign_qin_00089_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00090 == conv_Sgntin_row_00090_00000 ) begin
                    conv_qin_00090_00000  <= tout_00090_00000;
                    sign_qin_00090_00000  <=  0;
                end else begin
                    conv_qin_00090_00000  <=  ~tout_00090_00000 + 1;
                    sign_qin_00090_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00090 == conv_Sgntin_row_00090_00001 ) begin
                    conv_qin_00090_00001  <= tout_00090_00001;
                    sign_qin_00090_00001  <=  0;
                end else begin
                    conv_qin_00090_00001  <=  ~tout_00090_00001 + 1;
                    sign_qin_00090_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00090 == conv_Sgntin_row_00090_00002 ) begin
                    conv_qin_00090_00002  <= tout_00090_00002;
                    sign_qin_00090_00002  <=  0;
                end else begin
                    conv_qin_00090_00002  <=  ~tout_00090_00002 + 1;
                    sign_qin_00090_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00091 == conv_Sgntin_row_00091_00000 ) begin
                    conv_qin_00091_00000  <= tout_00091_00000;
                    sign_qin_00091_00000  <=  0;
                end else begin
                    conv_qin_00091_00000  <=  ~tout_00091_00000 + 1;
                    sign_qin_00091_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00091 == conv_Sgntin_row_00091_00001 ) begin
                    conv_qin_00091_00001  <= tout_00091_00001;
                    sign_qin_00091_00001  <=  0;
                end else begin
                    conv_qin_00091_00001  <=  ~tout_00091_00001 + 1;
                    sign_qin_00091_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00091 == conv_Sgntin_row_00091_00002 ) begin
                    conv_qin_00091_00002  <= tout_00091_00002;
                    sign_qin_00091_00002  <=  0;
                end else begin
                    conv_qin_00091_00002  <=  ~tout_00091_00002 + 1;
                    sign_qin_00091_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00092 == conv_Sgntin_row_00092_00000 ) begin
                    conv_qin_00092_00000  <= tout_00092_00000;
                    sign_qin_00092_00000  <=  0;
                end else begin
                    conv_qin_00092_00000  <=  ~tout_00092_00000 + 1;
                    sign_qin_00092_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00092 == conv_Sgntin_row_00092_00001 ) begin
                    conv_qin_00092_00001  <= tout_00092_00001;
                    sign_qin_00092_00001  <=  0;
                end else begin
                    conv_qin_00092_00001  <=  ~tout_00092_00001 + 1;
                    sign_qin_00092_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00092 == conv_Sgntin_row_00092_00002 ) begin
                    conv_qin_00092_00002  <= tout_00092_00002;
                    sign_qin_00092_00002  <=  0;
                end else begin
                    conv_qin_00092_00002  <=  ~tout_00092_00002 + 1;
                    sign_qin_00092_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00092 == conv_Sgntin_row_00092_00003 ) begin
                    conv_qin_00092_00003  <= tout_00092_00003;
                    sign_qin_00092_00003  <=  0;
                end else begin
                    conv_qin_00092_00003  <=  ~tout_00092_00003 + 1;
                    sign_qin_00092_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00093 == conv_Sgntin_row_00093_00000 ) begin
                    conv_qin_00093_00000  <= tout_00093_00000;
                    sign_qin_00093_00000  <=  0;
                end else begin
                    conv_qin_00093_00000  <=  ~tout_00093_00000 + 1;
                    sign_qin_00093_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00093 == conv_Sgntin_row_00093_00001 ) begin
                    conv_qin_00093_00001  <= tout_00093_00001;
                    sign_qin_00093_00001  <=  0;
                end else begin
                    conv_qin_00093_00001  <=  ~tout_00093_00001 + 1;
                    sign_qin_00093_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00093 == conv_Sgntin_row_00093_00002 ) begin
                    conv_qin_00093_00002  <= tout_00093_00002;
                    sign_qin_00093_00002  <=  0;
                end else begin
                    conv_qin_00093_00002  <=  ~tout_00093_00002 + 1;
                    sign_qin_00093_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00093 == conv_Sgntin_row_00093_00003 ) begin
                    conv_qin_00093_00003  <= tout_00093_00003;
                    sign_qin_00093_00003  <=  0;
                end else begin
                    conv_qin_00093_00003  <=  ~tout_00093_00003 + 1;
                    sign_qin_00093_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00094 == conv_Sgntin_row_00094_00000 ) begin
                    conv_qin_00094_00000  <= tout_00094_00000;
                    sign_qin_00094_00000  <=  0;
                end else begin
                    conv_qin_00094_00000  <=  ~tout_00094_00000 + 1;
                    sign_qin_00094_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00094 == conv_Sgntin_row_00094_00001 ) begin
                    conv_qin_00094_00001  <= tout_00094_00001;
                    sign_qin_00094_00001  <=  0;
                end else begin
                    conv_qin_00094_00001  <=  ~tout_00094_00001 + 1;
                    sign_qin_00094_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00094 == conv_Sgntin_row_00094_00002 ) begin
                    conv_qin_00094_00002  <= tout_00094_00002;
                    sign_qin_00094_00002  <=  0;
                end else begin
                    conv_qin_00094_00002  <=  ~tout_00094_00002 + 1;
                    sign_qin_00094_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00094 == conv_Sgntin_row_00094_00003 ) begin
                    conv_qin_00094_00003  <= tout_00094_00003;
                    sign_qin_00094_00003  <=  0;
                end else begin
                    conv_qin_00094_00003  <=  ~tout_00094_00003 + 1;
                    sign_qin_00094_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00095 == conv_Sgntin_row_00095_00000 ) begin
                    conv_qin_00095_00000  <= tout_00095_00000;
                    sign_qin_00095_00000  <=  0;
                end else begin
                    conv_qin_00095_00000  <=  ~tout_00095_00000 + 1;
                    sign_qin_00095_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00095 == conv_Sgntin_row_00095_00001 ) begin
                    conv_qin_00095_00001  <= tout_00095_00001;
                    sign_qin_00095_00001  <=  0;
                end else begin
                    conv_qin_00095_00001  <=  ~tout_00095_00001 + 1;
                    sign_qin_00095_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00095 == conv_Sgntin_row_00095_00002 ) begin
                    conv_qin_00095_00002  <= tout_00095_00002;
                    sign_qin_00095_00002  <=  0;
                end else begin
                    conv_qin_00095_00002  <=  ~tout_00095_00002 + 1;
                    sign_qin_00095_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00095 == conv_Sgntin_row_00095_00003 ) begin
                    conv_qin_00095_00003  <= tout_00095_00003;
                    sign_qin_00095_00003  <=  0;
                end else begin
                    conv_qin_00095_00003  <=  ~tout_00095_00003 + 1;
                    sign_qin_00095_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00096 == conv_Sgntin_row_00096_00000 ) begin
                    conv_qin_00096_00000  <= tout_00096_00000;
                    sign_qin_00096_00000  <=  0;
                end else begin
                    conv_qin_00096_00000  <=  ~tout_00096_00000 + 1;
                    sign_qin_00096_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00096 == conv_Sgntin_row_00096_00001 ) begin
                    conv_qin_00096_00001  <= tout_00096_00001;
                    sign_qin_00096_00001  <=  0;
                end else begin
                    conv_qin_00096_00001  <=  ~tout_00096_00001 + 1;
                    sign_qin_00096_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00096 == conv_Sgntin_row_00096_00002 ) begin
                    conv_qin_00096_00002  <= tout_00096_00002;
                    sign_qin_00096_00002  <=  0;
                end else begin
                    conv_qin_00096_00002  <=  ~tout_00096_00002 + 1;
                    sign_qin_00096_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00096 == conv_Sgntin_row_00096_00003 ) begin
                    conv_qin_00096_00003  <= tout_00096_00003;
                    sign_qin_00096_00003  <=  0;
                end else begin
                    conv_qin_00096_00003  <=  ~tout_00096_00003 + 1;
                    sign_qin_00096_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00097 == conv_Sgntin_row_00097_00000 ) begin
                    conv_qin_00097_00000  <= tout_00097_00000;
                    sign_qin_00097_00000  <=  0;
                end else begin
                    conv_qin_00097_00000  <=  ~tout_00097_00000 + 1;
                    sign_qin_00097_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00097 == conv_Sgntin_row_00097_00001 ) begin
                    conv_qin_00097_00001  <= tout_00097_00001;
                    sign_qin_00097_00001  <=  0;
                end else begin
                    conv_qin_00097_00001  <=  ~tout_00097_00001 + 1;
                    sign_qin_00097_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00097 == conv_Sgntin_row_00097_00002 ) begin
                    conv_qin_00097_00002  <= tout_00097_00002;
                    sign_qin_00097_00002  <=  0;
                end else begin
                    conv_qin_00097_00002  <=  ~tout_00097_00002 + 1;
                    sign_qin_00097_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00097 == conv_Sgntin_row_00097_00003 ) begin
                    conv_qin_00097_00003  <= tout_00097_00003;
                    sign_qin_00097_00003  <=  0;
                end else begin
                    conv_qin_00097_00003  <=  ~tout_00097_00003 + 1;
                    sign_qin_00097_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00098 == conv_Sgntin_row_00098_00000 ) begin
                    conv_qin_00098_00000  <= tout_00098_00000;
                    sign_qin_00098_00000  <=  0;
                end else begin
                    conv_qin_00098_00000  <=  ~tout_00098_00000 + 1;
                    sign_qin_00098_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00098 == conv_Sgntin_row_00098_00001 ) begin
                    conv_qin_00098_00001  <= tout_00098_00001;
                    sign_qin_00098_00001  <=  0;
                end else begin
                    conv_qin_00098_00001  <=  ~tout_00098_00001 + 1;
                    sign_qin_00098_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00098 == conv_Sgntin_row_00098_00002 ) begin
                    conv_qin_00098_00002  <= tout_00098_00002;
                    sign_qin_00098_00002  <=  0;
                end else begin
                    conv_qin_00098_00002  <=  ~tout_00098_00002 + 1;
                    sign_qin_00098_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00098 == conv_Sgntin_row_00098_00003 ) begin
                    conv_qin_00098_00003  <= tout_00098_00003;
                    sign_qin_00098_00003  <=  0;
                end else begin
                    conv_qin_00098_00003  <=  ~tout_00098_00003 + 1;
                    sign_qin_00098_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00099 == conv_Sgntin_row_00099_00000 ) begin
                    conv_qin_00099_00000  <= tout_00099_00000;
                    sign_qin_00099_00000  <=  0;
                end else begin
                    conv_qin_00099_00000  <=  ~tout_00099_00000 + 1;
                    sign_qin_00099_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00099 == conv_Sgntin_row_00099_00001 ) begin
                    conv_qin_00099_00001  <= tout_00099_00001;
                    sign_qin_00099_00001  <=  0;
                end else begin
                    conv_qin_00099_00001  <=  ~tout_00099_00001 + 1;
                    sign_qin_00099_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00099 == conv_Sgntin_row_00099_00002 ) begin
                    conv_qin_00099_00002  <= tout_00099_00002;
                    sign_qin_00099_00002  <=  0;
                end else begin
                    conv_qin_00099_00002  <=  ~tout_00099_00002 + 1;
                    sign_qin_00099_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00099 == conv_Sgntin_row_00099_00003 ) begin
                    conv_qin_00099_00003  <= tout_00099_00003;
                    sign_qin_00099_00003  <=  0;
                end else begin
                    conv_qin_00099_00003  <=  ~tout_00099_00003 + 1;
                    sign_qin_00099_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00100 == conv_Sgntin_row_00100_00000 ) begin
                    conv_qin_00100_00000  <= tout_00100_00000;
                    sign_qin_00100_00000  <=  0;
                end else begin
                    conv_qin_00100_00000  <=  ~tout_00100_00000 + 1;
                    sign_qin_00100_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00100 == conv_Sgntin_row_00100_00001 ) begin
                    conv_qin_00100_00001  <= tout_00100_00001;
                    sign_qin_00100_00001  <=  0;
                end else begin
                    conv_qin_00100_00001  <=  ~tout_00100_00001 + 1;
                    sign_qin_00100_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00100 == conv_Sgntin_row_00100_00002 ) begin
                    conv_qin_00100_00002  <= tout_00100_00002;
                    sign_qin_00100_00002  <=  0;
                end else begin
                    conv_qin_00100_00002  <=  ~tout_00100_00002 + 1;
                    sign_qin_00100_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00101 == conv_Sgntin_row_00101_00000 ) begin
                    conv_qin_00101_00000  <= tout_00101_00000;
                    sign_qin_00101_00000  <=  0;
                end else begin
                    conv_qin_00101_00000  <=  ~tout_00101_00000 + 1;
                    sign_qin_00101_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00101 == conv_Sgntin_row_00101_00001 ) begin
                    conv_qin_00101_00001  <= tout_00101_00001;
                    sign_qin_00101_00001  <=  0;
                end else begin
                    conv_qin_00101_00001  <=  ~tout_00101_00001 + 1;
                    sign_qin_00101_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00101 == conv_Sgntin_row_00101_00002 ) begin
                    conv_qin_00101_00002  <= tout_00101_00002;
                    sign_qin_00101_00002  <=  0;
                end else begin
                    conv_qin_00101_00002  <=  ~tout_00101_00002 + 1;
                    sign_qin_00101_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00102 == conv_Sgntin_row_00102_00000 ) begin
                    conv_qin_00102_00000  <= tout_00102_00000;
                    sign_qin_00102_00000  <=  0;
                end else begin
                    conv_qin_00102_00000  <=  ~tout_00102_00000 + 1;
                    sign_qin_00102_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00102 == conv_Sgntin_row_00102_00001 ) begin
                    conv_qin_00102_00001  <= tout_00102_00001;
                    sign_qin_00102_00001  <=  0;
                end else begin
                    conv_qin_00102_00001  <=  ~tout_00102_00001 + 1;
                    sign_qin_00102_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00102 == conv_Sgntin_row_00102_00002 ) begin
                    conv_qin_00102_00002  <= tout_00102_00002;
                    sign_qin_00102_00002  <=  0;
                end else begin
                    conv_qin_00102_00002  <=  ~tout_00102_00002 + 1;
                    sign_qin_00102_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00103 == conv_Sgntin_row_00103_00000 ) begin
                    conv_qin_00103_00000  <= tout_00103_00000;
                    sign_qin_00103_00000  <=  0;
                end else begin
                    conv_qin_00103_00000  <=  ~tout_00103_00000 + 1;
                    sign_qin_00103_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00103 == conv_Sgntin_row_00103_00001 ) begin
                    conv_qin_00103_00001  <= tout_00103_00001;
                    sign_qin_00103_00001  <=  0;
                end else begin
                    conv_qin_00103_00001  <=  ~tout_00103_00001 + 1;
                    sign_qin_00103_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00103 == conv_Sgntin_row_00103_00002 ) begin
                    conv_qin_00103_00002  <= tout_00103_00002;
                    sign_qin_00103_00002  <=  0;
                end else begin
                    conv_qin_00103_00002  <=  ~tout_00103_00002 + 1;
                    sign_qin_00103_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00104 == conv_Sgntin_row_00104_00000 ) begin
                    conv_qin_00104_00000  <= tout_00104_00000;
                    sign_qin_00104_00000  <=  0;
                end else begin
                    conv_qin_00104_00000  <=  ~tout_00104_00000 + 1;
                    sign_qin_00104_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00104 == conv_Sgntin_row_00104_00001 ) begin
                    conv_qin_00104_00001  <= tout_00104_00001;
                    sign_qin_00104_00001  <=  0;
                end else begin
                    conv_qin_00104_00001  <=  ~tout_00104_00001 + 1;
                    sign_qin_00104_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00104 == conv_Sgntin_row_00104_00002 ) begin
                    conv_qin_00104_00002  <= tout_00104_00002;
                    sign_qin_00104_00002  <=  0;
                end else begin
                    conv_qin_00104_00002  <=  ~tout_00104_00002 + 1;
                    sign_qin_00104_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00104 == conv_Sgntin_row_00104_00003 ) begin
                    conv_qin_00104_00003  <= tout_00104_00003;
                    sign_qin_00104_00003  <=  0;
                end else begin
                    conv_qin_00104_00003  <=  ~tout_00104_00003 + 1;
                    sign_qin_00104_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00104 == conv_Sgntin_row_00104_00004 ) begin
                    conv_qin_00104_00004  <= tout_00104_00004;
                    sign_qin_00104_00004  <=  0;
                end else begin
                    conv_qin_00104_00004  <=  ~tout_00104_00004 + 1;
                    sign_qin_00104_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00105 == conv_Sgntin_row_00105_00000 ) begin
                    conv_qin_00105_00000  <= tout_00105_00000;
                    sign_qin_00105_00000  <=  0;
                end else begin
                    conv_qin_00105_00000  <=  ~tout_00105_00000 + 1;
                    sign_qin_00105_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00105 == conv_Sgntin_row_00105_00001 ) begin
                    conv_qin_00105_00001  <= tout_00105_00001;
                    sign_qin_00105_00001  <=  0;
                end else begin
                    conv_qin_00105_00001  <=  ~tout_00105_00001 + 1;
                    sign_qin_00105_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00105 == conv_Sgntin_row_00105_00002 ) begin
                    conv_qin_00105_00002  <= tout_00105_00002;
                    sign_qin_00105_00002  <=  0;
                end else begin
                    conv_qin_00105_00002  <=  ~tout_00105_00002 + 1;
                    sign_qin_00105_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00105 == conv_Sgntin_row_00105_00003 ) begin
                    conv_qin_00105_00003  <= tout_00105_00003;
                    sign_qin_00105_00003  <=  0;
                end else begin
                    conv_qin_00105_00003  <=  ~tout_00105_00003 + 1;
                    sign_qin_00105_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00105 == conv_Sgntin_row_00105_00004 ) begin
                    conv_qin_00105_00004  <= tout_00105_00004;
                    sign_qin_00105_00004  <=  0;
                end else begin
                    conv_qin_00105_00004  <=  ~tout_00105_00004 + 1;
                    sign_qin_00105_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00106 == conv_Sgntin_row_00106_00000 ) begin
                    conv_qin_00106_00000  <= tout_00106_00000;
                    sign_qin_00106_00000  <=  0;
                end else begin
                    conv_qin_00106_00000  <=  ~tout_00106_00000 + 1;
                    sign_qin_00106_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00106 == conv_Sgntin_row_00106_00001 ) begin
                    conv_qin_00106_00001  <= tout_00106_00001;
                    sign_qin_00106_00001  <=  0;
                end else begin
                    conv_qin_00106_00001  <=  ~tout_00106_00001 + 1;
                    sign_qin_00106_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00106 == conv_Sgntin_row_00106_00002 ) begin
                    conv_qin_00106_00002  <= tout_00106_00002;
                    sign_qin_00106_00002  <=  0;
                end else begin
                    conv_qin_00106_00002  <=  ~tout_00106_00002 + 1;
                    sign_qin_00106_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00106 == conv_Sgntin_row_00106_00003 ) begin
                    conv_qin_00106_00003  <= tout_00106_00003;
                    sign_qin_00106_00003  <=  0;
                end else begin
                    conv_qin_00106_00003  <=  ~tout_00106_00003 + 1;
                    sign_qin_00106_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00106 == conv_Sgntin_row_00106_00004 ) begin
                    conv_qin_00106_00004  <= tout_00106_00004;
                    sign_qin_00106_00004  <=  0;
                end else begin
                    conv_qin_00106_00004  <=  ~tout_00106_00004 + 1;
                    sign_qin_00106_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00107 == conv_Sgntin_row_00107_00000 ) begin
                    conv_qin_00107_00000  <= tout_00107_00000;
                    sign_qin_00107_00000  <=  0;
                end else begin
                    conv_qin_00107_00000  <=  ~tout_00107_00000 + 1;
                    sign_qin_00107_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00107 == conv_Sgntin_row_00107_00001 ) begin
                    conv_qin_00107_00001  <= tout_00107_00001;
                    sign_qin_00107_00001  <=  0;
                end else begin
                    conv_qin_00107_00001  <=  ~tout_00107_00001 + 1;
                    sign_qin_00107_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00107 == conv_Sgntin_row_00107_00002 ) begin
                    conv_qin_00107_00002  <= tout_00107_00002;
                    sign_qin_00107_00002  <=  0;
                end else begin
                    conv_qin_00107_00002  <=  ~tout_00107_00002 + 1;
                    sign_qin_00107_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00107 == conv_Sgntin_row_00107_00003 ) begin
                    conv_qin_00107_00003  <= tout_00107_00003;
                    sign_qin_00107_00003  <=  0;
                end else begin
                    conv_qin_00107_00003  <=  ~tout_00107_00003 + 1;
                    sign_qin_00107_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00107 == conv_Sgntin_row_00107_00004 ) begin
                    conv_qin_00107_00004  <= tout_00107_00004;
                    sign_qin_00107_00004  <=  0;
                end else begin
                    conv_qin_00107_00004  <=  ~tout_00107_00004 + 1;
                    sign_qin_00107_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00108 == conv_Sgntin_row_00108_00000 ) begin
                    conv_qin_00108_00000  <= tout_00108_00000;
                    sign_qin_00108_00000  <=  0;
                end else begin
                    conv_qin_00108_00000  <=  ~tout_00108_00000 + 1;
                    sign_qin_00108_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00108 == conv_Sgntin_row_00108_00001 ) begin
                    conv_qin_00108_00001  <= tout_00108_00001;
                    sign_qin_00108_00001  <=  0;
                end else begin
                    conv_qin_00108_00001  <=  ~tout_00108_00001 + 1;
                    sign_qin_00108_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00108 == conv_Sgntin_row_00108_00002 ) begin
                    conv_qin_00108_00002  <= tout_00108_00002;
                    sign_qin_00108_00002  <=  0;
                end else begin
                    conv_qin_00108_00002  <=  ~tout_00108_00002 + 1;
                    sign_qin_00108_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00109 == conv_Sgntin_row_00109_00000 ) begin
                    conv_qin_00109_00000  <= tout_00109_00000;
                    sign_qin_00109_00000  <=  0;
                end else begin
                    conv_qin_00109_00000  <=  ~tout_00109_00000 + 1;
                    sign_qin_00109_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00109 == conv_Sgntin_row_00109_00001 ) begin
                    conv_qin_00109_00001  <= tout_00109_00001;
                    sign_qin_00109_00001  <=  0;
                end else begin
                    conv_qin_00109_00001  <=  ~tout_00109_00001 + 1;
                    sign_qin_00109_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00109 == conv_Sgntin_row_00109_00002 ) begin
                    conv_qin_00109_00002  <= tout_00109_00002;
                    sign_qin_00109_00002  <=  0;
                end else begin
                    conv_qin_00109_00002  <=  ~tout_00109_00002 + 1;
                    sign_qin_00109_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00110 == conv_Sgntin_row_00110_00000 ) begin
                    conv_qin_00110_00000  <= tout_00110_00000;
                    sign_qin_00110_00000  <=  0;
                end else begin
                    conv_qin_00110_00000  <=  ~tout_00110_00000 + 1;
                    sign_qin_00110_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00110 == conv_Sgntin_row_00110_00001 ) begin
                    conv_qin_00110_00001  <= tout_00110_00001;
                    sign_qin_00110_00001  <=  0;
                end else begin
                    conv_qin_00110_00001  <=  ~tout_00110_00001 + 1;
                    sign_qin_00110_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00110 == conv_Sgntin_row_00110_00002 ) begin
                    conv_qin_00110_00002  <= tout_00110_00002;
                    sign_qin_00110_00002  <=  0;
                end else begin
                    conv_qin_00110_00002  <=  ~tout_00110_00002 + 1;
                    sign_qin_00110_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00111 == conv_Sgntin_row_00111_00000 ) begin
                    conv_qin_00111_00000  <= tout_00111_00000;
                    sign_qin_00111_00000  <=  0;
                end else begin
                    conv_qin_00111_00000  <=  ~tout_00111_00000 + 1;
                    sign_qin_00111_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00111 == conv_Sgntin_row_00111_00001 ) begin
                    conv_qin_00111_00001  <= tout_00111_00001;
                    sign_qin_00111_00001  <=  0;
                end else begin
                    conv_qin_00111_00001  <=  ~tout_00111_00001 + 1;
                    sign_qin_00111_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00111 == conv_Sgntin_row_00111_00002 ) begin
                    conv_qin_00111_00002  <= tout_00111_00002;
                    sign_qin_00111_00002  <=  0;
                end else begin
                    conv_qin_00111_00002  <=  ~tout_00111_00002 + 1;
                    sign_qin_00111_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00112 == conv_Sgntin_row_00112_00000 ) begin
                    conv_qin_00112_00000  <= tout_00112_00000;
                    sign_qin_00112_00000  <=  0;
                end else begin
                    conv_qin_00112_00000  <=  ~tout_00112_00000 + 1;
                    sign_qin_00112_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00112 == conv_Sgntin_row_00112_00001 ) begin
                    conv_qin_00112_00001  <= tout_00112_00001;
                    sign_qin_00112_00001  <=  0;
                end else begin
                    conv_qin_00112_00001  <=  ~tout_00112_00001 + 1;
                    sign_qin_00112_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00112 == conv_Sgntin_row_00112_00002 ) begin
                    conv_qin_00112_00002  <= tout_00112_00002;
                    sign_qin_00112_00002  <=  0;
                end else begin
                    conv_qin_00112_00002  <=  ~tout_00112_00002 + 1;
                    sign_qin_00112_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00112 == conv_Sgntin_row_00112_00003 ) begin
                    conv_qin_00112_00003  <= tout_00112_00003;
                    sign_qin_00112_00003  <=  0;
                end else begin
                    conv_qin_00112_00003  <=  ~tout_00112_00003 + 1;
                    sign_qin_00112_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00113 == conv_Sgntin_row_00113_00000 ) begin
                    conv_qin_00113_00000  <= tout_00113_00000;
                    sign_qin_00113_00000  <=  0;
                end else begin
                    conv_qin_00113_00000  <=  ~tout_00113_00000 + 1;
                    sign_qin_00113_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00113 == conv_Sgntin_row_00113_00001 ) begin
                    conv_qin_00113_00001  <= tout_00113_00001;
                    sign_qin_00113_00001  <=  0;
                end else begin
                    conv_qin_00113_00001  <=  ~tout_00113_00001 + 1;
                    sign_qin_00113_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00113 == conv_Sgntin_row_00113_00002 ) begin
                    conv_qin_00113_00002  <= tout_00113_00002;
                    sign_qin_00113_00002  <=  0;
                end else begin
                    conv_qin_00113_00002  <=  ~tout_00113_00002 + 1;
                    sign_qin_00113_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00113 == conv_Sgntin_row_00113_00003 ) begin
                    conv_qin_00113_00003  <= tout_00113_00003;
                    sign_qin_00113_00003  <=  0;
                end else begin
                    conv_qin_00113_00003  <=  ~tout_00113_00003 + 1;
                    sign_qin_00113_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00114 == conv_Sgntin_row_00114_00000 ) begin
                    conv_qin_00114_00000  <= tout_00114_00000;
                    sign_qin_00114_00000  <=  0;
                end else begin
                    conv_qin_00114_00000  <=  ~tout_00114_00000 + 1;
                    sign_qin_00114_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00114 == conv_Sgntin_row_00114_00001 ) begin
                    conv_qin_00114_00001  <= tout_00114_00001;
                    sign_qin_00114_00001  <=  0;
                end else begin
                    conv_qin_00114_00001  <=  ~tout_00114_00001 + 1;
                    sign_qin_00114_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00114 == conv_Sgntin_row_00114_00002 ) begin
                    conv_qin_00114_00002  <= tout_00114_00002;
                    sign_qin_00114_00002  <=  0;
                end else begin
                    conv_qin_00114_00002  <=  ~tout_00114_00002 + 1;
                    sign_qin_00114_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00114 == conv_Sgntin_row_00114_00003 ) begin
                    conv_qin_00114_00003  <= tout_00114_00003;
                    sign_qin_00114_00003  <=  0;
                end else begin
                    conv_qin_00114_00003  <=  ~tout_00114_00003 + 1;
                    sign_qin_00114_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00115 == conv_Sgntin_row_00115_00000 ) begin
                    conv_qin_00115_00000  <= tout_00115_00000;
                    sign_qin_00115_00000  <=  0;
                end else begin
                    conv_qin_00115_00000  <=  ~tout_00115_00000 + 1;
                    sign_qin_00115_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00115 == conv_Sgntin_row_00115_00001 ) begin
                    conv_qin_00115_00001  <= tout_00115_00001;
                    sign_qin_00115_00001  <=  0;
                end else begin
                    conv_qin_00115_00001  <=  ~tout_00115_00001 + 1;
                    sign_qin_00115_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00115 == conv_Sgntin_row_00115_00002 ) begin
                    conv_qin_00115_00002  <= tout_00115_00002;
                    sign_qin_00115_00002  <=  0;
                end else begin
                    conv_qin_00115_00002  <=  ~tout_00115_00002 + 1;
                    sign_qin_00115_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00115 == conv_Sgntin_row_00115_00003 ) begin
                    conv_qin_00115_00003  <= tout_00115_00003;
                    sign_qin_00115_00003  <=  0;
                end else begin
                    conv_qin_00115_00003  <=  ~tout_00115_00003 + 1;
                    sign_qin_00115_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00116 == conv_Sgntin_row_00116_00000 ) begin
                    conv_qin_00116_00000  <= tout_00116_00000;
                    sign_qin_00116_00000  <=  0;
                end else begin
                    conv_qin_00116_00000  <=  ~tout_00116_00000 + 1;
                    sign_qin_00116_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00116 == conv_Sgntin_row_00116_00001 ) begin
                    conv_qin_00116_00001  <= tout_00116_00001;
                    sign_qin_00116_00001  <=  0;
                end else begin
                    conv_qin_00116_00001  <=  ~tout_00116_00001 + 1;
                    sign_qin_00116_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00116 == conv_Sgntin_row_00116_00002 ) begin
                    conv_qin_00116_00002  <= tout_00116_00002;
                    sign_qin_00116_00002  <=  0;
                end else begin
                    conv_qin_00116_00002  <=  ~tout_00116_00002 + 1;
                    sign_qin_00116_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00117 == conv_Sgntin_row_00117_00000 ) begin
                    conv_qin_00117_00000  <= tout_00117_00000;
                    sign_qin_00117_00000  <=  0;
                end else begin
                    conv_qin_00117_00000  <=  ~tout_00117_00000 + 1;
                    sign_qin_00117_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00117 == conv_Sgntin_row_00117_00001 ) begin
                    conv_qin_00117_00001  <= tout_00117_00001;
                    sign_qin_00117_00001  <=  0;
                end else begin
                    conv_qin_00117_00001  <=  ~tout_00117_00001 + 1;
                    sign_qin_00117_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00117 == conv_Sgntin_row_00117_00002 ) begin
                    conv_qin_00117_00002  <= tout_00117_00002;
                    sign_qin_00117_00002  <=  0;
                end else begin
                    conv_qin_00117_00002  <=  ~tout_00117_00002 + 1;
                    sign_qin_00117_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00118 == conv_Sgntin_row_00118_00000 ) begin
                    conv_qin_00118_00000  <= tout_00118_00000;
                    sign_qin_00118_00000  <=  0;
                end else begin
                    conv_qin_00118_00000  <=  ~tout_00118_00000 + 1;
                    sign_qin_00118_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00118 == conv_Sgntin_row_00118_00001 ) begin
                    conv_qin_00118_00001  <= tout_00118_00001;
                    sign_qin_00118_00001  <=  0;
                end else begin
                    conv_qin_00118_00001  <=  ~tout_00118_00001 + 1;
                    sign_qin_00118_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00118 == conv_Sgntin_row_00118_00002 ) begin
                    conv_qin_00118_00002  <= tout_00118_00002;
                    sign_qin_00118_00002  <=  0;
                end else begin
                    conv_qin_00118_00002  <=  ~tout_00118_00002 + 1;
                    sign_qin_00118_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00119 == conv_Sgntin_row_00119_00000 ) begin
                    conv_qin_00119_00000  <= tout_00119_00000;
                    sign_qin_00119_00000  <=  0;
                end else begin
                    conv_qin_00119_00000  <=  ~tout_00119_00000 + 1;
                    sign_qin_00119_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00119 == conv_Sgntin_row_00119_00001 ) begin
                    conv_qin_00119_00001  <= tout_00119_00001;
                    sign_qin_00119_00001  <=  0;
                end else begin
                    conv_qin_00119_00001  <=  ~tout_00119_00001 + 1;
                    sign_qin_00119_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00119 == conv_Sgntin_row_00119_00002 ) begin
                    conv_qin_00119_00002  <= tout_00119_00002;
                    sign_qin_00119_00002  <=  0;
                end else begin
                    conv_qin_00119_00002  <=  ~tout_00119_00002 + 1;
                    sign_qin_00119_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00120 == conv_Sgntin_row_00120_00000 ) begin
                    conv_qin_00120_00000  <= tout_00120_00000;
                    sign_qin_00120_00000  <=  0;
                end else begin
                    conv_qin_00120_00000  <=  ~tout_00120_00000 + 1;
                    sign_qin_00120_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00120 == conv_Sgntin_row_00120_00001 ) begin
                    conv_qin_00120_00001  <= tout_00120_00001;
                    sign_qin_00120_00001  <=  0;
                end else begin
                    conv_qin_00120_00001  <=  ~tout_00120_00001 + 1;
                    sign_qin_00120_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00120 == conv_Sgntin_row_00120_00002 ) begin
                    conv_qin_00120_00002  <= tout_00120_00002;
                    sign_qin_00120_00002  <=  0;
                end else begin
                    conv_qin_00120_00002  <=  ~tout_00120_00002 + 1;
                    sign_qin_00120_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00120 == conv_Sgntin_row_00120_00003 ) begin
                    conv_qin_00120_00003  <= tout_00120_00003;
                    sign_qin_00120_00003  <=  0;
                end else begin
                    conv_qin_00120_00003  <=  ~tout_00120_00003 + 1;
                    sign_qin_00120_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00120 == conv_Sgntin_row_00120_00004 ) begin
                    conv_qin_00120_00004  <= tout_00120_00004;
                    sign_qin_00120_00004  <=  0;
                end else begin
                    conv_qin_00120_00004  <=  ~tout_00120_00004 + 1;
                    sign_qin_00120_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00121 == conv_Sgntin_row_00121_00000 ) begin
                    conv_qin_00121_00000  <= tout_00121_00000;
                    sign_qin_00121_00000  <=  0;
                end else begin
                    conv_qin_00121_00000  <=  ~tout_00121_00000 + 1;
                    sign_qin_00121_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00121 == conv_Sgntin_row_00121_00001 ) begin
                    conv_qin_00121_00001  <= tout_00121_00001;
                    sign_qin_00121_00001  <=  0;
                end else begin
                    conv_qin_00121_00001  <=  ~tout_00121_00001 + 1;
                    sign_qin_00121_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00121 == conv_Sgntin_row_00121_00002 ) begin
                    conv_qin_00121_00002  <= tout_00121_00002;
                    sign_qin_00121_00002  <=  0;
                end else begin
                    conv_qin_00121_00002  <=  ~tout_00121_00002 + 1;
                    sign_qin_00121_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00121 == conv_Sgntin_row_00121_00003 ) begin
                    conv_qin_00121_00003  <= tout_00121_00003;
                    sign_qin_00121_00003  <=  0;
                end else begin
                    conv_qin_00121_00003  <=  ~tout_00121_00003 + 1;
                    sign_qin_00121_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00121 == conv_Sgntin_row_00121_00004 ) begin
                    conv_qin_00121_00004  <= tout_00121_00004;
                    sign_qin_00121_00004  <=  0;
                end else begin
                    conv_qin_00121_00004  <=  ~tout_00121_00004 + 1;
                    sign_qin_00121_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00122 == conv_Sgntin_row_00122_00000 ) begin
                    conv_qin_00122_00000  <= tout_00122_00000;
                    sign_qin_00122_00000  <=  0;
                end else begin
                    conv_qin_00122_00000  <=  ~tout_00122_00000 + 1;
                    sign_qin_00122_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00122 == conv_Sgntin_row_00122_00001 ) begin
                    conv_qin_00122_00001  <= tout_00122_00001;
                    sign_qin_00122_00001  <=  0;
                end else begin
                    conv_qin_00122_00001  <=  ~tout_00122_00001 + 1;
                    sign_qin_00122_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00122 == conv_Sgntin_row_00122_00002 ) begin
                    conv_qin_00122_00002  <= tout_00122_00002;
                    sign_qin_00122_00002  <=  0;
                end else begin
                    conv_qin_00122_00002  <=  ~tout_00122_00002 + 1;
                    sign_qin_00122_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00122 == conv_Sgntin_row_00122_00003 ) begin
                    conv_qin_00122_00003  <= tout_00122_00003;
                    sign_qin_00122_00003  <=  0;
                end else begin
                    conv_qin_00122_00003  <=  ~tout_00122_00003 + 1;
                    sign_qin_00122_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00122 == conv_Sgntin_row_00122_00004 ) begin
                    conv_qin_00122_00004  <= tout_00122_00004;
                    sign_qin_00122_00004  <=  0;
                end else begin
                    conv_qin_00122_00004  <=  ~tout_00122_00004 + 1;
                    sign_qin_00122_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00123 == conv_Sgntin_row_00123_00000 ) begin
                    conv_qin_00123_00000  <= tout_00123_00000;
                    sign_qin_00123_00000  <=  0;
                end else begin
                    conv_qin_00123_00000  <=  ~tout_00123_00000 + 1;
                    sign_qin_00123_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00123 == conv_Sgntin_row_00123_00001 ) begin
                    conv_qin_00123_00001  <= tout_00123_00001;
                    sign_qin_00123_00001  <=  0;
                end else begin
                    conv_qin_00123_00001  <=  ~tout_00123_00001 + 1;
                    sign_qin_00123_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00123 == conv_Sgntin_row_00123_00002 ) begin
                    conv_qin_00123_00002  <= tout_00123_00002;
                    sign_qin_00123_00002  <=  0;
                end else begin
                    conv_qin_00123_00002  <=  ~tout_00123_00002 + 1;
                    sign_qin_00123_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00123 == conv_Sgntin_row_00123_00003 ) begin
                    conv_qin_00123_00003  <= tout_00123_00003;
                    sign_qin_00123_00003  <=  0;
                end else begin
                    conv_qin_00123_00003  <=  ~tout_00123_00003 + 1;
                    sign_qin_00123_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00123 == conv_Sgntin_row_00123_00004 ) begin
                    conv_qin_00123_00004  <= tout_00123_00004;
                    sign_qin_00123_00004  <=  0;
                end else begin
                    conv_qin_00123_00004  <=  ~tout_00123_00004 + 1;
                    sign_qin_00123_00004  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00124 == conv_Sgntin_row_00124_00000 ) begin
                    conv_qin_00124_00000  <= tout_00124_00000;
                    sign_qin_00124_00000  <=  0;
                end else begin
                    conv_qin_00124_00000  <=  ~tout_00124_00000 + 1;
                    sign_qin_00124_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00124 == conv_Sgntin_row_00124_00001 ) begin
                    conv_qin_00124_00001  <= tout_00124_00001;
                    sign_qin_00124_00001  <=  0;
                end else begin
                    conv_qin_00124_00001  <=  ~tout_00124_00001 + 1;
                    sign_qin_00124_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00124 == conv_Sgntin_row_00124_00002 ) begin
                    conv_qin_00124_00002  <= tout_00124_00002;
                    sign_qin_00124_00002  <=  0;
                end else begin
                    conv_qin_00124_00002  <=  ~tout_00124_00002 + 1;
                    sign_qin_00124_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00125 == conv_Sgntin_row_00125_00000 ) begin
                    conv_qin_00125_00000  <= tout_00125_00000;
                    sign_qin_00125_00000  <=  0;
                end else begin
                    conv_qin_00125_00000  <=  ~tout_00125_00000 + 1;
                    sign_qin_00125_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00125 == conv_Sgntin_row_00125_00001 ) begin
                    conv_qin_00125_00001  <= tout_00125_00001;
                    sign_qin_00125_00001  <=  0;
                end else begin
                    conv_qin_00125_00001  <=  ~tout_00125_00001 + 1;
                    sign_qin_00125_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00125 == conv_Sgntin_row_00125_00002 ) begin
                    conv_qin_00125_00002  <= tout_00125_00002;
                    sign_qin_00125_00002  <=  0;
                end else begin
                    conv_qin_00125_00002  <=  ~tout_00125_00002 + 1;
                    sign_qin_00125_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00126 == conv_Sgntin_row_00126_00000 ) begin
                    conv_qin_00126_00000  <= tout_00126_00000;
                    sign_qin_00126_00000  <=  0;
                end else begin
                    conv_qin_00126_00000  <=  ~tout_00126_00000 + 1;
                    sign_qin_00126_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00126 == conv_Sgntin_row_00126_00001 ) begin
                    conv_qin_00126_00001  <= tout_00126_00001;
                    sign_qin_00126_00001  <=  0;
                end else begin
                    conv_qin_00126_00001  <=  ~tout_00126_00001 + 1;
                    sign_qin_00126_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00126 == conv_Sgntin_row_00126_00002 ) begin
                    conv_qin_00126_00002  <= tout_00126_00002;
                    sign_qin_00126_00002  <=  0;
                end else begin
                    conv_qin_00126_00002  <=  ~tout_00126_00002 + 1;
                    sign_qin_00126_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00127 == conv_Sgntin_row_00127_00000 ) begin
                    conv_qin_00127_00000  <= tout_00127_00000;
                    sign_qin_00127_00000  <=  0;
                end else begin
                    conv_qin_00127_00000  <=  ~tout_00127_00000 + 1;
                    sign_qin_00127_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00127 == conv_Sgntin_row_00127_00001 ) begin
                    conv_qin_00127_00001  <= tout_00127_00001;
                    sign_qin_00127_00001  <=  0;
                end else begin
                    conv_qin_00127_00001  <=  ~tout_00127_00001 + 1;
                    sign_qin_00127_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00127 == conv_Sgntin_row_00127_00002 ) begin
                    conv_qin_00127_00002  <= tout_00127_00002;
                    sign_qin_00127_00002  <=  0;
                end else begin
                    conv_qin_00127_00002  <=  ~tout_00127_00002 + 1;
                    sign_qin_00127_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00128 == conv_Sgntin_row_00128_00000 ) begin
                    conv_qin_00128_00000  <= tout_00128_00000;
                    sign_qin_00128_00000  <=  0;
                end else begin
                    conv_qin_00128_00000  <=  ~tout_00128_00000 + 1;
                    sign_qin_00128_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00128 == conv_Sgntin_row_00128_00001 ) begin
                    conv_qin_00128_00001  <= tout_00128_00001;
                    sign_qin_00128_00001  <=  0;
                end else begin
                    conv_qin_00128_00001  <=  ~tout_00128_00001 + 1;
                    sign_qin_00128_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00128 == conv_Sgntin_row_00128_00002 ) begin
                    conv_qin_00128_00002  <= tout_00128_00002;
                    sign_qin_00128_00002  <=  0;
                end else begin
                    conv_qin_00128_00002  <=  ~tout_00128_00002 + 1;
                    sign_qin_00128_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00128 == conv_Sgntin_row_00128_00003 ) begin
                    conv_qin_00128_00003  <= tout_00128_00003;
                    sign_qin_00128_00003  <=  0;
                end else begin
                    conv_qin_00128_00003  <=  ~tout_00128_00003 + 1;
                    sign_qin_00128_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00129 == conv_Sgntin_row_00129_00000 ) begin
                    conv_qin_00129_00000  <= tout_00129_00000;
                    sign_qin_00129_00000  <=  0;
                end else begin
                    conv_qin_00129_00000  <=  ~tout_00129_00000 + 1;
                    sign_qin_00129_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00129 == conv_Sgntin_row_00129_00001 ) begin
                    conv_qin_00129_00001  <= tout_00129_00001;
                    sign_qin_00129_00001  <=  0;
                end else begin
                    conv_qin_00129_00001  <=  ~tout_00129_00001 + 1;
                    sign_qin_00129_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00129 == conv_Sgntin_row_00129_00002 ) begin
                    conv_qin_00129_00002  <= tout_00129_00002;
                    sign_qin_00129_00002  <=  0;
                end else begin
                    conv_qin_00129_00002  <=  ~tout_00129_00002 + 1;
                    sign_qin_00129_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00129 == conv_Sgntin_row_00129_00003 ) begin
                    conv_qin_00129_00003  <= tout_00129_00003;
                    sign_qin_00129_00003  <=  0;
                end else begin
                    conv_qin_00129_00003  <=  ~tout_00129_00003 + 1;
                    sign_qin_00129_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00130 == conv_Sgntin_row_00130_00000 ) begin
                    conv_qin_00130_00000  <= tout_00130_00000;
                    sign_qin_00130_00000  <=  0;
                end else begin
                    conv_qin_00130_00000  <=  ~tout_00130_00000 + 1;
                    sign_qin_00130_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00130 == conv_Sgntin_row_00130_00001 ) begin
                    conv_qin_00130_00001  <= tout_00130_00001;
                    sign_qin_00130_00001  <=  0;
                end else begin
                    conv_qin_00130_00001  <=  ~tout_00130_00001 + 1;
                    sign_qin_00130_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00130 == conv_Sgntin_row_00130_00002 ) begin
                    conv_qin_00130_00002  <= tout_00130_00002;
                    sign_qin_00130_00002  <=  0;
                end else begin
                    conv_qin_00130_00002  <=  ~tout_00130_00002 + 1;
                    sign_qin_00130_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00130 == conv_Sgntin_row_00130_00003 ) begin
                    conv_qin_00130_00003  <= tout_00130_00003;
                    sign_qin_00130_00003  <=  0;
                end else begin
                    conv_qin_00130_00003  <=  ~tout_00130_00003 + 1;
                    sign_qin_00130_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00131 == conv_Sgntin_row_00131_00000 ) begin
                    conv_qin_00131_00000  <= tout_00131_00000;
                    sign_qin_00131_00000  <=  0;
                end else begin
                    conv_qin_00131_00000  <=  ~tout_00131_00000 + 1;
                    sign_qin_00131_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00131 == conv_Sgntin_row_00131_00001 ) begin
                    conv_qin_00131_00001  <= tout_00131_00001;
                    sign_qin_00131_00001  <=  0;
                end else begin
                    conv_qin_00131_00001  <=  ~tout_00131_00001 + 1;
                    sign_qin_00131_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00131 == conv_Sgntin_row_00131_00002 ) begin
                    conv_qin_00131_00002  <= tout_00131_00002;
                    sign_qin_00131_00002  <=  0;
                end else begin
                    conv_qin_00131_00002  <=  ~tout_00131_00002 + 1;
                    sign_qin_00131_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00131 == conv_Sgntin_row_00131_00003 ) begin
                    conv_qin_00131_00003  <= tout_00131_00003;
                    sign_qin_00131_00003  <=  0;
                end else begin
                    conv_qin_00131_00003  <=  ~tout_00131_00003 + 1;
                    sign_qin_00131_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00132 == conv_Sgntin_row_00132_00000 ) begin
                    conv_qin_00132_00000  <= tout_00132_00000;
                    sign_qin_00132_00000  <=  0;
                end else begin
                    conv_qin_00132_00000  <=  ~tout_00132_00000 + 1;
                    sign_qin_00132_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00132 == conv_Sgntin_row_00132_00001 ) begin
                    conv_qin_00132_00001  <= tout_00132_00001;
                    sign_qin_00132_00001  <=  0;
                end else begin
                    conv_qin_00132_00001  <=  ~tout_00132_00001 + 1;
                    sign_qin_00132_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00132 == conv_Sgntin_row_00132_00002 ) begin
                    conv_qin_00132_00002  <= tout_00132_00002;
                    sign_qin_00132_00002  <=  0;
                end else begin
                    conv_qin_00132_00002  <=  ~tout_00132_00002 + 1;
                    sign_qin_00132_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00132 == conv_Sgntin_row_00132_00003 ) begin
                    conv_qin_00132_00003  <= tout_00132_00003;
                    sign_qin_00132_00003  <=  0;
                end else begin
                    conv_qin_00132_00003  <=  ~tout_00132_00003 + 1;
                    sign_qin_00132_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00133 == conv_Sgntin_row_00133_00000 ) begin
                    conv_qin_00133_00000  <= tout_00133_00000;
                    sign_qin_00133_00000  <=  0;
                end else begin
                    conv_qin_00133_00000  <=  ~tout_00133_00000 + 1;
                    sign_qin_00133_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00133 == conv_Sgntin_row_00133_00001 ) begin
                    conv_qin_00133_00001  <= tout_00133_00001;
                    sign_qin_00133_00001  <=  0;
                end else begin
                    conv_qin_00133_00001  <=  ~tout_00133_00001 + 1;
                    sign_qin_00133_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00133 == conv_Sgntin_row_00133_00002 ) begin
                    conv_qin_00133_00002  <= tout_00133_00002;
                    sign_qin_00133_00002  <=  0;
                end else begin
                    conv_qin_00133_00002  <=  ~tout_00133_00002 + 1;
                    sign_qin_00133_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00133 == conv_Sgntin_row_00133_00003 ) begin
                    conv_qin_00133_00003  <= tout_00133_00003;
                    sign_qin_00133_00003  <=  0;
                end else begin
                    conv_qin_00133_00003  <=  ~tout_00133_00003 + 1;
                    sign_qin_00133_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00134 == conv_Sgntin_row_00134_00000 ) begin
                    conv_qin_00134_00000  <= tout_00134_00000;
                    sign_qin_00134_00000  <=  0;
                end else begin
                    conv_qin_00134_00000  <=  ~tout_00134_00000 + 1;
                    sign_qin_00134_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00134 == conv_Sgntin_row_00134_00001 ) begin
                    conv_qin_00134_00001  <= tout_00134_00001;
                    sign_qin_00134_00001  <=  0;
                end else begin
                    conv_qin_00134_00001  <=  ~tout_00134_00001 + 1;
                    sign_qin_00134_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00134 == conv_Sgntin_row_00134_00002 ) begin
                    conv_qin_00134_00002  <= tout_00134_00002;
                    sign_qin_00134_00002  <=  0;
                end else begin
                    conv_qin_00134_00002  <=  ~tout_00134_00002 + 1;
                    sign_qin_00134_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00134 == conv_Sgntin_row_00134_00003 ) begin
                    conv_qin_00134_00003  <= tout_00134_00003;
                    sign_qin_00134_00003  <=  0;
                end else begin
                    conv_qin_00134_00003  <=  ~tout_00134_00003 + 1;
                    sign_qin_00134_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00135 == conv_Sgntin_row_00135_00000 ) begin
                    conv_qin_00135_00000  <= tout_00135_00000;
                    sign_qin_00135_00000  <=  0;
                end else begin
                    conv_qin_00135_00000  <=  ~tout_00135_00000 + 1;
                    sign_qin_00135_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00135 == conv_Sgntin_row_00135_00001 ) begin
                    conv_qin_00135_00001  <= tout_00135_00001;
                    sign_qin_00135_00001  <=  0;
                end else begin
                    conv_qin_00135_00001  <=  ~tout_00135_00001 + 1;
                    sign_qin_00135_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00135 == conv_Sgntin_row_00135_00002 ) begin
                    conv_qin_00135_00002  <= tout_00135_00002;
                    sign_qin_00135_00002  <=  0;
                end else begin
                    conv_qin_00135_00002  <=  ~tout_00135_00002 + 1;
                    sign_qin_00135_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00135 == conv_Sgntin_row_00135_00003 ) begin
                    conv_qin_00135_00003  <= tout_00135_00003;
                    sign_qin_00135_00003  <=  0;
                end else begin
                    conv_qin_00135_00003  <=  ~tout_00135_00003 + 1;
                    sign_qin_00135_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00136 == conv_Sgntin_row_00136_00000 ) begin
                    conv_qin_00136_00000  <= tout_00136_00000;
                    sign_qin_00136_00000  <=  0;
                end else begin
                    conv_qin_00136_00000  <=  ~tout_00136_00000 + 1;
                    sign_qin_00136_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00136 == conv_Sgntin_row_00136_00001 ) begin
                    conv_qin_00136_00001  <= tout_00136_00001;
                    sign_qin_00136_00001  <=  0;
                end else begin
                    conv_qin_00136_00001  <=  ~tout_00136_00001 + 1;
                    sign_qin_00136_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00136 == conv_Sgntin_row_00136_00002 ) begin
                    conv_qin_00136_00002  <= tout_00136_00002;
                    sign_qin_00136_00002  <=  0;
                end else begin
                    conv_qin_00136_00002  <=  ~tout_00136_00002 + 1;
                    sign_qin_00136_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00136 == conv_Sgntin_row_00136_00003 ) begin
                    conv_qin_00136_00003  <= tout_00136_00003;
                    sign_qin_00136_00003  <=  0;
                end else begin
                    conv_qin_00136_00003  <=  ~tout_00136_00003 + 1;
                    sign_qin_00136_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00137 == conv_Sgntin_row_00137_00000 ) begin
                    conv_qin_00137_00000  <= tout_00137_00000;
                    sign_qin_00137_00000  <=  0;
                end else begin
                    conv_qin_00137_00000  <=  ~tout_00137_00000 + 1;
                    sign_qin_00137_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00137 == conv_Sgntin_row_00137_00001 ) begin
                    conv_qin_00137_00001  <= tout_00137_00001;
                    sign_qin_00137_00001  <=  0;
                end else begin
                    conv_qin_00137_00001  <=  ~tout_00137_00001 + 1;
                    sign_qin_00137_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00137 == conv_Sgntin_row_00137_00002 ) begin
                    conv_qin_00137_00002  <= tout_00137_00002;
                    sign_qin_00137_00002  <=  0;
                end else begin
                    conv_qin_00137_00002  <=  ~tout_00137_00002 + 1;
                    sign_qin_00137_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00137 == conv_Sgntin_row_00137_00003 ) begin
                    conv_qin_00137_00003  <= tout_00137_00003;
                    sign_qin_00137_00003  <=  0;
                end else begin
                    conv_qin_00137_00003  <=  ~tout_00137_00003 + 1;
                    sign_qin_00137_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00138 == conv_Sgntin_row_00138_00000 ) begin
                    conv_qin_00138_00000  <= tout_00138_00000;
                    sign_qin_00138_00000  <=  0;
                end else begin
                    conv_qin_00138_00000  <=  ~tout_00138_00000 + 1;
                    sign_qin_00138_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00138 == conv_Sgntin_row_00138_00001 ) begin
                    conv_qin_00138_00001  <= tout_00138_00001;
                    sign_qin_00138_00001  <=  0;
                end else begin
                    conv_qin_00138_00001  <=  ~tout_00138_00001 + 1;
                    sign_qin_00138_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00138 == conv_Sgntin_row_00138_00002 ) begin
                    conv_qin_00138_00002  <= tout_00138_00002;
                    sign_qin_00138_00002  <=  0;
                end else begin
                    conv_qin_00138_00002  <=  ~tout_00138_00002 + 1;
                    sign_qin_00138_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00138 == conv_Sgntin_row_00138_00003 ) begin
                    conv_qin_00138_00003  <= tout_00138_00003;
                    sign_qin_00138_00003  <=  0;
                end else begin
                    conv_qin_00138_00003  <=  ~tout_00138_00003 + 1;
                    sign_qin_00138_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00139 == conv_Sgntin_row_00139_00000 ) begin
                    conv_qin_00139_00000  <= tout_00139_00000;
                    sign_qin_00139_00000  <=  0;
                end else begin
                    conv_qin_00139_00000  <=  ~tout_00139_00000 + 1;
                    sign_qin_00139_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00139 == conv_Sgntin_row_00139_00001 ) begin
                    conv_qin_00139_00001  <= tout_00139_00001;
                    sign_qin_00139_00001  <=  0;
                end else begin
                    conv_qin_00139_00001  <=  ~tout_00139_00001 + 1;
                    sign_qin_00139_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00139 == conv_Sgntin_row_00139_00002 ) begin
                    conv_qin_00139_00002  <= tout_00139_00002;
                    sign_qin_00139_00002  <=  0;
                end else begin
                    conv_qin_00139_00002  <=  ~tout_00139_00002 + 1;
                    sign_qin_00139_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00139 == conv_Sgntin_row_00139_00003 ) begin
                    conv_qin_00139_00003  <= tout_00139_00003;
                    sign_qin_00139_00003  <=  0;
                end else begin
                    conv_qin_00139_00003  <=  ~tout_00139_00003 + 1;
                    sign_qin_00139_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00140 == conv_Sgntin_row_00140_00000 ) begin
                    conv_qin_00140_00000  <= tout_00140_00000;
                    sign_qin_00140_00000  <=  0;
                end else begin
                    conv_qin_00140_00000  <=  ~tout_00140_00000 + 1;
                    sign_qin_00140_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00140 == conv_Sgntin_row_00140_00001 ) begin
                    conv_qin_00140_00001  <= tout_00140_00001;
                    sign_qin_00140_00001  <=  0;
                end else begin
                    conv_qin_00140_00001  <=  ~tout_00140_00001 + 1;
                    sign_qin_00140_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00140 == conv_Sgntin_row_00140_00002 ) begin
                    conv_qin_00140_00002  <= tout_00140_00002;
                    sign_qin_00140_00002  <=  0;
                end else begin
                    conv_qin_00140_00002  <=  ~tout_00140_00002 + 1;
                    sign_qin_00140_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00140 == conv_Sgntin_row_00140_00003 ) begin
                    conv_qin_00140_00003  <= tout_00140_00003;
                    sign_qin_00140_00003  <=  0;
                end else begin
                    conv_qin_00140_00003  <=  ~tout_00140_00003 + 1;
                    sign_qin_00140_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00141 == conv_Sgntin_row_00141_00000 ) begin
                    conv_qin_00141_00000  <= tout_00141_00000;
                    sign_qin_00141_00000  <=  0;
                end else begin
                    conv_qin_00141_00000  <=  ~tout_00141_00000 + 1;
                    sign_qin_00141_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00141 == conv_Sgntin_row_00141_00001 ) begin
                    conv_qin_00141_00001  <= tout_00141_00001;
                    sign_qin_00141_00001  <=  0;
                end else begin
                    conv_qin_00141_00001  <=  ~tout_00141_00001 + 1;
                    sign_qin_00141_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00141 == conv_Sgntin_row_00141_00002 ) begin
                    conv_qin_00141_00002  <= tout_00141_00002;
                    sign_qin_00141_00002  <=  0;
                end else begin
                    conv_qin_00141_00002  <=  ~tout_00141_00002 + 1;
                    sign_qin_00141_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00141 == conv_Sgntin_row_00141_00003 ) begin
                    conv_qin_00141_00003  <= tout_00141_00003;
                    sign_qin_00141_00003  <=  0;
                end else begin
                    conv_qin_00141_00003  <=  ~tout_00141_00003 + 1;
                    sign_qin_00141_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00142 == conv_Sgntin_row_00142_00000 ) begin
                    conv_qin_00142_00000  <= tout_00142_00000;
                    sign_qin_00142_00000  <=  0;
                end else begin
                    conv_qin_00142_00000  <=  ~tout_00142_00000 + 1;
                    sign_qin_00142_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00142 == conv_Sgntin_row_00142_00001 ) begin
                    conv_qin_00142_00001  <= tout_00142_00001;
                    sign_qin_00142_00001  <=  0;
                end else begin
                    conv_qin_00142_00001  <=  ~tout_00142_00001 + 1;
                    sign_qin_00142_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00142 == conv_Sgntin_row_00142_00002 ) begin
                    conv_qin_00142_00002  <= tout_00142_00002;
                    sign_qin_00142_00002  <=  0;
                end else begin
                    conv_qin_00142_00002  <=  ~tout_00142_00002 + 1;
                    sign_qin_00142_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00142 == conv_Sgntin_row_00142_00003 ) begin
                    conv_qin_00142_00003  <= tout_00142_00003;
                    sign_qin_00142_00003  <=  0;
                end else begin
                    conv_qin_00142_00003  <=  ~tout_00142_00003 + 1;
                    sign_qin_00142_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00143 == conv_Sgntin_row_00143_00000 ) begin
                    conv_qin_00143_00000  <= tout_00143_00000;
                    sign_qin_00143_00000  <=  0;
                end else begin
                    conv_qin_00143_00000  <=  ~tout_00143_00000 + 1;
                    sign_qin_00143_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00143 == conv_Sgntin_row_00143_00001 ) begin
                    conv_qin_00143_00001  <= tout_00143_00001;
                    sign_qin_00143_00001  <=  0;
                end else begin
                    conv_qin_00143_00001  <=  ~tout_00143_00001 + 1;
                    sign_qin_00143_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00143 == conv_Sgntin_row_00143_00002 ) begin
                    conv_qin_00143_00002  <= tout_00143_00002;
                    sign_qin_00143_00002  <=  0;
                end else begin
                    conv_qin_00143_00002  <=  ~tout_00143_00002 + 1;
                    sign_qin_00143_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00143 == conv_Sgntin_row_00143_00003 ) begin
                    conv_qin_00143_00003  <= tout_00143_00003;
                    sign_qin_00143_00003  <=  0;
                end else begin
                    conv_qin_00143_00003  <=  ~tout_00143_00003 + 1;
                    sign_qin_00143_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00144 == conv_Sgntin_row_00144_00000 ) begin
                    conv_qin_00144_00000  <= tout_00144_00000;
                    sign_qin_00144_00000  <=  0;
                end else begin
                    conv_qin_00144_00000  <=  ~tout_00144_00000 + 1;
                    sign_qin_00144_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00144 == conv_Sgntin_row_00144_00001 ) begin
                    conv_qin_00144_00001  <= tout_00144_00001;
                    sign_qin_00144_00001  <=  0;
                end else begin
                    conv_qin_00144_00001  <=  ~tout_00144_00001 + 1;
                    sign_qin_00144_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00144 == conv_Sgntin_row_00144_00002 ) begin
                    conv_qin_00144_00002  <= tout_00144_00002;
                    sign_qin_00144_00002  <=  0;
                end else begin
                    conv_qin_00144_00002  <=  ~tout_00144_00002 + 1;
                    sign_qin_00144_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00144 == conv_Sgntin_row_00144_00003 ) begin
                    conv_qin_00144_00003  <= tout_00144_00003;
                    sign_qin_00144_00003  <=  0;
                end else begin
                    conv_qin_00144_00003  <=  ~tout_00144_00003 + 1;
                    sign_qin_00144_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00145 == conv_Sgntin_row_00145_00000 ) begin
                    conv_qin_00145_00000  <= tout_00145_00000;
                    sign_qin_00145_00000  <=  0;
                end else begin
                    conv_qin_00145_00000  <=  ~tout_00145_00000 + 1;
                    sign_qin_00145_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00145 == conv_Sgntin_row_00145_00001 ) begin
                    conv_qin_00145_00001  <= tout_00145_00001;
                    sign_qin_00145_00001  <=  0;
                end else begin
                    conv_qin_00145_00001  <=  ~tout_00145_00001 + 1;
                    sign_qin_00145_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00145 == conv_Sgntin_row_00145_00002 ) begin
                    conv_qin_00145_00002  <= tout_00145_00002;
                    sign_qin_00145_00002  <=  0;
                end else begin
                    conv_qin_00145_00002  <=  ~tout_00145_00002 + 1;
                    sign_qin_00145_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00145 == conv_Sgntin_row_00145_00003 ) begin
                    conv_qin_00145_00003  <= tout_00145_00003;
                    sign_qin_00145_00003  <=  0;
                end else begin
                    conv_qin_00145_00003  <=  ~tout_00145_00003 + 1;
                    sign_qin_00145_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00146 == conv_Sgntin_row_00146_00000 ) begin
                    conv_qin_00146_00000  <= tout_00146_00000;
                    sign_qin_00146_00000  <=  0;
                end else begin
                    conv_qin_00146_00000  <=  ~tout_00146_00000 + 1;
                    sign_qin_00146_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00146 == conv_Sgntin_row_00146_00001 ) begin
                    conv_qin_00146_00001  <= tout_00146_00001;
                    sign_qin_00146_00001  <=  0;
                end else begin
                    conv_qin_00146_00001  <=  ~tout_00146_00001 + 1;
                    sign_qin_00146_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00146 == conv_Sgntin_row_00146_00002 ) begin
                    conv_qin_00146_00002  <= tout_00146_00002;
                    sign_qin_00146_00002  <=  0;
                end else begin
                    conv_qin_00146_00002  <=  ~tout_00146_00002 + 1;
                    sign_qin_00146_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00146 == conv_Sgntin_row_00146_00003 ) begin
                    conv_qin_00146_00003  <= tout_00146_00003;
                    sign_qin_00146_00003  <=  0;
                end else begin
                    conv_qin_00146_00003  <=  ~tout_00146_00003 + 1;
                    sign_qin_00146_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00147 == conv_Sgntin_row_00147_00000 ) begin
                    conv_qin_00147_00000  <= tout_00147_00000;
                    sign_qin_00147_00000  <=  0;
                end else begin
                    conv_qin_00147_00000  <=  ~tout_00147_00000 + 1;
                    sign_qin_00147_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00147 == conv_Sgntin_row_00147_00001 ) begin
                    conv_qin_00147_00001  <= tout_00147_00001;
                    sign_qin_00147_00001  <=  0;
                end else begin
                    conv_qin_00147_00001  <=  ~tout_00147_00001 + 1;
                    sign_qin_00147_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00147 == conv_Sgntin_row_00147_00002 ) begin
                    conv_qin_00147_00002  <= tout_00147_00002;
                    sign_qin_00147_00002  <=  0;
                end else begin
                    conv_qin_00147_00002  <=  ~tout_00147_00002 + 1;
                    sign_qin_00147_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00147 == conv_Sgntin_row_00147_00003 ) begin
                    conv_qin_00147_00003  <= tout_00147_00003;
                    sign_qin_00147_00003  <=  0;
                end else begin
                    conv_qin_00147_00003  <=  ~tout_00147_00003 + 1;
                    sign_qin_00147_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00148 == conv_Sgntin_row_00148_00000 ) begin
                    conv_qin_00148_00000  <= tout_00148_00000;
                    sign_qin_00148_00000  <=  0;
                end else begin
                    conv_qin_00148_00000  <=  ~tout_00148_00000 + 1;
                    sign_qin_00148_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00148 == conv_Sgntin_row_00148_00001 ) begin
                    conv_qin_00148_00001  <= tout_00148_00001;
                    sign_qin_00148_00001  <=  0;
                end else begin
                    conv_qin_00148_00001  <=  ~tout_00148_00001 + 1;
                    sign_qin_00148_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00148 == conv_Sgntin_row_00148_00002 ) begin
                    conv_qin_00148_00002  <= tout_00148_00002;
                    sign_qin_00148_00002  <=  0;
                end else begin
                    conv_qin_00148_00002  <=  ~tout_00148_00002 + 1;
                    sign_qin_00148_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00149 == conv_Sgntin_row_00149_00000 ) begin
                    conv_qin_00149_00000  <= tout_00149_00000;
                    sign_qin_00149_00000  <=  0;
                end else begin
                    conv_qin_00149_00000  <=  ~tout_00149_00000 + 1;
                    sign_qin_00149_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00149 == conv_Sgntin_row_00149_00001 ) begin
                    conv_qin_00149_00001  <= tout_00149_00001;
                    sign_qin_00149_00001  <=  0;
                end else begin
                    conv_qin_00149_00001  <=  ~tout_00149_00001 + 1;
                    sign_qin_00149_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00149 == conv_Sgntin_row_00149_00002 ) begin
                    conv_qin_00149_00002  <= tout_00149_00002;
                    sign_qin_00149_00002  <=  0;
                end else begin
                    conv_qin_00149_00002  <=  ~tout_00149_00002 + 1;
                    sign_qin_00149_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00150 == conv_Sgntin_row_00150_00000 ) begin
                    conv_qin_00150_00000  <= tout_00150_00000;
                    sign_qin_00150_00000  <=  0;
                end else begin
                    conv_qin_00150_00000  <=  ~tout_00150_00000 + 1;
                    sign_qin_00150_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00150 == conv_Sgntin_row_00150_00001 ) begin
                    conv_qin_00150_00001  <= tout_00150_00001;
                    sign_qin_00150_00001  <=  0;
                end else begin
                    conv_qin_00150_00001  <=  ~tout_00150_00001 + 1;
                    sign_qin_00150_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00150 == conv_Sgntin_row_00150_00002 ) begin
                    conv_qin_00150_00002  <= tout_00150_00002;
                    sign_qin_00150_00002  <=  0;
                end else begin
                    conv_qin_00150_00002  <=  ~tout_00150_00002 + 1;
                    sign_qin_00150_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00151 == conv_Sgntin_row_00151_00000 ) begin
                    conv_qin_00151_00000  <= tout_00151_00000;
                    sign_qin_00151_00000  <=  0;
                end else begin
                    conv_qin_00151_00000  <=  ~tout_00151_00000 + 1;
                    sign_qin_00151_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00151 == conv_Sgntin_row_00151_00001 ) begin
                    conv_qin_00151_00001  <= tout_00151_00001;
                    sign_qin_00151_00001  <=  0;
                end else begin
                    conv_qin_00151_00001  <=  ~tout_00151_00001 + 1;
                    sign_qin_00151_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00151 == conv_Sgntin_row_00151_00002 ) begin
                    conv_qin_00151_00002  <= tout_00151_00002;
                    sign_qin_00151_00002  <=  0;
                end else begin
                    conv_qin_00151_00002  <=  ~tout_00151_00002 + 1;
                    sign_qin_00151_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00152 == conv_Sgntin_row_00152_00000 ) begin
                    conv_qin_00152_00000  <= tout_00152_00000;
                    sign_qin_00152_00000  <=  0;
                end else begin
                    conv_qin_00152_00000  <=  ~tout_00152_00000 + 1;
                    sign_qin_00152_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00152 == conv_Sgntin_row_00152_00001 ) begin
                    conv_qin_00152_00001  <= tout_00152_00001;
                    sign_qin_00152_00001  <=  0;
                end else begin
                    conv_qin_00152_00001  <=  ~tout_00152_00001 + 1;
                    sign_qin_00152_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00152 == conv_Sgntin_row_00152_00002 ) begin
                    conv_qin_00152_00002  <= tout_00152_00002;
                    sign_qin_00152_00002  <=  0;
                end else begin
                    conv_qin_00152_00002  <=  ~tout_00152_00002 + 1;
                    sign_qin_00152_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00152 == conv_Sgntin_row_00152_00003 ) begin
                    conv_qin_00152_00003  <= tout_00152_00003;
                    sign_qin_00152_00003  <=  0;
                end else begin
                    conv_qin_00152_00003  <=  ~tout_00152_00003 + 1;
                    sign_qin_00152_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00153 == conv_Sgntin_row_00153_00000 ) begin
                    conv_qin_00153_00000  <= tout_00153_00000;
                    sign_qin_00153_00000  <=  0;
                end else begin
                    conv_qin_00153_00000  <=  ~tout_00153_00000 + 1;
                    sign_qin_00153_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00153 == conv_Sgntin_row_00153_00001 ) begin
                    conv_qin_00153_00001  <= tout_00153_00001;
                    sign_qin_00153_00001  <=  0;
                end else begin
                    conv_qin_00153_00001  <=  ~tout_00153_00001 + 1;
                    sign_qin_00153_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00153 == conv_Sgntin_row_00153_00002 ) begin
                    conv_qin_00153_00002  <= tout_00153_00002;
                    sign_qin_00153_00002  <=  0;
                end else begin
                    conv_qin_00153_00002  <=  ~tout_00153_00002 + 1;
                    sign_qin_00153_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00153 == conv_Sgntin_row_00153_00003 ) begin
                    conv_qin_00153_00003  <= tout_00153_00003;
                    sign_qin_00153_00003  <=  0;
                end else begin
                    conv_qin_00153_00003  <=  ~tout_00153_00003 + 1;
                    sign_qin_00153_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00154 == conv_Sgntin_row_00154_00000 ) begin
                    conv_qin_00154_00000  <= tout_00154_00000;
                    sign_qin_00154_00000  <=  0;
                end else begin
                    conv_qin_00154_00000  <=  ~tout_00154_00000 + 1;
                    sign_qin_00154_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00154 == conv_Sgntin_row_00154_00001 ) begin
                    conv_qin_00154_00001  <= tout_00154_00001;
                    sign_qin_00154_00001  <=  0;
                end else begin
                    conv_qin_00154_00001  <=  ~tout_00154_00001 + 1;
                    sign_qin_00154_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00154 == conv_Sgntin_row_00154_00002 ) begin
                    conv_qin_00154_00002  <= tout_00154_00002;
                    sign_qin_00154_00002  <=  0;
                end else begin
                    conv_qin_00154_00002  <=  ~tout_00154_00002 + 1;
                    sign_qin_00154_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00154 == conv_Sgntin_row_00154_00003 ) begin
                    conv_qin_00154_00003  <= tout_00154_00003;
                    sign_qin_00154_00003  <=  0;
                end else begin
                    conv_qin_00154_00003  <=  ~tout_00154_00003 + 1;
                    sign_qin_00154_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00155 == conv_Sgntin_row_00155_00000 ) begin
                    conv_qin_00155_00000  <= tout_00155_00000;
                    sign_qin_00155_00000  <=  0;
                end else begin
                    conv_qin_00155_00000  <=  ~tout_00155_00000 + 1;
                    sign_qin_00155_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00155 == conv_Sgntin_row_00155_00001 ) begin
                    conv_qin_00155_00001  <= tout_00155_00001;
                    sign_qin_00155_00001  <=  0;
                end else begin
                    conv_qin_00155_00001  <=  ~tout_00155_00001 + 1;
                    sign_qin_00155_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00155 == conv_Sgntin_row_00155_00002 ) begin
                    conv_qin_00155_00002  <= tout_00155_00002;
                    sign_qin_00155_00002  <=  0;
                end else begin
                    conv_qin_00155_00002  <=  ~tout_00155_00002 + 1;
                    sign_qin_00155_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00155 == conv_Sgntin_row_00155_00003 ) begin
                    conv_qin_00155_00003  <= tout_00155_00003;
                    sign_qin_00155_00003  <=  0;
                end else begin
                    conv_qin_00155_00003  <=  ~tout_00155_00003 + 1;
                    sign_qin_00155_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00156 == conv_Sgntin_row_00156_00000 ) begin
                    conv_qin_00156_00000  <= tout_00156_00000;
                    sign_qin_00156_00000  <=  0;
                end else begin
                    conv_qin_00156_00000  <=  ~tout_00156_00000 + 1;
                    sign_qin_00156_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00156 == conv_Sgntin_row_00156_00001 ) begin
                    conv_qin_00156_00001  <= tout_00156_00001;
                    sign_qin_00156_00001  <=  0;
                end else begin
                    conv_qin_00156_00001  <=  ~tout_00156_00001 + 1;
                    sign_qin_00156_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00156 == conv_Sgntin_row_00156_00002 ) begin
                    conv_qin_00156_00002  <= tout_00156_00002;
                    sign_qin_00156_00002  <=  0;
                end else begin
                    conv_qin_00156_00002  <=  ~tout_00156_00002 + 1;
                    sign_qin_00156_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00156 == conv_Sgntin_row_00156_00003 ) begin
                    conv_qin_00156_00003  <= tout_00156_00003;
                    sign_qin_00156_00003  <=  0;
                end else begin
                    conv_qin_00156_00003  <=  ~tout_00156_00003 + 1;
                    sign_qin_00156_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00157 == conv_Sgntin_row_00157_00000 ) begin
                    conv_qin_00157_00000  <= tout_00157_00000;
                    sign_qin_00157_00000  <=  0;
                end else begin
                    conv_qin_00157_00000  <=  ~tout_00157_00000 + 1;
                    sign_qin_00157_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00157 == conv_Sgntin_row_00157_00001 ) begin
                    conv_qin_00157_00001  <= tout_00157_00001;
                    sign_qin_00157_00001  <=  0;
                end else begin
                    conv_qin_00157_00001  <=  ~tout_00157_00001 + 1;
                    sign_qin_00157_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00157 == conv_Sgntin_row_00157_00002 ) begin
                    conv_qin_00157_00002  <= tout_00157_00002;
                    sign_qin_00157_00002  <=  0;
                end else begin
                    conv_qin_00157_00002  <=  ~tout_00157_00002 + 1;
                    sign_qin_00157_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00157 == conv_Sgntin_row_00157_00003 ) begin
                    conv_qin_00157_00003  <= tout_00157_00003;
                    sign_qin_00157_00003  <=  0;
                end else begin
                    conv_qin_00157_00003  <=  ~tout_00157_00003 + 1;
                    sign_qin_00157_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00158 == conv_Sgntin_row_00158_00000 ) begin
                    conv_qin_00158_00000  <= tout_00158_00000;
                    sign_qin_00158_00000  <=  0;
                end else begin
                    conv_qin_00158_00000  <=  ~tout_00158_00000 + 1;
                    sign_qin_00158_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00158 == conv_Sgntin_row_00158_00001 ) begin
                    conv_qin_00158_00001  <= tout_00158_00001;
                    sign_qin_00158_00001  <=  0;
                end else begin
                    conv_qin_00158_00001  <=  ~tout_00158_00001 + 1;
                    sign_qin_00158_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00158 == conv_Sgntin_row_00158_00002 ) begin
                    conv_qin_00158_00002  <= tout_00158_00002;
                    sign_qin_00158_00002  <=  0;
                end else begin
                    conv_qin_00158_00002  <=  ~tout_00158_00002 + 1;
                    sign_qin_00158_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00158 == conv_Sgntin_row_00158_00003 ) begin
                    conv_qin_00158_00003  <= tout_00158_00003;
                    sign_qin_00158_00003  <=  0;
                end else begin
                    conv_qin_00158_00003  <=  ~tout_00158_00003 + 1;
                    sign_qin_00158_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00159 == conv_Sgntin_row_00159_00000 ) begin
                    conv_qin_00159_00000  <= tout_00159_00000;
                    sign_qin_00159_00000  <=  0;
                end else begin
                    conv_qin_00159_00000  <=  ~tout_00159_00000 + 1;
                    sign_qin_00159_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00159 == conv_Sgntin_row_00159_00001 ) begin
                    conv_qin_00159_00001  <= tout_00159_00001;
                    sign_qin_00159_00001  <=  0;
                end else begin
                    conv_qin_00159_00001  <=  ~tout_00159_00001 + 1;
                    sign_qin_00159_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00159 == conv_Sgntin_row_00159_00002 ) begin
                    conv_qin_00159_00002  <= tout_00159_00002;
                    sign_qin_00159_00002  <=  0;
                end else begin
                    conv_qin_00159_00002  <=  ~tout_00159_00002 + 1;
                    sign_qin_00159_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00159 == conv_Sgntin_row_00159_00003 ) begin
                    conv_qin_00159_00003  <= tout_00159_00003;
                    sign_qin_00159_00003  <=  0;
                end else begin
                    conv_qin_00159_00003  <=  ~tout_00159_00003 + 1;
                    sign_qin_00159_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00160 == conv_Sgntin_row_00160_00000 ) begin
                    conv_qin_00160_00000  <= tout_00160_00000;
                    sign_qin_00160_00000  <=  0;
                end else begin
                    conv_qin_00160_00000  <=  ~tout_00160_00000 + 1;
                    sign_qin_00160_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00160 == conv_Sgntin_row_00160_00001 ) begin
                    conv_qin_00160_00001  <= tout_00160_00001;
                    sign_qin_00160_00001  <=  0;
                end else begin
                    conv_qin_00160_00001  <=  ~tout_00160_00001 + 1;
                    sign_qin_00160_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00160 == conv_Sgntin_row_00160_00002 ) begin
                    conv_qin_00160_00002  <= tout_00160_00002;
                    sign_qin_00160_00002  <=  0;
                end else begin
                    conv_qin_00160_00002  <=  ~tout_00160_00002 + 1;
                    sign_qin_00160_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00160 == conv_Sgntin_row_00160_00003 ) begin
                    conv_qin_00160_00003  <= tout_00160_00003;
                    sign_qin_00160_00003  <=  0;
                end else begin
                    conv_qin_00160_00003  <=  ~tout_00160_00003 + 1;
                    sign_qin_00160_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00161 == conv_Sgntin_row_00161_00000 ) begin
                    conv_qin_00161_00000  <= tout_00161_00000;
                    sign_qin_00161_00000  <=  0;
                end else begin
                    conv_qin_00161_00000  <=  ~tout_00161_00000 + 1;
                    sign_qin_00161_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00161 == conv_Sgntin_row_00161_00001 ) begin
                    conv_qin_00161_00001  <= tout_00161_00001;
                    sign_qin_00161_00001  <=  0;
                end else begin
                    conv_qin_00161_00001  <=  ~tout_00161_00001 + 1;
                    sign_qin_00161_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00161 == conv_Sgntin_row_00161_00002 ) begin
                    conv_qin_00161_00002  <= tout_00161_00002;
                    sign_qin_00161_00002  <=  0;
                end else begin
                    conv_qin_00161_00002  <=  ~tout_00161_00002 + 1;
                    sign_qin_00161_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00161 == conv_Sgntin_row_00161_00003 ) begin
                    conv_qin_00161_00003  <= tout_00161_00003;
                    sign_qin_00161_00003  <=  0;
                end else begin
                    conv_qin_00161_00003  <=  ~tout_00161_00003 + 1;
                    sign_qin_00161_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00162 == conv_Sgntin_row_00162_00000 ) begin
                    conv_qin_00162_00000  <= tout_00162_00000;
                    sign_qin_00162_00000  <=  0;
                end else begin
                    conv_qin_00162_00000  <=  ~tout_00162_00000 + 1;
                    sign_qin_00162_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00162 == conv_Sgntin_row_00162_00001 ) begin
                    conv_qin_00162_00001  <= tout_00162_00001;
                    sign_qin_00162_00001  <=  0;
                end else begin
                    conv_qin_00162_00001  <=  ~tout_00162_00001 + 1;
                    sign_qin_00162_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00162 == conv_Sgntin_row_00162_00002 ) begin
                    conv_qin_00162_00002  <= tout_00162_00002;
                    sign_qin_00162_00002  <=  0;
                end else begin
                    conv_qin_00162_00002  <=  ~tout_00162_00002 + 1;
                    sign_qin_00162_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00162 == conv_Sgntin_row_00162_00003 ) begin
                    conv_qin_00162_00003  <= tout_00162_00003;
                    sign_qin_00162_00003  <=  0;
                end else begin
                    conv_qin_00162_00003  <=  ~tout_00162_00003 + 1;
                    sign_qin_00162_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00163 == conv_Sgntin_row_00163_00000 ) begin
                    conv_qin_00163_00000  <= tout_00163_00000;
                    sign_qin_00163_00000  <=  0;
                end else begin
                    conv_qin_00163_00000  <=  ~tout_00163_00000 + 1;
                    sign_qin_00163_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00163 == conv_Sgntin_row_00163_00001 ) begin
                    conv_qin_00163_00001  <= tout_00163_00001;
                    sign_qin_00163_00001  <=  0;
                end else begin
                    conv_qin_00163_00001  <=  ~tout_00163_00001 + 1;
                    sign_qin_00163_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00163 == conv_Sgntin_row_00163_00002 ) begin
                    conv_qin_00163_00002  <= tout_00163_00002;
                    sign_qin_00163_00002  <=  0;
                end else begin
                    conv_qin_00163_00002  <=  ~tout_00163_00002 + 1;
                    sign_qin_00163_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00163 == conv_Sgntin_row_00163_00003 ) begin
                    conv_qin_00163_00003  <= tout_00163_00003;
                    sign_qin_00163_00003  <=  0;
                end else begin
                    conv_qin_00163_00003  <=  ~tout_00163_00003 + 1;
                    sign_qin_00163_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00164 == conv_Sgntin_row_00164_00000 ) begin
                    conv_qin_00164_00000  <= tout_00164_00000;
                    sign_qin_00164_00000  <=  0;
                end else begin
                    conv_qin_00164_00000  <=  ~tout_00164_00000 + 1;
                    sign_qin_00164_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00164 == conv_Sgntin_row_00164_00001 ) begin
                    conv_qin_00164_00001  <= tout_00164_00001;
                    sign_qin_00164_00001  <=  0;
                end else begin
                    conv_qin_00164_00001  <=  ~tout_00164_00001 + 1;
                    sign_qin_00164_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00164 == conv_Sgntin_row_00164_00002 ) begin
                    conv_qin_00164_00002  <= tout_00164_00002;
                    sign_qin_00164_00002  <=  0;
                end else begin
                    conv_qin_00164_00002  <=  ~tout_00164_00002 + 1;
                    sign_qin_00164_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00164 == conv_Sgntin_row_00164_00003 ) begin
                    conv_qin_00164_00003  <= tout_00164_00003;
                    sign_qin_00164_00003  <=  0;
                end else begin
                    conv_qin_00164_00003  <=  ~tout_00164_00003 + 1;
                    sign_qin_00164_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00165 == conv_Sgntin_row_00165_00000 ) begin
                    conv_qin_00165_00000  <= tout_00165_00000;
                    sign_qin_00165_00000  <=  0;
                end else begin
                    conv_qin_00165_00000  <=  ~tout_00165_00000 + 1;
                    sign_qin_00165_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00165 == conv_Sgntin_row_00165_00001 ) begin
                    conv_qin_00165_00001  <= tout_00165_00001;
                    sign_qin_00165_00001  <=  0;
                end else begin
                    conv_qin_00165_00001  <=  ~tout_00165_00001 + 1;
                    sign_qin_00165_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00165 == conv_Sgntin_row_00165_00002 ) begin
                    conv_qin_00165_00002  <= tout_00165_00002;
                    sign_qin_00165_00002  <=  0;
                end else begin
                    conv_qin_00165_00002  <=  ~tout_00165_00002 + 1;
                    sign_qin_00165_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00165 == conv_Sgntin_row_00165_00003 ) begin
                    conv_qin_00165_00003  <= tout_00165_00003;
                    sign_qin_00165_00003  <=  0;
                end else begin
                    conv_qin_00165_00003  <=  ~tout_00165_00003 + 1;
                    sign_qin_00165_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00166 == conv_Sgntin_row_00166_00000 ) begin
                    conv_qin_00166_00000  <= tout_00166_00000;
                    sign_qin_00166_00000  <=  0;
                end else begin
                    conv_qin_00166_00000  <=  ~tout_00166_00000 + 1;
                    sign_qin_00166_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00166 == conv_Sgntin_row_00166_00001 ) begin
                    conv_qin_00166_00001  <= tout_00166_00001;
                    sign_qin_00166_00001  <=  0;
                end else begin
                    conv_qin_00166_00001  <=  ~tout_00166_00001 + 1;
                    sign_qin_00166_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00166 == conv_Sgntin_row_00166_00002 ) begin
                    conv_qin_00166_00002  <= tout_00166_00002;
                    sign_qin_00166_00002  <=  0;
                end else begin
                    conv_qin_00166_00002  <=  ~tout_00166_00002 + 1;
                    sign_qin_00166_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00166 == conv_Sgntin_row_00166_00003 ) begin
                    conv_qin_00166_00003  <= tout_00166_00003;
                    sign_qin_00166_00003  <=  0;
                end else begin
                    conv_qin_00166_00003  <=  ~tout_00166_00003 + 1;
                    sign_qin_00166_00003  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00167 == conv_Sgntin_row_00167_00000 ) begin
                    conv_qin_00167_00000  <= tout_00167_00000;
                    sign_qin_00167_00000  <=  0;
                end else begin
                    conv_qin_00167_00000  <=  ~tout_00167_00000 + 1;
                    sign_qin_00167_00000  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00167 == conv_Sgntin_row_00167_00001 ) begin
                    conv_qin_00167_00001  <= tout_00167_00001;
                    sign_qin_00167_00001  <=  0;
                end else begin
                    conv_qin_00167_00001  <=  ~tout_00167_00001 + 1;
                    sign_qin_00167_00001  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00167 == conv_Sgntin_row_00167_00002 ) begin
                    conv_qin_00167_00002  <= tout_00167_00002;
                    sign_qin_00167_00002  <=  0;
                end else begin
                    conv_qin_00167_00002  <=  ~tout_00167_00002 + 1;
                    sign_qin_00167_00002  <=  1;
                end
             end
             if (start_d5) begin
                if (sgnprod_00167 == conv_Sgntin_row_00167_00003 ) begin
                    conv_qin_00167_00003  <= tout_00167_00003;
                    sign_qin_00167_00003  <=  0;
                end else begin
                    conv_qin_00167_00003  <=  ~tout_00167_00003 + 1;
                    sign_qin_00167_00003  <=  1;
                end
             end
       end
   end


   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
            sum0_00000                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic93835a022c46b7aa00a465c407d7da2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I92cb615e2c439914e72ce001256518e4  <= 1'b0;
            I2e30088bf29cedd7debc15b1e6ec4ada        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iad799775eb657f8973e6dfcf70a9875c  <= 1'b0;
            I38f512bfb84094d1e92a10a345d5505f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifb064c69c7110c014593149ae69c75fb  <= 1'b0;
            I1e878f00f056f637625cb013a93325a8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7f7b30f2acbb8e31f50b58096b738254  <= 1'b0;
            I25db27464b31fee41ccd7a3cfe4d403e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iefe4099ff7e457f6b9fefc83e176c1a0  <= 1'b0;
            I19417a224c5cdf1211e9790aa29c4c5c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icddb43f9b760a4597a0bb637fb405616  <= 1'b0;
            I16dcafa854ea9c67d8a080feb2ba9166        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic76e72b434b47c10ebac3fac4ea50bde  <= 1'b0;
            I7f63338eee2663fbe61fffd248433310        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9eb87e62d23bc87d7cd82c0f329f247f  <= 1'b0;
            Icb1e3c56c8729c32d43c69710e345db2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2eac5b39c6f485c9ae0bd341f894633d  <= 1'b0;
            I6ece8e3c1e89613879336936f77d732f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I76992221b1edff5684c482df7ac4693d  <= 1'b0;
            I72a646ae7e32a16af0f5930a6e95b36a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iada5bc4a51dc1bf57bb9cca11326bdff  <= 1'b0;
            I7e72d119dd93a6ab05a23fde0a865866        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I364ed3f83c49626bc3b939e53524d9c7  <= 1'b0;
            Ied4fdf5805039cd2fcd042fd13755fdc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic2b000c3b2ca3beff2d427caab04701a  <= 1'b0;
            Id44c2293b765cff450dd1d747c47c1f3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8e873fb2321eea82bb590a92411e2e2c  <= 1'b0;
            I8f4ed02f7aeb823b745040f7f3f43ac7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If4cb744ee52b6ae793431cd038069b57  <= 1'b0;
            I6488b9b8f405d7d81a4874fab2678102        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7741e239c16828889d488cc87647c154  <= 1'b0;
            Ifff612d16828ec907a348479e19ddf31        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7979161aa1e2262ebea862004c387697  <= 1'b0;
            I268262076f22bc6b1507bc8f91b98a0a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic62fc602da3d16fe13d03a49a21269d0  <= 1'b0;
            If1f732841adb7c0cad1ba37c0f5fd517        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I94009bb7239be96243902ab0f0abea7e  <= 1'b0;
            I0df8a24f31c027756d248c3bd1b9bf7b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iae7b72abf4d3c536330a229e3836b441  <= 1'b0;
            I8ef901e733b12e76412eb36684e2b575        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie5d9cc18b2dd300132470f206452ff17  <= 1'b0;
            Ia48916a02f68b1b8f5fc7fece04677bb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7c791c854d0bc28e8dd787545f8fbda0  <= 1'b0;
            sum0_00001                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia37409944d9fdd3b16e7007e13d82a79        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5b177dd5c14ad082516b47f550875682  <= 1'b0;
            Idd65f149afe9d5f63ddaf34b82b11e95        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I55e4ad2d71a29ad63b4999d64ac0dc4f  <= 1'b0;
            If2886d560854faed32ebd8e33d868973        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I59c5da6338f431a626c86a065a355c35  <= 1'b0;
            I77778118bb3ea900c080754ff4c49c26        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia098bbeda8b755ece6b88eac83d03e55  <= 1'b0;
            I7292ed752d8741594d757730950feea4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie7470dd75b54d14038de19e4d3043ba9  <= 1'b0;
            I68cfd7868e061793ee8a41e69e80219b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie95662d4faf6b5a4cd5ecfa41697b983  <= 1'b0;
            I667ead814b303fca64ef047bb8246b19        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia1b617e3d141263b51e58c5ef0bd7a89  <= 1'b0;
            I4f25c7edb12e868cb5532e42b4ba5133        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If9a5d830e3ade0fd96b98f5949f165f0  <= 1'b0;
            I5aed2d82717f359bb5ac5a0ab91b7beb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id3de87169c440f95d406693ef77cacd6  <= 1'b0;
            I92835fd54631deaefa7b214e2c4b9bff        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3751f191f5009322acb7c9be4f8d7129  <= 1'b0;
            I67e067da565635fcff166e3a7d0c446b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic1927bb3335f6a28c0816eba12d3975e  <= 1'b0;
            Ifdb0f307b1b9458c0487a1574ccc094b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia659126b51468cfef48c97a135a71500  <= 1'b0;
            I5c6b7d143e42fd3b8bcdb7d7ed4da2c2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3c3c22bf63e55a81ae91b1dd1ef615a0  <= 1'b0;
            Ie679a21d0136a08cc5e6526e9f8d1843        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia62832d325f86160285c4d1a790a32cb  <= 1'b0;
            I611942a72a5e12f6afaea6bde6699ef6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I83c7d177eec2dad0a924557cdc91ba77  <= 1'b0;
            Ica9883c97f823a4491cbee5b45c43590        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7050adb9d06f767549b7f35c4679e391  <= 1'b0;
            I8e6addfc61f5bfb7af74fc2993639565        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I04aacd95d9e44657f616e01c9053f0fb  <= 1'b0;
            I9d53619f10e2a426f7297bbf7c81158a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2ff317d57f59747c4524ef4278d51092  <= 1'b0;
            I8a055c27778913287ad951183fa0d4d6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8bd2a9d90074500698b302cb8db7f03a  <= 1'b0;
            I8f6ae5c80bb2f50084b5f5ee5ab0ffc3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3b8cdfb1440732ce98cd1676e05a2af1  <= 1'b0;
            I3db8b3a342e8e2f13a448246aa001c2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I671de3d408b5b783541663c7f1e3a6fa  <= 1'b0;
            Ibbee0996ea0f5e16b1f711345be7f2ae        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I446857735e680cae93a24dccb59b1924  <= 1'b0;
            sum0_00002                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Idb777f1eb4c3cbba103b9b43f948ccf9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I77b05a8aa92c66a235195a66dc13c0cc  <= 1'b0;
            Id5e46b1f8844c7587f99d22170581a24        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie92110d19f4886cdfcfacd0920c06a4e  <= 1'b0;
            I67aadabd3cf49456cace7392a1e7a35a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I36ba87b69b5b9dd919319230f697dfad  <= 1'b0;
            Id5635595d6b7b6dd7e6d510a27ad6702        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id20e72ac258d1d1b6cdca1e6c9e3596d  <= 1'b0;
            Ice783314a4868f0bba8bc3c5e3b65ae4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifc34f5d6b7a7d0533439794958959856  <= 1'b0;
            Ib2d9b7f58cf571b904be02e6073f9b94        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I849ee5d34760be03d4285185136aa52e  <= 1'b0;
            I61b6effae91ae4bdcce4550eb5cf0796        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia3559d98eb372b7307f30ad1f7c4c7cd  <= 1'b0;
            If5cf6e81b0e3b77f6a45f2555201acc2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7332e088bbff69db19c62685e033d26a  <= 1'b0;
            I62fae5bf51588f28c3521715b834909d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I44daa5992b00e7af19adbee70bf01f2b  <= 1'b0;
            If5cbdab78a4cf86b6285a400d0e0ac90        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie517386cb5832e406fefc5e85eb2e7d1  <= 1'b0;
            I6e481cc49441c08bcd9fdcabbe90a000        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9b096ce09467c10f448496fda13987d2  <= 1'b0;
            I3aa663be3dd604564ef68b9a2b9d7319        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If1c0a3726041f70e508d68cbf6e40e04  <= 1'b0;
            I8031632ee8700c63c207e2d6a6bdb630        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaf36ce8598a29573979c683a5e2cf9fd  <= 1'b0;
            If9be2701858da0bdffbf2dff7bcfd7e1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ice82cfe55a5f226746e59e5c8beb46be  <= 1'b0;
            Ief209532f4cbf1c6a41bea414577f825        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iea1297491d1dfe98f395d8c73808a893  <= 1'b0;
            I1c8953ad3f64f3c3cc506808aad29dab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If43dd31198c8a0da6fabd194cf13bb70  <= 1'b0;
            I1b519d88bbf86cfb080a50ea0480a128        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibeb8c72b90b50c6897224ca1a792fa56  <= 1'b0;
            I5b8258f35d889071109216b464abb2a4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8e87530a131b5a73cad6df68b9e4967f  <= 1'b0;
            Id9681d4e0e4d375f9279de115a4337a3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idf8d15c7bd7705b9aafbda09c3a5b46c  <= 1'b0;
            Ib42144ece00b82debd70011724a29c91        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2aea17846a53e2eb2968581ee2c48226  <= 1'b0;
            Ic5717058a1815f63f164de1b1defe8cb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I169d8f2bb5fde5b202b4239b7a7f1ed5  <= 1'b0;
            Iea41672f012f225d64d9c75b198c812f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I40a223380fb4414a3f26a08cb90025ec  <= 1'b0;
            sum0_00003                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I7a070bd014e1d2c5e55e5fcba88a5664        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie117f6ec475f5d6444998af151ce4e69  <= 1'b0;
            I4a0a8b28429b708363458c74230b0fc2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If7f3174da35dd39af7f4792aaa649bf1  <= 1'b0;
            If585e4075ac1740f3b141ae6a50200f7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I719a892ad54e63b217c7271741b29cc5  <= 1'b0;
            Ie1a68cf09bb21a1629369fde87f51bea        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4acf6d84471cd237f65c9b2391b7a20c  <= 1'b0;
            I72b8547125d0ad6c1ad39a68b55c818c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7a387a1f887c32e9d0f8e89912a8618c  <= 1'b0;
            Ie14ba4a8657740f9a8d057258db2cb09        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib862ac63c230ccde7fae0e62f9d047fe  <= 1'b0;
            I27490a69fb2a1f6f298639254c37cf9e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8f1a8a22637d37c3692e808d5eb3d543  <= 1'b0;
            I49b9c212fbe74a5dd8b087e417296186        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6f420c64640dfb0c001f57df7e3b4504  <= 1'b0;
            I0a8e6f5cc8b6ea599b7605abe6479bec        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3600031716c2b4e21c9f577d34e033dc  <= 1'b0;
            Ib6d94b34d3886717e4016fec196f277f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I002820a37fa7c6c504c487df4368e2cf  <= 1'b0;
            Id7e53d36da7171e036ebfc984dbcea6e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8a4c1f23212ff846400651b100add502  <= 1'b0;
            I2ec254d80fd0683d782302cf3839559b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ice1ce5b4c30841dd92268559ebadafcf  <= 1'b0;
            Ibbedaef61051d5df82cd6d55e05c80da        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3eeeb1949945032d6c1759875426b733  <= 1'b0;
            I501336bb7ba172c05dd5840036e6228c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I384d5377ee6b8f7eb2db23a2e444ddbc  <= 1'b0;
            I8e5c4c6c63e42054359cee697cc0d026        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I30d615203b697787ead37394953925cc  <= 1'b0;
            Id3daa6db921871b752bf92366446afcc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib16548d471f0a4f4625852ea04335dcc  <= 1'b0;
            Id8367ec60787bfad0da8aa76c6ed8ddb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0987c561670b7b2b6683303c1be39561  <= 1'b0;
            I533649312ec995f1f9e514c59a8675b1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2bdf4736022e5da7294a0e851006a124  <= 1'b0;
            I0621d0b2c83e70b4afd65eb9dca4b514        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic6fd9592d2ffcb8f4ca83c6f0bd19975  <= 1'b0;
            I2ae01892a3cd0432618d7280b31daddb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I14bf11ad80890227e47fda26ae1b9c24  <= 1'b0;
            I5ed8a2f30bd2ea269341c2267ae3fe83        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8ca17b6cf35e1b1f8f601604575d3f27  <= 1'b0;
            I2c819e7f62c0dc0aac650074b203163b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I275cd09649a750edb8ae8313e4e1e279  <= 1'b0;
            sum0_00004                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I30e20b58913d6fbe5817e1956ba8e570        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7d6a6026eb3c4d06e682523424f9628f  <= 1'b0;
            I1b922bed7f3c4a6705f3ce7a885a68cd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia0c192e590d8c914555b434ce5a634a8  <= 1'b0;
            I2f65f0917713ecc8585392d3b557c1bf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic98c8641d2022080297c54ff2539e75d  <= 1'b0;
            I3301533e7d9e527118a67c462f1b4357        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I87f34821cd0b58f8855b25c75f2dd32d  <= 1'b0;
            I52a88bdb1f03da82730f7579b7b5305d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I87211ac14d832ad3205d47fb83cf256a  <= 1'b0;
            I644c730662b3725d26cd46fb46106104        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib81431cfb3b281555fa7e5b4582a2524  <= 1'b0;
            I3da3e36c76c4123bec6879bccb39e933        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I835b902949c2c4c09b757d4d35574a76  <= 1'b0;
            Iebde55cddc8170f7dd8855ea55eff0ce        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8510240df7dc41f85ad58a39868a1fd7  <= 1'b0;
            Ie673e2d92a7090b2fa1c5e14a2e03be3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1b6abc8fbab3849b285e9f88a4fe867b  <= 1'b0;
            If90afe75714f8660ad0eb9f9ea06cd6b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied638fee34f8baed4154b0b72e43a21e  <= 1'b0;
            Ifd96e3a6e0050c30a4308328cfecb21f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I14fa7aebb608d4a3d67176ba27d34d9a  <= 1'b0;
            I68b92cc2d83e9a718edd2aea82314016        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iad90879acba3fc2101829549264960f3  <= 1'b0;
            I6bdbb92363f0e072ed04654e9aad17a5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ife0952b85f14a960007b67646b0cd969  <= 1'b0;
            I87a4267db59b97ef1b9bca8743cb0322        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If876ca6a14ffb4323503ed46666bc25f  <= 1'b0;
            I44eacb2bea725efab7c0dd560279f0f8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If2dfcbf493b761fb5d7c622e739b23f3  <= 1'b0;
            I87a2736466c5ee62b7cc55f17e715ffa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2c8f4a147b363d9c5ef0e080d9a9ed40  <= 1'b0;
            I7a66c7713ba126fdc24940cd92f7e10b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I485f9d1104a965d5d035feef912a2ca8  <= 1'b0;
            I1f11c579f34c41aade41c53f53468057        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I10fca5f2cbf5e2bc3433c0dda579a051  <= 1'b0;
            I651a438f70583d476ae10f066e035435        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If8572800d5d80cc92dd917b60447b63b  <= 1'b0;
            Ibdf17fa73794c846e15fe0a915b071e5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I24645082ef16129eed1c574f5fc601ca  <= 1'b0;
            I76d3221fbcefc0ee08655f7ba4919f3c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I207a0f6184a0b3be71766a8b47ea5535  <= 1'b0;
            I3458f69c90ea8b20b3d1f67e9a13ec2e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5cac08dabbb6de3b01c821d4db93a8e3  <= 1'b0;
            Ia2d6e9e1e92a30c7028af50ddfbb9bf9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibe6b8c57d7ff47b6fdad5fadf1f6b841  <= 1'b0;
            sum0_00005                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I66c91b5133d9812a03daecc0b14211f8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I477326720157df2503149125a43ee987  <= 1'b0;
            Ifb5986949e88167526d9fcfe07b417ca        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2c741a5fed7d88e9bdd6b7459feac649  <= 1'b0;
            Iedada801ca6cd173ee523ef335e91ff6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17a6511072c7fb4846be5844decf17d6  <= 1'b0;
            I4e2722e547586da7565b2d91a7fc91e7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5ebc3047985651f4b9a957d502a97e95  <= 1'b0;
            Ib321a8ceda62c64ab25dc1c718301bda        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifa09fc1b009d073d5a9973b430c63469  <= 1'b0;
            I58daeebec4873e6c1c07c090ff81235c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie6212a29c7c6b035cfff4c869f945b68  <= 1'b0;
            I3f103fbbe49c86c9db46129bd4632cab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If343015b4815b01dae88bbb6f2017b3d  <= 1'b0;
            Id6697ca17f1bd6ddd112951b9d89a8ea        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia0116a3cebf94318ed5b287960957ad6  <= 1'b0;
            I445ede2983c7470b4418a2ec0cbbd5e1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id75c23e80cdf25d883806ed20d4ae783  <= 1'b0;
            I034e56cd77ee400ed81b78177b202930        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1b43f29e0ddb72467befd6f3a9c1c829  <= 1'b0;
            I08edadbd9366786f96b44268d096b4aa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3fd0fa3b774d30a267d61e9427d09f3f  <= 1'b0;
            I8f86a7af86eb04c5df18e09888cdce7b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2eb08ebaa07a1004638cdd61a7209b7d  <= 1'b0;
            Ic00d037a11f8a27ab34e4daab8c9c2e6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I258c45897919cec5c6acaddee7f3a41b  <= 1'b0;
            I4d95ceccc6c3ad37f13c98339c59e5c4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib42d37576e3aff3d205f1f8822cc58b5  <= 1'b0;
            I1ea967d377f462a0e06d7d0d4d95b342        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1c2ee281cd47a8414851c5e1c758ea65  <= 1'b0;
            Ib0feec63123e66bd6ad6935e9b7fa6bf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie644d131c4f2c603e8e64c5581fdf822  <= 1'b0;
            I7d120060ddae9ff8f7206b3ef63eda50        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9b76f0121a3f7e887e7121db50024ab4  <= 1'b0;
            Ib47f8f72386e2e65a88fbadd3a705225        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9eaf4e9ebe07717503ff69b51f0e1905  <= 1'b0;
            I4e0efc35346e2934f5bb4c34a4bc5f90        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icb0841ecf142687c3aa23e68f01c927c  <= 1'b0;
            I3ca1014802f58087e3434a1e0df19c01        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie8c0fac00a9de74870e59cbf9e87a39b  <= 1'b0;
            I688a3879b7be1544e6f94b4221c03213        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iae5d6faac1f5685cb1d400ee2b1d85e0  <= 1'b0;
            Ic22988138610c8671ec342f65f34c7ae        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib62b02ddf0f57bee49838d19783ef6c3  <= 1'b0;
            I0b85fdd83569e5cbb7d71eed50cb32fd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibd59d0e5a062f149bd0e91ba76985a13  <= 1'b0;
            sum0_00006                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Idf55390c11e5b41ebc2a28e0af109913        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I876fdba97e755b74532f7ab191fbac14  <= 1'b0;
            I6b48935ea25672ee9a42f49eae9e519f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8edf1a08ef943f06ee28771c6e140e28  <= 1'b0;
            I6a9e6c39c20e45773dab7823a7ff9486        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7e12ad8a8ef857e02f4563b2f3a7f0ca  <= 1'b0;
            I42907182010c5889ddb7a700ead16525        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17b3a9df6752da6cc987e902e6bbad48  <= 1'b0;
            Ib6c26f3e3358cc2ed6fbda83eabd4bd3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I487496233a32f657171b3789590d0522  <= 1'b0;
            Ia50d85808790790450f87a5246874b3f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie34534dfd435b3d1cf35e82ca71e83ba  <= 1'b0;
            Id4a1744702d7808a80bc40697c864765        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0e8679271ba733bb87c44b6b9f0b6ed2  <= 1'b0;
            I0cf3d2f3e6793a2dcf15949da16ad28d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic14760b65c6fe150c3c48e64389a41d8  <= 1'b0;
            I90bd9107f4c931fa1ccb92998ea8cdeb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied6c684cdd280b41ffab93a026d27282  <= 1'b0;
            Ida1c729e6bfcec2c31a92aa9002f2c68        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id0f4dbb72da33748d8baf723c5a32567  <= 1'b0;
            Ib848feeccd0ea78ebc8ba8368534c3d1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib0bb71b1f8829347b3a9a7543f9dd964  <= 1'b0;
            Icc11970bbae3adcfa33a0e5dba3e78f4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I47cbb92d2284aef7b9e56e88f0ba6f7e  <= 1'b0;
            I86bb4ef4bdd7af8861280ef30fbeeeea        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic69094123b75ae36e3e54f179a9f2cb5  <= 1'b0;
            I7e0c259c6c7bacdff5edc44a22e005ba        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I07abbbd75d91018ac53f53e64cffafb9  <= 1'b0;
            I897ddba059b27f7ed009b0cb70cfb46f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib02268d5048c7c8e83118070e927453f  <= 1'b0;
            I4496243eb0542a514b551b4d09bffd7d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc2a9c6dd8d2aa912548c918c8a488f4  <= 1'b0;
            Ic931fb08b2e8441321ebdeed84576a0d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5ad7eb9d3ce7c712515254f892d1670d  <= 1'b0;
            Ieb6af5390b98e893ee05a939c16d2ffd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ife25829fb3c5023b7d69bbaadf9cf77e  <= 1'b0;
            Ic2a54bad4c5a8885dd24b8687c6db0de        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8b2a79aa4ac88e6b4ca8188a7852022e  <= 1'b0;
            I6ecbad763d2b48b78a0584beaefc78ee        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I081e2595b18f306a74d070203447ecf6  <= 1'b0;
            I20556d23c873c71c7ebc8a961bf40251        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I68b152a599887c0039dd9d45c528c219  <= 1'b0;
            I79012e6351e6320c22437aa216ea4df1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id051f1d5454802e0eb37e22248efe8ca  <= 1'b0;
            Ibf74ab9af877d27c3a6f3881f00ddaf1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic4c6f707f461cebbc4c93f2ba664ae7b  <= 1'b0;
            sum0_00007                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I843d35db35d7b42a87ce78d3772cec2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia538dadbd6ae3711740595a18c89b65d  <= 1'b0;
            I2b1398b4bfd374d7221b0a68da28e979        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie7d9730b191781c78391141d95d4f8bd  <= 1'b0;
            I6f615d6e74b0c02f8e4265523ad16404        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I12f2f886517647044cc251861721bbb9  <= 1'b0;
            Iae8a98dd4a7cbfbc56c1404b6a2020af        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I615053b36a1851a06125e2ed5ec7f880  <= 1'b0;
            Iad53375a54d01c559c74981bf279dfb5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifbc6aa14cd448bbe416897a3671ba857  <= 1'b0;
            I5db1307f922e0c742d7d9f3a79a4a4f3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie596289582a73e37f78f4ca4cab21e3c  <= 1'b0;
            I9f78172ed5bf73752196f9a8810005f3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifad8c7bacf72583f91be27fbe5b7a1e1  <= 1'b0;
            If85a22d670d47f491dd7568d0453ba1d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie74c72742807ae4243748fd27d80d626  <= 1'b0;
            Ib9e529170b2896e930a839295796fd31        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie7a68c2b368a295f95571bc4a109b9f1  <= 1'b0;
            Ib7af536846bac40c1f221d1f72c6c25c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id88a7edf897eea1b4a137141789a04f5  <= 1'b0;
            Ib0eb61a2cb831dd35ce9850994e7c2da        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib13436ad16a37d656d6b1ee95b9aee20  <= 1'b0;
            I89d338f59960af7a47595d6afa206abc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc07dc30c0a957e474546ac7a60df38f  <= 1'b0;
            Ib3c1176eb8991e3e85855a9fe845c303        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I595665d8128bb87ab62741d7ac520a4b  <= 1'b0;
            I93073d05d509b821a743998cf32c58ee        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I256050251d23250854ff337bef28e460  <= 1'b0;
            Iab6dac1909c1564c3890ffecc13418df        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I82f0e5a32d1bcd761a74f1f9ce8c88ba  <= 1'b0;
            I1b75eeb29167a171d89f6e67039436d5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I98febac90cccb5fc1f3d966b6e38c4d3  <= 1'b0;
            I3a31adc52a1405555017b2ddf219b407        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib534288c2cf976b6ec85db743bc2a823  <= 1'b0;
            Iaadba89c6a370240fc0758029f7d8db0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If988b82b86db1f4ff6d3695f7b0197e4  <= 1'b0;
            I4f4a64fb3ced7d9f7ee4513178e9655a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6ef260ef75e47b011a46ba2080ac3684  <= 1'b0;
            I0c76ca58f69c91758e755cd581241284        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifc1da524e7670772834d521a6fc4c96f  <= 1'b0;
            I2312bce18958346149c868846e04643b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I852d5295a32984af00c95f6d9389555e  <= 1'b0;
            I3e154098cb0a48f1c23234f46613f406        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3c0a621dbef864fd1f566bc2e47f32c6  <= 1'b0;
            I1645c1c588bcbf15dd62d47e08b8e139        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic04828ba2db8239b093043c27476d345  <= 1'b0;
            sum0_00008                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4c25de66590e1745d37112e08d8c8e2c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I319012bc6fe93d78de57bcace0caaef5  <= 1'b0;
            Ia03092ac621b8dd1c206fea1e8b0215f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibb35bace971548c9fc98d773d1aff712  <= 1'b0;
            I5c9bdb033436dc9f6069baca31f24c2d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I90023493600924a76d2192080cf6194e  <= 1'b0;
            I8f07cf4865480f18ad6945974ec2231c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia9f5ce4603af279bbd9b486b67016482  <= 1'b0;
            I4a7119e8862fe4a6a4100dd9ac67dd24        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I05721e06a1acdcc0571907c7d853f18c  <= 1'b0;
            Id78fcfc6724a05f46d44d7c3e7d0c756        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibfcfd3151af0d82bfce293ada44059b3  <= 1'b0;
            I7cbd9d619623cbabf8ed6b1fece8f012        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9539fcc40d26b13015a864718b116d5b  <= 1'b0;
            I58951165d251e370b0f3b3fb537aed18        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5490039998187a1a2efc3549e3dee7d6  <= 1'b0;
            I21daac106f526d84cb8fa5239c19499d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2b97a79c90f6578c8b2f321f8d598cc8  <= 1'b0;
            I178029cec3a5d6141abdfa91b91fdbf4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0c616f736879c28a5222de3d6f49a587  <= 1'b0;
            sum0_00009                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I96dfb2efbb55a644616e3474ed07c364        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5590d801fd7fb496019d4c31b7c6d898  <= 1'b0;
            I7a17d8f0e2d16c441044db68ee037731        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I27e1d2e0e980216b27b90ea48c061025  <= 1'b0;
            I2ced9bb3ae6bdc5b5ef2865fb46abf07        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I474f6bd977f4197742d0bddb3bece684  <= 1'b0;
            I89a93384020d93cf4d26b3902e06cd9e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaa1e981134f5a5c02983c49562683bc5  <= 1'b0;
            Ibbb47d29b9a45559c13ffa3b046c66f5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib051eb1091a85f85a1e50007f1b27cab  <= 1'b0;
            I0034177eb1049577a3578b371527f34b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6b5645cdde4b35a16fe3e91d90caaa4e  <= 1'b0;
            I22d9ea7bb5a1a3405bcd04b9af40fa62        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8850ab26807dcd55fefadf6310729ca7  <= 1'b0;
            I8a632e7a911bf5726fee587189cb6f16        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic5cb81c821716a8aabf8cc2283ff73ba  <= 1'b0;
            I3765afc490b34e8a310998a4ebcff8cb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9a6923c6368526a53ef70e16471386ef  <= 1'b0;
            I7607e800ae46a96e016b303120da4247        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I620b8ecdcaccc1ec80ebcf9fa6af0017  <= 1'b0;
            sum0_00010                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I29b2f1fddee5e32f217d25410bcfce4f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I141cda06bae0c5666e3bc61c6fe5ad66  <= 1'b0;
            Iba5f8a31a81f6aa06f5e38c03dc6db54        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia9c273b32d0701c7f185ab2de9e57829  <= 1'b0;
            Ifcb5c907ad503331317599e4e0ce7be8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic3fb524ab434e80b3289c9241b65d224  <= 1'b0;
            I62d6f2ab4ec8b6ecfa544ad4d90eb30b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I23c8b64e433af0bd00cef44e38df99f8  <= 1'b0;
            Ide65414c51b3cb182c0f2f238903d60a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If6a5dc79c0f6ce348956286737a369d8  <= 1'b0;
            I03a8dc2288eaeb619e746990e20cc868        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I34e6e9d2153e4a70ee36ab85e72d5318  <= 1'b0;
            Id81c1b44d16ddbcd466382c60fe84986        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifdabf743a8cb46b7053000ff48ea0c60  <= 1'b0;
            I503d72f4a2fd20dbf35aa27321d2ede7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I22f5bb821a2571d1764978fd76c8f1d0  <= 1'b0;
            Id6595a4cf33062d1f05cbcee2d0685f1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1b695aa715615662eff7065c742b0859  <= 1'b0;
            I83ebdd7331ca8fbcf5250851b346c0b0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iec91b3ca3b54010755d57f8b8ea4a544  <= 1'b0;
            sum0_00011                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I7f6ea26cdfe5986065e7b5aa6842cc1c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I06ad520cb02e46d34c45f207d42a9243  <= 1'b0;
            Idab1ec32c20f93c4cc1acb38158f92d5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9d18ff3465afd8cae63abba68487542e  <= 1'b0;
            I0738add83419502e73674ded2f1ad6c7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I914dedc1d5e5e21c9b8d07ec0ecc01f9  <= 1'b0;
            I6c93e63a8e5a2dbd598f1565c7323b39        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3375fff5ee0d4b4b12c5a70fbdee59fe  <= 1'b0;
            I4aa57a9d46371f1680d5f95596f60b5d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia8e304ca12c82e41cb8e4de7be199394  <= 1'b0;
            I5369a7203b78951a3c006c2d3b22507c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3566f2779e860008b1a5d305366a07c9  <= 1'b0;
            Ie72a79a6966cf198687b7c8a8bcdeb13        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie68b31360c12a83c6095254b6f14603c  <= 1'b0;
            Ie917ae4c44ab0f9c2f1747ff0d2a754e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I42ae0c42360c977b35429ce290516a6f  <= 1'b0;
            I0b1a31ccb34a742552c11b1945e23dd8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibe01835305315fab50269c72ef849b61  <= 1'b0;
            I9a65a845cf2eced39050e8481665f557        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id806a2df1c4519bbbe811791cb4072f9  <= 1'b0;
            sum0_00012                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I3b402b35d38a9fde312c89b82297c1a5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifb70a30f8bade95f402e71f95fe6644b  <= 1'b0;
            I309fa33562370e339c19e2377e6a6a7a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I592a495aecc800236c3470ff8e6adbb5  <= 1'b0;
            I7d06aed81222a030837cad2074c68e19        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1c8024aa9d81704d2dcf63e34853f8cf  <= 1'b0;
            I835cc6af0cd8189035f2441c2e0d3100        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ief03713f5cf37200373a20d42c7fc9eb  <= 1'b0;
            If6f768d12f04087246a0d65de1aef99b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic3cb34aae74c5f1a870b3635f8a40764  <= 1'b0;
            sum0_00013                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie4b180e1e2cadb865b0eaf6509f99dbb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifa3df8b249467cc1e827c69925ef415f  <= 1'b0;
            Ie329a11fc3f6f59f6f1790612fde3250        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icf3ad912aaeaa0c5cd1ab0edb898d6e8  <= 1'b0;
            Idb7ddbee4076f7bf49177e69f5e4d112        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib774f380e3d7cfd1f5f064e93d8134b4  <= 1'b0;
            I614d66a7dca2d08efdfdc157ca803d5c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic07c650e6e49892a41cfaf3a37471426  <= 1'b0;
            Iea16eb0ab70ebb1bc47ae55e11ced62d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib1073489d63ea33d7f3892f4ff875358  <= 1'b0;
            sum0_00014                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ifa8db43284d5bbebaed4f72d65cf9f92        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I174b6c36f2af82f8047cc76543a3b4ee  <= 1'b0;
            I365d9f3e8b2a9890427f07386deeb093        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I953b975a89adcc88039284970e9b3404  <= 1'b0;
            I466aaa0b6cde2ade1901797b8c11e32c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If2b40d249c531e10cc22d1335f350441  <= 1'b0;
            I7057e329a65ab240ed6cfa824307af65        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I44ccc3ae897109dd51f9afeef93daca4  <= 1'b0;
            I624e50e3457d33d12680eaf8e7c34aa3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie9236599cea94cfb603c6b977fdbb44a  <= 1'b0;
            sum0_00015                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9f356fd6820c33fdb5baff05a781e192        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I25f1ee9cee4d04bd8fec1fe601d016d7  <= 1'b0;
            I39b9c7c664fe7017731877d145d55b44        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5ec1e530b9007a75a778af4d82ab427b  <= 1'b0;
            Ic62ffbb9e58e0d08b0dec24bba1dc6f2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8a9e516aa824260998d10db758642bb0  <= 1'b0;
            I8da2a532288fb817e7dc0cb7b4e3761c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I70dd1350d65155ee7b562f4c79024a3d  <= 1'b0;
            I6a6e559f5c98f846014e8107fea5a5d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic9146d8b3dd0c612073b70b8a8791e8c  <= 1'b0;
            sum0_00016                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ibef9219f577b1a62dfdd77296fbfb24d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I857d3155df0b6dd704514b039c66fa97  <= 1'b0;
            I52e6688b5bfff75529d18e20b22832ce        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc1b8aa2f81a7fbd87e4f5821d14bf01  <= 1'b0;
            Iff22c49354eefca0ea3c5959c14b782c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I68b585571699a57bc6ba5e8955467119  <= 1'b0;
            Ie5377bbdb4111ed00356d5b7737102f3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib70e99c3acc76286a6811bcacc9284de  <= 1'b0;
            I55bf0f3379a8c44634b8f0a3d06c049e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iee17ece482d04964d3c21a092ec955a4  <= 1'b0;
            sum0_00017                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9bc9541607f4f6aedb686cdde297bcda        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5a247475beb737d470f03507e55f5b24  <= 1'b0;
            Ia4620554fbb1d81a71a15a846e4be2f5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I13b0c9578f7b6b3b7e6704d7b44079c4  <= 1'b0;
            Ibb31b35388ba8ba2ecf98449308ee67d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I41eff06fe1dea8be4613945de596d3ca  <= 1'b0;
            Ia20410fb3d56587f89a54c00b943b305        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I08f22261d5713c0636d77c7938f592d6  <= 1'b0;
            I9d268f3da12e35b9a4229b7340c0f018        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1c7e41b9cb1bdb6f649c88c0ed3f4100  <= 1'b0;
            sum0_00018                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2fce29bd666082eedb2fb3ec8b5ae4dd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idd59a5357d4c835379ed180ac0924bf1  <= 1'b0;
            Ia1e8b61e2579a90f5c88ded11c7322c2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibe7e5c2cb9c50eca34a3859d13e83a92  <= 1'b0;
            I8cf3718ba65b7fed72e3955f190e34d1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibf5c141c5cc0a6a20c05b52bf8282476  <= 1'b0;
            I7e802d300af54d394b4ee041798c0513        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0038305f94aaefe2cd1a243580d95932  <= 1'b0;
            Id4fd5a4b97cfa1e176a26f3a823c5516        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5364deb983adc2ae505ed2b8c57f876d  <= 1'b0;
            sum0_00019                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Icbf8d4e75fc66c05eb49c5075696fb07        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifdb5589982db805a0416e1c01276249a  <= 1'b0;
            I746a7e90adb2f213b75ae12a161aca0d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8bb5522183b65583fda83067990b3e94  <= 1'b0;
            Icb1029aaaaed8c698862ea9c5e22132c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1e77fe6aeaba852aba34ed37dd53add6  <= 1'b0;
            Ib93ea7028c172373b53cdafecae32a67        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9171019227f35760d02d0c8ce786f4d3  <= 1'b0;
            If9628275b000e418f3903daebfdace92        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6e92a48aaab94074a555efa9bd1e7243  <= 1'b0;
            sum0_00020                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I830202fb6f08f98c7f71893a881bd555        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3bc094d67805664859fdcb66f1360e64  <= 1'b0;
            I6f38bc9359562f57c1603355e9ee312b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2518ccf385b3b677d95983bc550282e8  <= 1'b0;
            I4701b732d59c26e3790a63c1936f9a24        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7547c56b32513ad45d775b4502596d9d  <= 1'b0;
            Ib5d28d8f73d17ab6df6a1291e50c04ab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I013d84bfd582acc7accf07ec522961fa  <= 1'b0;
            I81259f391db792339824ad5dd1a0057b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0ec27b590ee6dcdd9c1086105e3b6c23  <= 1'b0;
            I6f09ac63effe67a86798b9b4e1690664        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4cdc955fa9afc75c2c977de4ec540e1e  <= 1'b0;
            I370b4b3a0048a93ba374a40e170c75a3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ieefbb5d6f4ac1e586832c5c0f513c5a2  <= 1'b0;
            I3f8476d0aa0ea2439b67ea1a4adf36c5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic828cdd5dfde844df4c150921af2a443  <= 1'b0;
            I35b52dba10a8a5b22b518388fecac82d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idf1ecab26889c4adcb835fda6b1cb368  <= 1'b0;
            Ic7db274ed18e6fdecf30381a31238777        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I00d3f14b20e1ea7d726533386e0eba27  <= 1'b0;
            I2c4e538a8db759e9799541d9178ec61e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7f720a18542528f0c9bfb14f699ff4da  <= 1'b0;
            Ief6d4c3f5ef8663e111ef99347b023f5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia98a6f01e4eb5bc74d50d350e79be426  <= 1'b0;
            Id95e964e5faecb52c72669b0d28a4bf5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I182b43872d50de6f7afb700f178b160e  <= 1'b0;
            I0fcef4538102ac6d24aa7090d5405afa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic9b72b2a91d951cf08cf54ed215ecaa8  <= 1'b0;
            sum0_00021                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I055019e38eec6badd1739033d43d7d97        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I93084ccf5b5e4efaee968b497bb2a775  <= 1'b0;
            I35c20a6e823da77a870b421eef2e0a95        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id38852415486e6989b89a0d85ad6771b  <= 1'b0;
            I32cc12cdacef1a4ef64577e0fa977f46        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17cf58ef5326978c62c03c56090a299f  <= 1'b0;
            I26b3f2360ca4a8caee61b2f3a3a08267        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie41ca18c7d11a47e274f9c33f75393ec  <= 1'b0;
            I5ef9b7dc0c63e9ca6a5fb5f7ffa06041        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7b80b4902fe98c10dd72c9eb082346e5  <= 1'b0;
            If881473b05090f40a027d7eeee7f7ed9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I20ffba20af04b99954bf719589e90d1a  <= 1'b0;
            I23bd59ab5b038935301396aaf2acefc1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If8fe5af7e5c3c97b5a713f6bcf919f1f  <= 1'b0;
            I874386d94dacf84e699d159af1a49836        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc5fb0f3a04ab32948e249e088a11b11  <= 1'b0;
            I95bfe51a759bf4165168e5e3b99d6b34        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia9f1e580e8f441394d719d52a7bad688  <= 1'b0;
            I4ba5b2f9b7ec0937ecd2c9945cf6de87        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I02849282dd1bd663fd39baccf41762f9  <= 1'b0;
            I0b08fb8db0e8a1de3d416907c87fe700        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie4cda4648f6ceb76b8fb74f290ab6439  <= 1'b0;
            Ie030d12e5acf9ef4975a17c83b2481c1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I24135210c23b2422a42c90ee25594191  <= 1'b0;
            Ia7a0e852d3dfcef950804ea0ebb0c80a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib08897f9216599042f7b97b137e07fe1  <= 1'b0;
            Iaa4c38d030eab2b7899399aa0d7886d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I51e14ece9ab6607f83e6ba27f3f046a9  <= 1'b0;
            sum0_00022                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Icce7ff1d652d4d9c2be5ecf679059bbe        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7a626ec321bf963a5401892a7e3891c7  <= 1'b0;
            If816bc5eacaea23443602e575ddf60b8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If76f04fe0baf171d7df2c0cd849aea2b  <= 1'b0;
            I3b224a4ded05446cc5300d430bdd1947        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia9c8cc5e3becf3d48feedec8fa2c93a4  <= 1'b0;
            Ia5fc5cfb0e52237b407b37a3858fccb5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If3b77c41fabcdb283f2c6fdacaa5e9a4  <= 1'b0;
            I92f8ba6e7f8e9b30fb5b6973eb8fd03e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie5373b01a92f2ff85be8077cfef2175a  <= 1'b0;
            Icdfa60d2a024dd934f7e6639c6cb2c28        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5109afc4dc91780e05704ea5e1399e3e  <= 1'b0;
            Ifff70b976513eaa42b6bd4b80c98611e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3e0b41bee4c76eb5f3340ad23bfa01ad  <= 1'b0;
            Ica12fa8b631b70a6bbe9f6e92bf73ea0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic0732810fd355d59a3168be896a0f9ac  <= 1'b0;
            Ie69c255335760f706c644b115887269b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I220e32641265b46527ca61111f7ebf1b  <= 1'b0;
            Idb06676b41de19bc86eae34c292183d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ice59d2af73d0b0f2ae91a2ef0c2b7f04  <= 1'b0;
            Ib21d2306d5ded3406fac754e69a10d20        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic308610ea8bb62ecb6094192e02dbdba  <= 1'b0;
            Ib41d1aa2dcf81879976fb8964cbf6f79        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I33ee415d85e2bcd8f975d34b880f6ea7  <= 1'b0;
            I5f8f5e246f008b8d8c75f72828337bab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie61f299252b8fecfd3e8634b64df5a90  <= 1'b0;
            Id6625e78da0e14d2eeb19cc8ac6520e0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icc67656ad2dd3fffae4e5abe02f8fff9  <= 1'b0;
            sum0_00023                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6d9ddc6afa559ac35c042df1a9390ce9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0c47ccef4b55410286248884a7249703  <= 1'b0;
            I9334055c7833676469670372d3c5cc31        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I94e4041b482064334fd0ed92b91bde89  <= 1'b0;
            I0c97d772c737c6ff85b584bf69ccaf93        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I39d3bce4060032a81e6b6a1c1805cfe8  <= 1'b0;
            Ic6ce97ae85d91dd8a79f3f9d0da375a2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifb422c30663eb4824caa72326b238df6  <= 1'b0;
            I83ff9a2750b298b0f7c9b6ce13f574af        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I41ab6fb6ec6ef7ffff70e50f25f217b6  <= 1'b0;
            I85699a2a05c343a6a9e828af6d445e9e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3ce10718a2211184999663c3c2493cc1  <= 1'b0;
            I51f6e39b24b2554884e381be79f47ff2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I877e8d94236c3d8b0a31858a98fba5d6  <= 1'b0;
            I9f65fd05c6929300860c8cbbde5607f2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iff2f1716cbd73b406d8f07c22dc79fc8  <= 1'b0;
            If09761d8f06051d4287ee29ac9c9fa19        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibc48fabc172f27ebce18d0a9b5120dc5  <= 1'b0;
            I33bfbe0bcca6d32c86b9576577e3f265        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie562ebb336e476a81f20a652d4cb20f1  <= 1'b0;
            If2921210b1c05ecbf00af3a2bcb96ef4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib5ee5a6ffc45ed1fece0822dc4619b57  <= 1'b0;
            Ib074e38e280474a782da831a3e0028b4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I86ba73ee348f80e2f9891d2ebc8a02ed  <= 1'b0;
            I507449dde0bc0c8f53a10759436ec731        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1e96d5af3d0e3fdce39530dfd0131a7d  <= 1'b0;
            Id55a3e3f2d75baeba71a345fad695c69        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I38352b363fa37f6f822fbc1a39100968  <= 1'b0;
            sum0_00024                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I20984f43d22671639a7a178ad15aec04        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4ba41864bb1d2130c6971e0b2903027a  <= 1'b0;
            I59f88336d6bdd50ded87d353fb5ce3e9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib68deeb7bec4ca3585d1a4dcbf8793f1  <= 1'b0;
            I488635e3f7ed77ea88199f5bffd4b1d6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ida3d808d100e0bba290f96ed9e744e65  <= 1'b0;
            Ie6893017d21c050ba10d206854f4a9f4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4d4901ff372f6820ca9c8c29cefa664a  <= 1'b0;
            Id3f68b4dc0ab60673208b7d2081f3533        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib99e1b93fb7fbda260d93eea3d24c3e9  <= 1'b0;
            I433756b944e061a824a89bda241e879f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I019e399a1cef87745e025a7d74e94db0  <= 1'b0;
            I2eb60a922aa4f7482dd92b9351d53a2d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia8974083bfd064f2c27dcd421490fcfd  <= 1'b0;
            sum0_00025                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0867979e1b159c8ceae548930376f482        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8fd5787ebf758919e7cb75d7419441e8  <= 1'b0;
            I4accfbeae8a5ee0dbeab23ef3a116145        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id14074d5230885c38b89b09b130ecf68  <= 1'b0;
            Ic7570b0b7c5bef5758f68562ae4c90f6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I86fefad34d3c864dd0e725133f303b4f  <= 1'b0;
            Iceadadc4456881fdeea85934a9bf4d6c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1ca188bcdebbf41d84f7a5220bd1d195  <= 1'b0;
            I7b2b617ae67424f54961eebce42de77e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifc640243288c9b37b7eb9e00351b23f0  <= 1'b0;
            I953f0f8af76f89b2d9ab4abf19fb411d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3d149293f106ae8680c7f4702daa0bd6  <= 1'b0;
            I915b4736dcb20f831d02e48f4e79f008        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie232799bd6c4ec99e24c78f3ad798265  <= 1'b0;
            sum0_00026                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ib7eec587348ae1ca1f00c0a3ad10ad27        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifebcf64858d5e2d07ad7894d6182eb11  <= 1'b0;
            I001a212686304248c8359e5fc01227c0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibab55499323660588ec82ebd07ab0572  <= 1'b0;
            Ibb7554e012c0fc1223c29b759c900666        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I89af7644c48a80d7d22f50b008d35841  <= 1'b0;
            I9aeb9c42b54a05be6bf9b7b88b6860ba        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0152dc6e6a7acd72a2144623e63998ef  <= 1'b0;
            I6a5a5966965b0790b906c6fda71aef80        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I951dedd7af44c3865a8f36888432d0c9  <= 1'b0;
            Ic943083ca65ace6c42d73f4234739a06        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8188dd7cb03854c6f709de06ff785d91  <= 1'b0;
            Id0b321686d4c39621024cf0dd99822dc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3b30b4ab00a49e10a75587aa324d6132  <= 1'b0;
            sum0_00027                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0839dd3787442f1b79b87e02436bfdce        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie50aca688b3433fad7565998cb900155  <= 1'b0;
            I89e6a9fd97d8aa4dd3b832c3be4697b2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3342fe0c5d3ee5021892d53eb45bde21  <= 1'b0;
            I93d4157f48b132642752220059861e98        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5134b762ac428bed07ce102d8927a418  <= 1'b0;
            I8fc4faa2891d7fd3479ac1f788f481dc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic14f948884da19a272a4760ffaab9ea9  <= 1'b0;
            I440f30e9cb4bc89233b46ea00b4cbeb4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I46e1047bca2b38e62b4de80d1d2249de  <= 1'b0;
            I6568bfd8780c11e0b1b049a01f92abd8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I866b30a63b3b5fb708934a1cbb0e1d9a  <= 1'b0;
            Ibf7dc4da07f9955d5d4c7e1f63f1ad68        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaddc1f2e822fd2fe9d9046d759a82cb4  <= 1'b0;
            sum0_00028                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I7ec1a328587b72a39c462083efea0ee0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If9285bf7611bcc5ea6432215c349e021  <= 1'b0;
            Iaf028e7ab4dc77a7649f15d603834b5f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id277f5f05551eeb5dec1701056330da1  <= 1'b0;
            I58db79a8e9f0cd1ded379897ba2f27ae        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9963d0b24763ed8038b1f3922b8f9548  <= 1'b0;
            I6d3cb4ccb4e51c7e6603d0abd1a082c4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia98de3691917dfb63bebdc3f8655c8be  <= 1'b0;
            I79f75f49ea8a29d684af396014b2f3ab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0bce960fcc58938e6a1e01b912eabbf2  <= 1'b0;
            I9c5ecd86bedb189fada40fae9d751a68        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ice5f7168aeb940d48093cc9df7cba36b  <= 1'b0;
            Iad5f06e1989ead7d306c70a3b02cb8f4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I859d795a7d141eb777c1f3c038203794  <= 1'b0;
            If6d1a410df5a4aea6a01337a6074fbd9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0dccb8eaad52ce4d780696a8485420f1  <= 1'b0;
            I3bc40a4db14566b5099b14cee5f61135        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6d4fc81ced37c159303c243af04d345e  <= 1'b0;
            I7e683fd8235d7cfbf4ff407a286f07de        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iefdb8bd28839af9413a3906cbfe715e6  <= 1'b0;
            I97afcedf05e588b7976d6005191dc916        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0615acb0f7cf79b5f6ae8e91cb525dc9  <= 1'b0;
            Ib8d8eec0aaa662adf2837c9b705fce7e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ieed4c810a5bb69de112522dcf00b16ed  <= 1'b0;
            Icbd765be950123705955e2c5d7ace84b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If533578cacb685a95afbb8e1c05d3c07  <= 1'b0;
            sum0_00029                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I706e8f5617cfae1e6fc83db18c8b5fe3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia858ff5551286beffd4cf82f876d30ac  <= 1'b0;
            I1dd8f8c7f1b673898096b1f3ae383197        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4c66570630a650fa7b9bec543f685487  <= 1'b0;
            I10ca8978cf4659265ed25a27d09acc1c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If10f33385e236eaba56cbab8c2883399  <= 1'b0;
            Iec4656b32460def4a608b6b0f6486af9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7cb58e4c486e683faa4acad4756815d5  <= 1'b0;
            I5f4475897d1d58965da1b35fe0ef8c01        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I452e51cca9acec44e36e4efd21b43034  <= 1'b0;
            Ife61469306df3cf220666b187f1496a9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ice0234f25de4ab1f03a3cb01a2d61dbf  <= 1'b0;
            Ib49319b9dfa4914f92f423ceaf840014        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I12a18a1f8d4416e9bc8abee6ac3dacfc  <= 1'b0;
            I93ff2f879233cac9b9f0dd2f4c082c09        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id17ada8dae3f9810d1892d34f2288859  <= 1'b0;
            I44597d694e9c5d29280e503d72a27c8d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia2c5fe53cb5b318fa63d09881609655f  <= 1'b0;
            I04a19448c5e75af8021ad02d1a708bb0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I579c7926e7b78f4ffc606adc10522f53  <= 1'b0;
            I71a3093121c2f19dcd1412b468652fa8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iffa06a336949f56f4e5a88a06d8b7e60  <= 1'b0;
            I3ae09c82029c617034fe6aacbe9e94e6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaf82668eb49248709540f2f529f1b3e4  <= 1'b0;
            Ie7af6b3b441f910b000a333afad6c76f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I90b3708abdf742370f06cc513ee307e1  <= 1'b0;
            sum0_00030                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4d71dfea8407aa5b5cbb991bc4fea963        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia17906696bd0e095d7a5297da2e049ea  <= 1'b0;
            I1a082caecc831a90e74674ba35da4183        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I180d4f3b23b518271d7cb8189fbeadc5  <= 1'b0;
            Iec1de44616a2354a56ab1f681059d4c5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id79636d195efff260c430978f0bcee9c  <= 1'b0;
            Ie3c2318e64d0e218c3db557404c4aac8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idbf4ad11ab2a27044193448c8739fec6  <= 1'b0;
            I9a251d50f41e51b1a5cc2475f267e8a0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3051f561a5e1131ebf167cb6ccb5adf4  <= 1'b0;
            I9b5767a49f7b9dcb8fdaea924835033c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9322a2a61900943075bbc23c72a3f65d  <= 1'b0;
            I6ca1e6700a19d03621a193c7240bff54        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iedc463e359dd3003d9f7e50f3e858e93  <= 1'b0;
            I931c597ff12bffce581f653346202f83        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie7cfdd25541414ff3f8d6e5d7677fbe5  <= 1'b0;
            Ia3a2c5d59f6340917ca3933c05ba4678        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1e93f0470d2818249f1c28ef2a399a0e  <= 1'b0;
            Ie83d0a8ee5ed214bc7577467748aaa04        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5d6e576b0fa7e3219aaf9ccc345085b8  <= 1'b0;
            Iaac29552e5fc65aaf4f0116f917b707c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id962beade26396738ba0e97f67d5e261  <= 1'b0;
            Ie2c8eac7204b98139c03b6fbfff9af36        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id0ab747d92288f23cef793567b2363d1  <= 1'b0;
            Ied7fcdaec662cb3c2f89f131986fa102        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie536879e6fa9be65376d7f00e0fc40d0  <= 1'b0;
            sum0_00031                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ib16a17d6430570b45a304d847ee2b11c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibf312ae4f51fbc44b43848f9df62a45f  <= 1'b0;
            I42169e454756fe4d1c5f17f2eeb2e091        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icfc03646b36b971b9fa57d04a26dbfc4  <= 1'b0;
            I6fde38a3a92e06fa77123e3279813c41        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4f134c0669b5a6a8c7e03be7eee30c6c  <= 1'b0;
            Id8ee16437e8d6d6da6d37440e04097b6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6c765e677f42fe600b848698c8a78349  <= 1'b0;
            Ibf249d8e5acced9b064132575f40e001        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I284b23051c85300c2a1e3afe8f25e99e  <= 1'b0;
            I580659084e3d17b48de6b1c66154fcf5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9b560d9baf8a7422b0dd84720e924ced  <= 1'b0;
            I7a14e45d43ab77b265501902152c8616        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I457ae11ad90c8478751eb4b42764e158  <= 1'b0;
            I81ba868784103e0eb05a44d981d4d666        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2b7822d5d77aaed61eee87570564df76  <= 1'b0;
            Ic6b88783957cbaf253648a30b22f6b1c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibdad0ab78e4404c852e60a2b04c3a5f6  <= 1'b0;
            I4103c218a85a1d08db5c4f4b5686b2e5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic4efba3932e598784f5b9ad6ad04772d  <= 1'b0;
            I0e6c0958af503e4a120a49d02a432863        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia03836a4e93d2f36513227d1dfaea0fa  <= 1'b0;
            I8f76b31e8f15c0e5fe24dcb723418111        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I138fb0c48f2d27e3315e237d9e61d653  <= 1'b0;
            Id1457221b58344b60070aa026436df2c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id0b1c46fa4caa63a4c63a44ba3c5ef8a  <= 1'b0;
            sum0_00032                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Icc31966508e03d8869e81d8aeb243705        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3566033cf5c9a06977c9182925750707  <= 1'b0;
            I9dcccf542ba434b6e0fde6f012f98f92        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I02812a8a833bb69eb168a1004b6fafdf  <= 1'b0;
            I51ccbb824a5e1e340eefd173c4491728        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie886c5effc85f1fe0b6411db4a2cde77  <= 1'b0;
            Ib7ae1730dcd8bc708bbfcc6a9f97ac66        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibab1d13cd6a4f7b0c79c9f845339e53f  <= 1'b0;
            I4714f5c91203fcfa552f0fcf71b87442        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7b813d83b13bb7bc13940cf5714c06ba  <= 1'b0;
            I3b6d1e84fdd1019249886fa5fe65895b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I09031235f61238b0e32ff52641aab70e  <= 1'b0;
            sum0_00033                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia8a7d4207dbabc7970bf36f3fe74f72d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5402fd208dc7ca81dfd2920a9cfa2715  <= 1'b0;
            I84047457b43ef33874f4550c3b773460        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia01c82761aeb124cd92fb15ee367ee8b  <= 1'b0;
            I5e51563c3e69beca0b463742e6e5f9ee        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib1a40247057324b0bd810c844bf11f51  <= 1'b0;
            I6c8d14e31c80811ccab1b6ab09d28089        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied8bd4b6fd0e4fbcced6d20eb7435f55  <= 1'b0;
            I50b3b7490c9b65b6e662cc86b163a2df        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4ee312036de8c08300c358edcff1e1e9  <= 1'b0;
            I8351a2110a3d73ad8803cf17e3317017        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I477a920e2326828bf026b0a6b6a18e2b  <= 1'b0;
            sum0_00034                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I1e6c696951688d581f21ab2302593335        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic11a6b77b84c44180eb99220a0c4c9f6  <= 1'b0;
            Ie9840e28133eebdca0be313552195c7b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If0970d9f7b053fce3ced3521b4885588  <= 1'b0;
            I82812258a8032e273cab7139266be1b6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic7ebdc317c978eb275eca41d5b9106a5  <= 1'b0;
            I27ab6fd9927518e29ed36d7a7a241498        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibe3d3e6bc58efc2e9d9eb1f96cdfe424  <= 1'b0;
            I05b0f33a3808ac53b29d8d8309447650        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1dd4671765f8826c2fe20c592c5e32c8  <= 1'b0;
            If150ebf242231f0d22c996a71552f6eb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6cde57127c5bd2732e71ecb7738fad6d  <= 1'b0;
            sum0_00035                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If2d0a2b58510715e74787cb60719cb5b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If6ce2fa9f0b8bc74442ed8262b5089cf  <= 1'b0;
            Ib6745a6d17034a29501e022bd846bf2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib0001d7298ad1f3b1c7603173a70d8b5  <= 1'b0;
            Iae09c127dfe86c9f7bdbeff447c777f5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I05e739fc87e962848f265e2c73338cac  <= 1'b0;
            I742128de6b237ed48e3a7ccd3788f0d7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaaaf373f7e6f55214915b93da9bd71d3  <= 1'b0;
            Id5e8fda13ba8f6d95d694d0f30da75bb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I47b0847946b0e00961233ac0101fa2a7  <= 1'b0;
            I1aa5a04e40f9b1685c77e4d101c3ccf4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2f23d4cdb6f5f827513aa60266936e4f  <= 1'b0;
            sum0_00036                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ife1adea26d13bc299bb2de241ad4a6ea        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia67f9b902a21de0414eb8dda52171991  <= 1'b0;
            Ifcf6c761f0f253921710af87ab1d2247        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I87b10521099179c18652c86d5887c908  <= 1'b0;
            I1478e6a9113c124bdc4361908af6643f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I84057a3b319ab3d6a2ed8f2310f970fc  <= 1'b0;
            I0afd42151925883835844cf5deef6156        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I67d57e38df8cb35ca686ac2eb44e233e  <= 1'b0;
            I2b4ab0aadffb3a1bb86f45ebc8acf085        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I23955b54e486f0f0d21a2809a9472b86  <= 1'b0;
            Iffa867719ba9c31a8756cc5e6bf81147        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1e11f0088959aa40b4ad1a047b59caf4  <= 1'b0;
            Ibb62b6cb003f0d5549c864075f23d19b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I68c35d63dc95baff41b4dc27a86d2342  <= 1'b0;
            I3690d101ae99f258cc58b4482cc378c8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I837183265ee22d080e81fea468ab0887  <= 1'b0;
            sum0_00037                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id597e95ce8a168ab67890085a26870d0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I413b1c1985a6c9c6f202e85ff901e3a8  <= 1'b0;
            I98df60eb8f65641f9cccce4023be905c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic32c6734132776c290155a80025fe366  <= 1'b0;
            Ibcb4fbdee372353b79c460cdeafdfe4e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I624958486d181501c7a8ec2642cb503c  <= 1'b0;
            I74dbf75966d047a4a9e91c1bc793666f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I04864c28351edb33b61a103add6fb875  <= 1'b0;
            I79b8d9f9447c4c1b551ec6c1e8903040        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ida3dd5e990ce3c237e9628a9a090901e  <= 1'b0;
            Ib34b66548621fabe0753223712b1369f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id182a776b03f48fb139c28194ae7ab6b  <= 1'b0;
            Ie5b3eb4c00bedfaecc3215d43ff28362        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0c5539373b3868d0664a92157b4b4226  <= 1'b0;
            Icf3a1b0b6dbcf959b44379024f3c4169        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic0191941cb968bbd7644c21767423d2e  <= 1'b0;
            sum0_00038                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I918c2bbe7c71f8c6a07b0bad8811f4e7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I163cf58b9a308e0439a8dc7c1526e6b5  <= 1'b0;
            Iedd960a21b1c08b4a5293cff200218b3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie08ad9bd71329858c1742c8f571a1c36  <= 1'b0;
            If9722c28747df3a59b0ecf8200907e98        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3c10d579f80bd0106506ad047d75f188  <= 1'b0;
            Ib83df72c8b73a333d0699a8bbbec16be        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ieca2767ac27170058499d83016447aa7  <= 1'b0;
            Ide3798a77f709a9f694523338b081f70        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib9c194ec16f435a9357cb344cf25bdcc  <= 1'b0;
            I0a9722a805604433562f85c62b168b96        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic920452d5997a8477724fa78c86c0fba  <= 1'b0;
            If9480ec13cd538ed03a43e56bd6264a6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6eea5fde8e2517554ad6ba25018572dc  <= 1'b0;
            I433ecf86b7704c5552e5fb5cafe0d529        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9ad2f6fd2d7f68011fc926ec9abd5c34  <= 1'b0;
            sum0_00039                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8326f0b2d25139609e2c5e466724f224        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied33f18cbb778d5ba744d249f91c950b  <= 1'b0;
            Ibbe211d9955cdf2810c9003d1fb78074        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibabf61085ca7af8dfc7927b3656a76f7  <= 1'b0;
            If15e950b569a92b590127d0ca6f20a16        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddc5b5b4501f9f13bcaf22081e5a70f4  <= 1'b0;
            I03e0532841ba39eb1d4ae823c4de2f7d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I67f87fbb746dd937fffc534c596f36c4  <= 1'b0;
            I1be81a7b73987ee023e396cec87312d1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I45bdd0cfe107da0d57cad1333bf95e3b  <= 1'b0;
            I4ce1a767a78673590c4074f3f03bad8d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4d54dd2ee2f32909098d3cc2b6689220  <= 1'b0;
            I57806bb7da625881e68ae315543f70d6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7bfb4c5d9e22d1bd8811844d9c74dff8  <= 1'b0;
            I8b0ab476b4790150575abb06bcdce2b3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib9d58222da98f29fa302b4896594fe26  <= 1'b0;
            sum0_00040                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8846a8961b7d557df4fc62dada679c33        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iea3e35ece9fdb3aff3b9ff5369e9a7e0  <= 1'b0;
            I7909a0f96a92e93f95023cddc742a5eb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic44eab478be232721e7a43d14beca32f  <= 1'b0;
            I43ac4857544c0fb79d04e850435ef673        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifab075b1437495268b6a3be4cb022e71  <= 1'b0;
            Ia6dfa47c465325c1d9fb9b9c5ce08f01        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2919272e9ae3996a3e1d602ff72ba86d  <= 1'b0;
            I2e9eda5bea0cc3d88359ce8a7a82f21f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib6fbe376477afa58bfcc17a8564f78b2  <= 1'b0;
            I53ec2486418e41b2ccfa8fd82777eaf0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I659322a9fd0d5eac514437b02e0491b3  <= 1'b0;
            I18387c05cef21970ecbc39c20a87aafb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic68f500938d80460ffdb33a0adc48298  <= 1'b0;
            I2b23eae78cb925008ad59f45e80e165b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If5ae6fbf843fdeee17945bc5ce81aec8  <= 1'b0;
            Ic69eb7677638a90b7a54389d47be46de        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I94460b6ce7b776bcc5eca149eab80c26  <= 1'b0;
            sum0_00041                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8cb9a216f4da7c27f678386cb214c59d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3347717ba9556e69de30ce7533d4f5a4  <= 1'b0;
            I48cb720a6323697084ac3bbd8fcadfcb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2db290170ddae8dc52ce07edaf48b365  <= 1'b0;
            Ib8dc3c1885c92cdcce7fcb58d65d03e7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idd775d9fe6fa8dbdbfb07d4071b9caa5  <= 1'b0;
            Ic3aa51a5c758405fa6e2dbed707555b2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6cbc06919b9c695d99621db6f8d768cb  <= 1'b0;
            I4d418179c859feb8bc7d750416bb1004        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5b8a1e1a6b904b0f6822c224ee0486e3  <= 1'b0;
            If207b2adc6f668f85cb76bf54673fe18        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3f5053e519a928640ae49cf4e5b39d1e  <= 1'b0;
            Ib08b8067ea75e210e83526ca4a37217e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7c965c047d862c973d09a81abe03a845  <= 1'b0;
            I95b30f641cbf7bec1886643c4468017d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9b8023f4dced915cd52c91bc9d4ed78f  <= 1'b0;
            I1978531a6f8d1d25ee6d404025ec4753        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc6b6357741c9887a9db1037ccc2d922  <= 1'b0;
            sum0_00042                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6c9698ba88db16b8d22ccebd58cc541d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibe97860165dc5d9a076ebd935385ae51  <= 1'b0;
            I0d8ac5e09b200a55bf5ba6f834cc9174        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I777ee54ff20d0544af18ad8a870d6915  <= 1'b0;
            Ib58b7d3d77a54ff1a180c6fa5f1400e6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id18c5a1d4eaa73a94e699e5f9e3c3d35  <= 1'b0;
            Icf6b990098b7ab91800bfcf1e643153c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I72939e49bf2d9c6a84e404419fc644a1  <= 1'b0;
            Ie4308b9ac6fb6de9329ba02b1eeb0e8a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I57b7b48f13436b19a8d6a47e014eb41f  <= 1'b0;
            I01d4f02a356c51d7e4e1993de0d8eebd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia3ef2f70c5abaa852586a33c505aee0d  <= 1'b0;
            I36c351e3641b01cc43e1dd5de0a649e5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6d423a7d17e05a3c597ec6ef6c5a7cba  <= 1'b0;
            I4fc983e94c5b8f7bafca61fb0d351c08        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I48e3309c61918c3991852b45d9c72ea5  <= 1'b0;
            I1fcb82fdf96cda14a55fa6358cb62c1e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I472352e7027b9df2fa957d9fd68443ff  <= 1'b0;
            sum0_00043                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I665e54ea6bdca483149d3b7f3ee42a2b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idbbf2ce4a30787c5f07c3b908a73da75  <= 1'b0;
            I925df2307b5af6d1b166e5435641d3bd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibc9a860879ccc58c815b9f6caa23320a  <= 1'b0;
            I9b14f48aa357d09e460a445da86cdf89        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia71cf07b645c58cffe33be1a9a960eb2  <= 1'b0;
            I78e94ecb6c92fa8ee24edaff33b6f82d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0ceb14ac0187d804f9692e0c55b8e941  <= 1'b0;
            I5ebeb9ce5adee72a7c9527ea6d3a3028        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ief18a19d451f05f6051e3cc8de16d73c  <= 1'b0;
            I90d7b28ec09142ca8086836fc0c5ea0d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I30be0b18e4415ca50f2d8149efaaafe6  <= 1'b0;
            I27d9985415e6d0b117e5a4c2863aa7f8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7ec15b73b2811b44e1e50c74a9f921e9  <= 1'b0;
            Idf9b563e5d10c2bdbcc07e81d74467eb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0fd2f706e374a4eb57ee26ab50201e15  <= 1'b0;
            Ie351922194483938302ff6cafc477e4a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I44f170d02bae7fe044456e125a98451d  <= 1'b0;
            sum0_00044                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ifb2da5faf236ca8636677bc1dc35c4db        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I30c0fcd89e0cc7c5fa348df7b4fa2ccf  <= 1'b0;
            Ie15825d216685ae241b528fa9c158ff3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I13a98f98c54b2e412cd88c96f016c41b  <= 1'b0;
            Id92c2d8bc61245c0c8e40bec2424c3c8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9890f7fc708c7b8cf460849b4a30025b  <= 1'b0;
            Icd9fd8d7114b6e894dbee493b6797df6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5e69e930a318dcb0594a823b3129d650  <= 1'b0;
            I29ff688c085f2b18e7a3af969f18af76        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I403303228c0df825f67436f4a7e64061  <= 1'b0;
            I6d56db9fcfe69dfcd747521a1ff62297        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I946246be5b4745508b7d4b578f83aaa2  <= 1'b0;
            I2f17f7c79a0118b39a63894917c6affa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I95f0acd4f955058041c035789c3a4d99  <= 1'b0;
            I7350af5d5ee09ad28c459e3674a829ab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4082b3564c1949a19ed35bd5a88e1ef4  <= 1'b0;
            I67b6415c5135e3d6a41d56d98d3f8315        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia7606050c683ecefc510ba92ac539a9c  <= 1'b0;
            I4a6fffd8bb7244599383f2aa3a1c8916        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5446c1c323774715371c73bd1be66697  <= 1'b0;
            I7dbcd21016231546b76aab175cac9f74        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3a8e9e7d2cd6751e8500a5567cef5acc  <= 1'b0;
            I9aeff3dc44ed0d0f32518590a900dcc9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I621b20d29d3a9a9f41065bc3c3bbd2d8  <= 1'b0;
            I988b7d5d56d22d2c77c5c8c125129a50        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I263aad78110a1136eb7012c6983b2a8d  <= 1'b0;
            Iff35cd97f2a6d37a7861b9cc1a655ef5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If4308ed204e33952c9931f8fe257aca4  <= 1'b0;
            Ifb3f2a1bedfe41c73d198046a2a3f177        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddcfab4a7022e0f12fd20cb34e9b9d02  <= 1'b0;
            I37ddc6ccbc188a3eb8c33a501de820be        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I759409e242eaeb144a53e630a8cfd514  <= 1'b0;
            sum0_00045                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ica608f1136da397e2ab61bd4a5d83201        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5f96a68d20e3ebc71dad4b43305baa20  <= 1'b0;
            I80636a3df4541bf29780bcb4d0ee48f9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5d92fdff96b9cd64f3af2b28b13e9956  <= 1'b0;
            I9ad99d544187db3cc7090b92c9933a31        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iab2f643f81921ed8464e1bbd9fa8c68e  <= 1'b0;
            Iaa8a2b6fcd469869efcf0b75ca38e68f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17d7f36fdade16dbcf621fe302bd7e57  <= 1'b0;
            I9a171d2d8eee362a0073ab7b139d3037        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I23afd747ecece714e32fbb896b5c022a  <= 1'b0;
            I84cdcba86bc5991feb391003cd7be40b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I388528eaf83566cc56b23485a9c05962  <= 1'b0;
            If9e5c3a848acce5daf570458f78f6aad        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iea424dd9d8916c4951b8746408b8a521  <= 1'b0;
            I73247d4348333f67a491fc607b15af0e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I73bbf90b625d56f663ad10f9d21d8e76  <= 1'b0;
            I021c745eee4b85a2cd91d9d8d2b18b2c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I41796b587316c600bf583edc62649bd8  <= 1'b0;
            I1381c0a0bd28b1c5542992084635b355        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7009c18515dd43d8dd2e5d1ee6779641  <= 1'b0;
            Ie74eeddc21428254a8fc4c3e293b5eb7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I797c9cb725f88c07be28f017871d17f8  <= 1'b0;
            Ib1d0f94258b45de4bfe610086d8990c5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I06b48093d4c9b0327c3efc6fa4ca7daf  <= 1'b0;
            I138d6d5d60df37870cdbb1d9c51a94af        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I04c734eb876aa722e84d6b9edd297978  <= 1'b0;
            I706378735e63e15c8d5395446ea41db8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifb89e7ad8ef661959d82b7c22f187243  <= 1'b0;
            If8680a7fc4f5532a660006bf4ca6a66e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id1dce2b9eafc35fa71df33ada4aac539  <= 1'b0;
            Ic59d1ff3051a95166c3c2d5a2881221b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied19cb51636bfb029ba8a2c390f97105  <= 1'b0;
            sum0_00046                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I54a551af28c505601cdfaf8faaa94afb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie46b71f55aef4d00168202431d47dce0  <= 1'b0;
            I6a3124c03eb83d41c16704133bd1cfde        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8c0c1a0a35f4f7a688f516c567242d39  <= 1'b0;
            Ie9ee27b9761af611ab96f0010abd47a3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I53222c82827cab7c770e057ae91bc10e  <= 1'b0;
            I305436919f84066a22ab1417ebabd737        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8015717cd36aabbf2cf4aa3a5c234690  <= 1'b0;
            I78e63717f436493b756efa32d66cdefd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic0c13c9a929c8c46e8702cef74de8955  <= 1'b0;
            Ic965ba971642db19ca773eb68dc0b9bf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I71d7f72d83b7410de31e09ea96adb95c  <= 1'b0;
            I579480a66a5f6331fb46de13090ce888        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1db4ea6916125702e7fb09d0f742e60a  <= 1'b0;
            I38d78b447217271a63f30f78b424e2ae        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc445d3f5b3b62562b0ac83e5f17e92a  <= 1'b0;
            I4c8d7e5474b19a7c63444d0cb6143728        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iee6e52d75c093a24eb4e5e0b45feb256  <= 1'b0;
            Ia4bc4b7414bf31305ec8f63e7eda61e7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id48fe0672aa98f987162931527e9f9bc  <= 1'b0;
            Ibbebe287d56c7d627f3ffcf706575e77        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idce46f6d03376bea1ba361e8c59f8bd1  <= 1'b0;
            I83867e6ee369fff7e39ef5c8d5398fef        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie79ce8adeef2c3c24a3386f054d0cf5b  <= 1'b0;
            I1d40df7dbf99674f987bd06db714a702        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0d41bef808860bde56d48792764612d5  <= 1'b0;
            I92f42789cb81760ff2973e3a5fe915c3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib6ae81df8db1dae269437861ee11ec0d  <= 1'b0;
            Idbd5f2a25ab05808721cf9c403017565        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I33ddee677715877c11a1df45cbfb01ac  <= 1'b0;
            I7ca5f07d6d3c2a045dfd55ae5214dd65        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I433dd5092cf1851cd196feade3cfa6d8  <= 1'b0;
            sum0_00047                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I7f4e1445c68abbadce23944b99d206f9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I71d3a999d88e591e102398409b3adebf  <= 1'b0;
            Id9f28016678e5e2127d9f0aa93e0b534        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iebecd2d19f9174d87deedc1a273e7baa  <= 1'b0;
            I6b939c57a8b7c7c51ab43e1b1df12f6a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I168afc1863f909dbcb6a9230db9f3e00  <= 1'b0;
            Ic5d0df586d56bf4cb322d4c3ad677385        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1c4b29e48d0effac4839037ae5688334  <= 1'b0;
            I2e287724873cf6761799eaf464ed6302        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I431fc2e9533012c8571d8158d4777dea  <= 1'b0;
            Ia7a10cffe31a53aafa1104b97543280b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ief72606c77113ae37845e4aa4a2ae5e7  <= 1'b0;
            Ieeb089c6a18791a2227c8571913d689a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I641539560711ff1824bd90baa0f21f96  <= 1'b0;
            Ib29b00328971c3cd67209a5ea5b63b0a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3ac0799861144b599995318bdade2114  <= 1'b0;
            I517e0868f2bb9a22c287a1f3eeaad2f3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie83fa8157a7cce44c2e25f46ce897dbb  <= 1'b0;
            I2bc9f76469e2a3f9846560ad1975cf54        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8be4711146486fea913843e497065b50  <= 1'b0;
            I9f089315e435cd69d2929fdd936a8a77        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I65171c9ee8449407484e5c82d13c6751  <= 1'b0;
            I9b54c9fb4179423c731217286e329930        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7353ebf3a1cde89d2bb3fa667f7f5485  <= 1'b0;
            I82fb41ab743146badfd2e82258afb310        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I669d34b955d2991ebbb31c149ad1b6f8  <= 1'b0;
            I5619b91de99eead78befdcba1c62411e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iabb01dc9980b4879a7356712b51df0d6  <= 1'b0;
            I83dd2047dece99cd841b2e7955819d57        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I373841aa2bcbad8232d54ac9035a3ef9  <= 1'b0;
            I8c927e66ccbf4d19f07af5ef9fbfe3fb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib6124faff821158c6a2c9a9c454ab68c  <= 1'b0;
            sum0_00048                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0793fa8938acdf65486e5582d01b9e5a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6f7a45fe64ffeda9ed120be3a4519aea  <= 1'b0;
            Ied68d7ba0ee9974eb33767e737760b4d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id1dafb7e45b860d506e0c2c91b28142e  <= 1'b0;
            I95ba37056659b29fd4318a68d85445e8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5f1609647f1e71cef4ba2d605c6c8445  <= 1'b0;
            I08d7051a18f358d08728f1c401c15c47        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If17c0096ce34b88007247bf4c429d5c4  <= 1'b0;
            I768b6f55827ac49eb6ac2655e9397be1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifc2963762403a00c4f3662b2863c991e  <= 1'b0;
            Ic66f737fe60c55d4c10e5d72b307a061        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5fdd8e1550feaecd81b82069fe73ed7e  <= 1'b0;
            I5653779f15c6c9b0f3b26927c48d6234        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I85654bd3a07b4329aba17d8b27777f4e  <= 1'b0;
            Iac550729fc437fd67151fab57134ec88        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibf2a253afde05c905d0b2404c5a808a0  <= 1'b0;
            I853b03c5826eedc3c67a2fae7a640212        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3ade5535a79ce83857481ac771cd8618  <= 1'b0;
            sum0_00049                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If46a6b47c1c52243cc0bc92d1edb594f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I221524a69e18854f029cad30e8f94e8a  <= 1'b0;
            I75b36a9b429cd657afc8151b9613aca6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied764ee7730ad129b6f62837ef50774a  <= 1'b0;
            Ife682dd9f677da4d27294fb61b141948        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic98f33c6a4613534bcc9b6bc4b4f2d17  <= 1'b0;
            Ic2b6177a9c586b274b68b25584e6df2c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I92eb6f60c14ee9eecb01718b01ea980f  <= 1'b0;
            I0d23011c4381496a19cced7bf7960546        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I97e82e5f6775d1e31537b891597223bd  <= 1'b0;
            Ic5992d5eaeafd5dded641a7d9801e763        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iba1c0ebd9cefeb0dd7f690bdbbbfec58  <= 1'b0;
            Ic9e7fe68b9045c6c9eb86185b5f5872e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I235c3a9fd3e8ea1cee762c10bc8e2c53  <= 1'b0;
            I51ad746720b5e6e09ab50f0283552f1a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idd474d80b50992537d6f527faf279800  <= 1'b0;
            I0c8964888a1315507f5d71959dd24cf0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I88a89b2d938552458dab9bc34728959b  <= 1'b0;
            sum0_00050                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id4d4f814a0bb3418cbf70c306acf048f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib105151d91678f81978495ff94b1e651  <= 1'b0;
            Ic91bd7b4bd148e526ca21d4a5ba87be9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4edd64d1f1da865b1eb886e22726a033  <= 1'b0;
            I7959dddc32f0f181b3ba39149afe1016        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia7c9c24f8e993526e76c6915e56908c4  <= 1'b0;
            I087263600b5f38be072a4f1db787aea7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib0dadebad37d9ea9d01350054872863c  <= 1'b0;
            I78d17a56de5cbe08191ef23b9731c485        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I76fd9005abd511c3c5bf6c77de8bf2f3  <= 1'b0;
            I82f713a43596df3b935d6da6f8041dc2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic124975d36a292816146a2fe61ab3ab9  <= 1'b0;
            I422987396853a6a39dabb6e7ddbf91fb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I70a4926e9e6a05fa9ee51a26988862fe  <= 1'b0;
            Ibb6556671e104141dd33188ea5fc024d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc5e98f6958786ccf95d39b922b42ea9  <= 1'b0;
            Ie42ce76076a2a5e887e0112086012da6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8879df010bbdf6e5fc9370e2fb3289b4  <= 1'b0;
            sum0_00051                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4aea430599b9c0702b3bebd5960b5c91        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I94a9de743d5bedbea3876de954f479bd  <= 1'b0;
            Icbe11a3970136e485eee1bc5053e7273        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17c9d8f658dd6b2916b645d103f4702a  <= 1'b0;
            I0a7f1ea1719c1f5ff104445a4130a5a8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I384e50fa8daa639124f083dda56fac00  <= 1'b0;
            I1802d759f26dd919bc315bfd4156238d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie165d0729542c81ca89f45d15e0afd3d  <= 1'b0;
            I2148493e253783fad70f4f2807b83008        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie8e29053f122a9247b0dec291c6ef4f3  <= 1'b0;
            I39e7f78d33aa7f50264908d2efe23634        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I453dd7d7c0a2f003f0b67e909630d641  <= 1'b0;
            I844be5874def16af98de935019f35fe8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5707d30ca29842b6a96cfaeb44ac6668  <= 1'b0;
            Iee5172ba70a6e368b4903f9ff1d93471        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3fbd40faa4c3b78b547b8348c466fd1f  <= 1'b0;
            I1f34b473283291e0970879465c005e2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9a403c511fe2d44472ab319a9477199c  <= 1'b0;
            sum0_00052                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie1e0b5120737a7f4bf845618ccd22239        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9db50007841762c9a10f6b7e9d40f858  <= 1'b0;
            I8abec3020ee5358f8768e5595e9992b4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I89c5af1a6176cefa1f77ee69996473cb  <= 1'b0;
            I6fe683073211a484cb6e3c416b365d9f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5ede62333e0f7ddc5446b653ba9a2382  <= 1'b0;
            Id7d764da58ade36853e8a45b5ee19dc3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I69d82ab774d52c219509e993e7cc4deb  <= 1'b0;
            I3cee2fdf353643deac7d6bca20c8fb52        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0eaa22f5eca8f33dd254fe241017a098  <= 1'b0;
            Ie9b8f8f0434fe3783c3d8f68fef30e50        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I570c036d0237c53bb069c52d621e539e  <= 1'b0;
            I68cba8ad7742cbb34d0b1fb16be4a58a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9d7614d286377329eb3999213889b707  <= 1'b0;
            Idcea56657d40e0fdf9a1c2d920938fd6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3eab1582cc42db0ac7739386cce2a712  <= 1'b0;
            Ic549ffab8f0ce161a177faa2ffd1326d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie4827dc0983c1a63053c08de6e36d375  <= 1'b0;
            I4d463d500f93f74b2724972ec1d62439        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2eed3d32a27d51036e17c4a21382b4c1  <= 1'b0;
            Iba2f362e263953331649c726afa9c481        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie039ab562e9cf90289047b5425186123  <= 1'b0;
            I6a053d931fb030e03d4882856d3bda75        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iefbdf686d9452a62cb99cf023a4d9fe7  <= 1'b0;
            sum0_00053                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I27ede93004e0c240efaa56cc8c570910        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc5dd6caa4ed17a63746d30d381a944e  <= 1'b0;
            I61a11c1711ca10eefea3438722b40bff        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17086dc5193aa55e5c6f56ecd365cc00  <= 1'b0;
            Ia7924c88692cfddf24fb1eff66eacb7e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib2fe0f68044c11f879e512a200f8099e  <= 1'b0;
            Ibcfd01e622f7f5a5156dd9b335b4e5e0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I768720af835b02a8dab376ef23d17a15  <= 1'b0;
            I7f6f418ea51b4298da8758bda3f6a21b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1d98943b01a6a2d8c4db18b98dd62f5c  <= 1'b0;
            I7185da8937449e23abdd0f39a4b3ed7d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id3b089fb6edd5bcfdbca142fddd5ff89  <= 1'b0;
            Idc3e3ffa31d9b76c7cf9358a5b2e65d7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5196382b75d16892d550f17893de15ec  <= 1'b0;
            I31fe8c887c4aff7c69336676cd31aaa1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6387919f2426c283e2d70e471cda54a6  <= 1'b0;
            I59684d5fe6bbb4b54ac097bd25fceef5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3b84dad6d0dd8730312b3e20c6d5a2a8  <= 1'b0;
            I86a7cd69148f9590ce91d0aa270d6c54        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2a4bbedf880a9a7b4e1bf946f9f96c0e  <= 1'b0;
            Iabce1ccdd968980f622f0e137b159d11        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I49d35ec6369de10afb15be8e0cf135c3  <= 1'b0;
            Iff02977d7b4c733cca1794246f630931        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic3ba4531855366e9a060cec1c7694844  <= 1'b0;
            sum0_00054                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9026c904e5ead7ff2994c4f781d61466        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4dbabfd592b74aef93b819163130ef5e  <= 1'b0;
            I99d7489ba87c629c6dd9702a9bbfd3c8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9ece87047aec25abc02a5eea72f0e647  <= 1'b0;
            Ifaf191e0d00ba6da7019c2efcf08e1d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3ed6426fbdba8aaf1c948cca7442b3a6  <= 1'b0;
            I4c295991fb08c90862a2f3ba6489000a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I24075f37c6bbd90c83370de1a2e58af2  <= 1'b0;
            Iee61d179da125934298400256788cbb8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3175159add7b814df637c2db8feb43f6  <= 1'b0;
            If87c84440426fb24070372dc1d4bf315        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0a569f6536789efb7ad2377c11842830  <= 1'b0;
            Ib9259a807b31c1b7a528d336bfc403ee        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iae6ed7748692f2edf1aa9d73380075f0  <= 1'b0;
            I411c4d909b2a571e685cd703245516d7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib4ae1cedd09d72c235765a6cd7e91366  <= 1'b0;
            If8425453cca8fc8623cb85375c4b8a1d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie2d946edaddd3c87f328e861f3e72c0a  <= 1'b0;
            I654b497f62df75fa283127b5de29b1ad        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id6b508145cd21ba088ab8fda34577c35  <= 1'b0;
            I2768519342f7b8a1ee40c1d5ac502b66        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifa6e3541f5e12bf9677ffc51d0392749  <= 1'b0;
            I8e354c1c5ba44fe5430887248ce0c43b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I21e72a7e5870151c3247d15121e5fb4f  <= 1'b0;
            sum0_00055                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8970d8a8aea29913e8696c14c153d16e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iba283e99a57d0a3b78ad2e309c316b65  <= 1'b0;
            I3555c6e2fd480a6be11549bf95a9b0b1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifba3e46933049cb093d2c1809f3a8a3e  <= 1'b0;
            I8d5600a352e8ba4756f917f912fda6dd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4af3e2bf2ebc913ac902b48da672c5b6  <= 1'b0;
            I7e99d73c95e7ae5c3fe07a3c60ef52eb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifbadefd3a7ab50719a703400ddd742c6  <= 1'b0;
            I831633aebe5c6a52b98d630205376f3a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If2042aede3390bd208a281f0380c95a4  <= 1'b0;
            I82e35482de74223be0d2558334ac2dfb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I19b73c5c93a71e90f620572f23f0e6d2  <= 1'b0;
            Iae2a6f9649ef1bb193e4f0ab5ecbc3e3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4b99891bed4f5c149cd4a5b4f1dde0f0  <= 1'b0;
            Ie8eca65d791ad2f6e8f4ed244f22ae3d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3472ee8c06644490252e606b62bf9bd5  <= 1'b0;
            Ic24146b01094df9b9ccd455a791f239d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idb1efe99b5d7fd567a7f82cfd52f7eb8  <= 1'b0;
            I1c9031fd54ff9417d44c9fb17dc1fc63        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I24f82a3f2c0e8df486fe495dd95cf8bc  <= 1'b0;
            Idefa20487bc5ba6daff03e6b327d76c6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I83ecf12f3b38fc14c3b75e47b71ecc09  <= 1'b0;
            I6f984fd9ea27b40ab3afeac8afd29ade        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I74cbc0ec3bb682e0f927890eef8d7a58  <= 1'b0;
            sum0_00056                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0be92debced4961df5f461fe81e80bf1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I989dda9add29306d7b3c0f376822763a  <= 1'b0;
            sum0_00057                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia7bdaba4c6601b7146498aea6c9a3e07        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibc929201e2eeb3e61cc8f0acbade497a  <= 1'b0;
            sum0_00058                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id450c0a1cabe087be051fbf4158e6016        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib0dfbbbca2d3d264065f73b4241caed5  <= 1'b0;
            sum0_00059                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I656d0d69f6e243746b87ad67764dbc3d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I339786aa60d4c71d12c65db27ac420fe  <= 1'b0;
            sum0_00060                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iab9d870dc1ad159bbaecb20a9b72f005        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3ade020bbdf8f954821f737439513043  <= 1'b0;
            sum0_00061                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id53b60854f19e095c38f2c255dc57f29        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia50526cd3a3174bebc5a7a0889fda661  <= 1'b0;
            sum0_00062                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If9ba44a2e4a8f0b61692fc69ebeb82bd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie9f37dba0791359bc426a73639ce33ad  <= 1'b0;
            sum0_00063                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ief95e8620a1c8ddfd6df673a3a223bd8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9518532a8617fc8290eb6a5e981dea94  <= 1'b0;
            sum0_00064                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I61519bc0aa02ed461dbb91851d0ae19e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If66524125bfde5aa48ac70c4e448b38f  <= 1'b0;
            sum0_00065                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie0c11d584811174a66ca221baf87c36b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic3ec6375998b05a3e48f6c5fe7b3910b  <= 1'b0;
            sum0_00066                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If10f4f45ff0fd17541735934ad20f187        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0ac421af6e311b6005c3e02e93ff94ce  <= 1'b0;
            sum0_00067                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I445919f07a6fa8654211301a9a6126bd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib9db80f43718305a8a8774d8d80c86c9  <= 1'b0;
            sum0_00068                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I64102b82893352549abd2e2132b19476        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3b775b06b5d78fcd7373c966a62f44ad  <= 1'b0;
            sum0_00069                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I1fc1933fe891ac26f35a42a1b242d919        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If2372a5956f21f97eeb9c76281b6675e  <= 1'b0;
            sum0_00070                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I84dfba8bcf8ad3b85f9472fd60d607b5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7b32c2b108e24750e2a24785668af3ea  <= 1'b0;
            sum0_00071                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4302fccefe5ee13161f9ad49f9ddf43c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8ec99197a7d823f5745d382c10161430  <= 1'b0;
            sum0_00072                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I59d7153724d3b3805af799692fbe245a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib895fec0b3756932b85962c1d129a03e  <= 1'b0;
            sum0_00073                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id1650d0e39be078027493f58e9bbcbdd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I76aab345d13c6678fe37a4a7133cfd7d  <= 1'b0;
            sum0_00074                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If40ad4aca8dbb3bf7dde8c2ff2e5b8f2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib4f368fa3d3ec11d9ffb2ae9a2ae6310  <= 1'b0;
            sum0_00075                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie49f173549396caeab1d13da36e37c65        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idd0f3cfc5599481c954a2bfe69f044e5  <= 1'b0;
            sum0_00076                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I3002a0e0cdf8e79bc7186a876410d106        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie624c4dad5036a25ca314b94cf3c4b95  <= 1'b0;
            sum0_00077                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2b50fa03f584d10e9af3be085a02a12c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibf4b3caa5655cfb6663f9b7e2383bbbf  <= 1'b0;
            sum0_00078                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If473d172a7bff5aeae99245bbb72978d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I049d1c09c15def12ba7bae95fc1c3d55  <= 1'b0;
            sum0_00079                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ib89f7b5625995290a64bcfb143d978ca        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ide06ba186ddb179b489ba6e3e209e3e8  <= 1'b0;
            sum0_00080                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iebe0c9b4a87d58a1c55e2ee6b01603c4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1b78785ebe2e7f77a3125a6334c4dc54  <= 1'b0;
            sum0_00081                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I104411bb641d2445c7e1385a809bb682        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie79c93f1703121713fb9401617f349a8  <= 1'b0;
            sum0_00082                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I47dd28b4ae4f7151aff5bb271e35b716        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icf25f076eec2bf81c899c66f6cfbebc0  <= 1'b0;
            sum0_00083                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I3a27d5573b748df459b90a5a347f9d09        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic5c837a0556d1cb66edbf0294d08283a  <= 1'b0;
            sum0_00084                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2dbef85d2b2b95af39c3a98c4e143253        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I51ff4bda38746682e3cd4c68118c3216  <= 1'b0;
            sum0_00085                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I510d39830ae7b0a857ac11baa7c144d3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1c074a53e6c0f2467bcdd7c952f51670  <= 1'b0;
            sum0_00086                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2751a94a66ea4cb44c512df4c509937f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I37c49c5a2af240496f5a5706b0d42ea6  <= 1'b0;
            sum0_00087                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic9a003bfb70ac2da6c229fcad09246d4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia94c439131e1df5c95fc8ad3cfdba473  <= 1'b0;
            sum0_00088                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I34ed986182a3311a8cb005b3dccc224b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I723a6fee3b2496f23c48b3584f8bf9ce  <= 1'b0;
            sum0_00089                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic79281755397f6099ff30c5d07d7e6de        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I648b62fa0bc2185c1756ee531e8e34de  <= 1'b0;
            sum0_00090                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8d6559ccc33cbc663584923a55b928b5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ife631f9a3c4c64a3d92aa9586ae75f3c  <= 1'b0;
            sum0_00091                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4f0a4c241844e390318f11899a0f2c5a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaac1d82f0846fce1bd88ebf8e60300ac  <= 1'b0;
            sum0_00092                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I45fffa266ce3838f82d755b59216a4d6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I48cd09f035f668536cd288a23010b07b  <= 1'b0;
            sum0_00093                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8f0e65f5db47d5460d4ec2172807a3e1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I119b2e5c2fea5338244c4019884af26f  <= 1'b0;
            sum0_00094                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I34127c0d1af2438e13b6f4709ece80ba        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2bd34b2fd12f12bc301fd0d5d69c0fb6  <= 1'b0;
            sum0_00095                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I3a67de0e76bbf29d8c77c21865abda2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib715b1e0061b84ce614a30d961a83e7e  <= 1'b0;
            sum0_00096                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic64e64aeb754249b868e14311ea19759        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ief8c2838abac83370fd7ec25c06d509b  <= 1'b0;
            sum0_00097                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic4aa0dc9014c8445f8d9a7723d7263f5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I561d79eb079915c0b1732cbddb119c2d  <= 1'b0;
            sum0_00098                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I47b988d017580bdfe8f443904b1f3aac        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8bb75bf828d5ef337fa6a965808e4638  <= 1'b0;
            sum0_00099                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ica9ff13e8c3850be6c70b0b06c1d9fbf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I11ba339c8250d07b497c88a39a6df1ac  <= 1'b0;
            sum0_00100                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If2efeb489911f295dd7722cb22ea521d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I173aa69cf52114e223ac1410d90b4bfe  <= 1'b0;
            sum0_00101                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iaa16dffcc01e41e6ff17e92bdefe3df5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia4e89e99acb95f4183474b94798ca35d  <= 1'b0;
            sum0_00102                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie8857b9841fbd795a4192976ef7ecc25        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If4c36727ab1c29bf78f72e8acfc00d7c  <= 1'b0;
            sum0_00103                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If12aef69eea28052aa3bdb6ac31af205        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6426943b4ab66f17c2b7b399ccc7a6a9  <= 1'b0;
            sum0_00104                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0b3c6162ae2b9221738a18a29489887f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddcffa815489773b3688fd68dba18bd8  <= 1'b0;
            sum0_00105                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I08211bba29e87faf4079152bcc973e7d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id00642563679fa9a6696f8e7bbdf6576  <= 1'b0;
            sum0_00106                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ibff3da265f1c3f21548f5b019e1a9dc1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifda1c55899cd3506853cc82b450b3936  <= 1'b0;
            sum0_00107                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie9fa1762d7844b0d781afdfb0771cea9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib5d1a7cdbcba0b654c12063d4f1768e1  <= 1'b0;
            sum0_00108                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia677d504b9f7fc2698c0345f236428ba        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5e8ed024e2f2548bb375a2ecf1918a5f  <= 1'b0;
            sum0_00109                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Idebce29121c0481df83d755b60ff632c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id25deba967318f049de8163e67262f4b  <= 1'b0;
            sum0_00110                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iad2c780a6386674d50cca54d8c4ebd86        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I925f6b549a25cdc8f85152eb21ea3b58  <= 1'b0;
            sum0_00111                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If1d7944e7c4828ddb91ffea28609cbc7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9b49e1acb81ef5b088b808d2e4ce9954  <= 1'b0;
            sum0_00112                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I843a68ceb0adab829091f31d0de56eb6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6386a4dd26e7c36165dc265b3a2c93cf  <= 1'b0;
            sum0_00113                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I59701b9eb54dda2744a79cebe7d73f3b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia20709f08cfff3a51d4af1e81d640400  <= 1'b0;
            sum0_00114                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If63cf5e8f47e4e51176401f0d954ea23        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1ff042bdb52aac5d69791e96e2f9706c  <= 1'b0;
            sum0_00115                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id09454844b525697de3e3727d89551e4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaa2cbf59f6f61198b4fcf5a741cd5bc8  <= 1'b0;
            sum0_00116                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6d1b2ce4368945b56eee7814638471cc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I01c94743a11042e75638ba6618356203  <= 1'b0;
            sum0_00117                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6079945faa57335b1c902ccf7f960a70        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0a0340a0e52145f3597accfe4a4e8624  <= 1'b0;
            sum0_00118                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie7752906ac55cf51f3e96e8c0046f1aa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3bb4d24caaa0882a75125e466070f0b1  <= 1'b0;
            sum0_00119                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2d7d4135a94f5df949283c043228791f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I44ead0ab5ccc53226fccc03024643771  <= 1'b0;
            sum0_00120                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I99c75e3d26c5d01f6ae9abcd05407d8c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaded125f7fd5c833e7206dd7071069be  <= 1'b0;
            sum0_00121                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I81e6f97621dbfb2fed6fc236005a2b19        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I373be7c3f9511a2906584e33e5048abf  <= 1'b0;
            sum0_00122                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ieac60532dcfc916a65054e35cf31d6d2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie0b5f51835ebdb508a596eeebf0e4847  <= 1'b0;
            sum0_00123                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ib7eb83ba73e0dc17f69c357b6ca555bf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddb75e0197b9a76b36a59ac2a7ccdf3a  <= 1'b0;
            sum0_00124                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I5139d8a7a099e3c619c60647c15b7420        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I08c03198b9599b2f4590e3022e398f7c  <= 1'b0;
            sum0_00125                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6ccd2e11ebd5b2de80b120e20650a602        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia4f3cff223e24815ee1d86bf41756f06  <= 1'b0;
            sum0_00126                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie669cebe5fe39e1a841f8dd3c1f6bc57        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I56592e1452c4b559af19465b30230ec0  <= 1'b0;
            sum0_00127                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If32acb9fc212c4af34099acf6df2bc5a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I213ce488e5345fa405a9c5df297d6f74  <= 1'b0;
            sum0_00128                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I075ce236a181bf925c8ccce91d9bc8cd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iefac1e428116a797c2c0803410ac5601  <= 1'b0;
            sum0_00129                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I541d4e422b999a0dfca44d275178e1d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8b419d5827e5b1af9649d602401c189a  <= 1'b0;
            sum0_00130                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I3e02657f3d9f79338cd083ed024bf96c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie989550c9101de382056dd60d5da0e01  <= 1'b0;
            sum0_00131                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia5e5537405ab8edcc7cd43c86837d43d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I259010e323e1e8dcd9dd719091131f6c  <= 1'b0;
            sum0_00132                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I07ff388e3b6c7288f0f6c35a345023fe        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I389ac86954fd70464c9550e3fed4ed33  <= 1'b0;
            sum0_00133                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I56cb3b3e193ca5068734417fd0ec4e02        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I77371f0e55b4684d1af196ed52d3d997  <= 1'b0;
            sum0_00134                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I5bbf1765d8f81581d0cf31c0bc755fb3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5a21996f5724a2a49fcf8e928c01b062  <= 1'b0;
            sum0_00135                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iaa1643095e518846cdede4d5a90dff84        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id46108963921efa50aff64d4dd7d1701  <= 1'b0;
            sum0_00136                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iee6e12f4717a3279dd31b874eabae69e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8da50e5093acefb6f809aed64564a53e  <= 1'b0;
            sum0_00137                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic52a9edbbc5283844d2514ea142ca6e2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I03b0694777d0160a83cbc82ac1397736  <= 1'b0;
            sum0_00138                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ice3e978c8da2a7de5b28542a5589f0a2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I85c2bffb93569d9fe1b1bcb10b98bcac  <= 1'b0;
            sum0_00139                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I336a425aed221c85ca80b9a97d21d6b1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id00274c88b93867a80606343add1cdab  <= 1'b0;
            sum0_00140                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie477c0f3b77bb299ba8b1a410d211ef7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I61e829cbf7d6c0ef8ddc11677981e2cf  <= 1'b0;
            sum0_00141                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie62920d089ae762603cd33fbf97d92bb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9e8ae2aed048068b01b3bd46f30baae8  <= 1'b0;
            sum0_00142                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2ca952e4e676537fd5a8fc71ecfa10e9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7dab71adbe62687846fc027d2789451d  <= 1'b0;
            sum0_00143                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iefd31e7ff3c829c88f60bc89d70afcf7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If1295608bd218ed60922a0b95bf1d098  <= 1'b0;
            sum0_00144                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iafa987a413fd8fcacfe872bc0f5bc2d6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idf04e08c120ed116af14a62659675b44  <= 1'b0;
            sum0_00145                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I305c1ea420d666f258e38c5a65847367        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ieb7614ad1b1bfed3e2b0089a72fe214a  <= 1'b0;
            sum0_00146                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9f040c4088bfab72d74e5332e9710d1a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I589062eca318b25dfe5735da455b6fe1  <= 1'b0;
            sum0_00147                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia2f41f9778324a06daeb185c736516a4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If3db87afb3ea184c9e4020c5e45cb161  <= 1'b0;
            sum0_00148                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id9778ba5fbdbed4d33a092da6b68c414        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia14bc1fcd5bbdcb60b8e68298f7d716a  <= 1'b0;
            sum0_00149                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I27c2c79d0d719c71c8e28218d1174a13        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I268b60cb371b3d46dc3f8b0009f541b1  <= 1'b0;
            sum0_00150                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2a9d6a774769b12ae20bc0cee0c36f5c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If2cd93b57cd1c2b91ee7a73a97dd19f2  <= 1'b0;
            sum0_00151                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2c567b75f1399c069b95284f4c36b6d1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id81305359a07db527e49fda05cd2784f  <= 1'b0;
            sum0_00152                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If3d3eb609abfd6e315eec803d2e94490        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id8292eca087c1a17dc8b5a572a76f21f  <= 1'b0;
            sum0_00153                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9c58aea7ce986b1d28f5808b347c015d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddb19725b093506e5e521d8d68dcb8e1  <= 1'b0;
            sum0_00154                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id139c7a783196941100003b6cb0cd1e7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0b573d3a86a3111451da661e46384876  <= 1'b0;
            sum0_00155                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I524d7614b01460778da3ce98f6aaa3d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0ff479e61d1a0cede88ebffb073c60be  <= 1'b0;
            sum0_00156                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8acda65f116d5c91cbe2662ac282aa31        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icd6f8f5df6b4ca4c81855e974db76526  <= 1'b0;
            sum0_00157                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If67dbe22f8d22b3430215fb0deae8204        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7ce064a756dad56d37684d5d7d168047  <= 1'b0;
            sum0_00158                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9a35cd7512787263abedd6d9913cf507        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied2ea62cfb21602645babc36e27b8218  <= 1'b0;
            sum0_00159                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If9cca23469c5e6001650f1f8b1360ae8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I79b85da6e5ce0b02ebd1619115c98e24  <= 1'b0;
            sum0_00160                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Icc2606ae8f9a3b425225ae7339112b9d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8e1ddd7e4185c28caa71d30bc28138f3  <= 1'b0;
            sum0_00161                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I34aa1802d24e074ae54563898929abfa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iab0bff1633e2f3ea0bfbc291f3ab5d29  <= 1'b0;
            sum0_00162                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Icb85b3464dc40e8504c53c377e889c45        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5f0751fceaa008feba5c6867ced453dc  <= 1'b0;
            sum0_00163                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie595a7d10b5ac84c0301fb55bebd3680        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9f6751c15237c20b0cf2175575195ea7  <= 1'b0;
            sum0_00164                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9c217a672cabc05efbdff218637123ba        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6ea50be10bc990a1206cdc9e28e0c4c2  <= 1'b0;
            sum0_00165                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If20f3780b4af857ffe8083056085517a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I43c2fab87f70ea883321ab82de85f133  <= 1'b0;
            sum0_00166                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic2e275bfa8ab3d2002d2aa374ac9bfe2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1af02ed6cf00d4cb0704b5e44c83bfa3  <= 1'b0;
            sum0_00167                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iac5798fd9915b6778700da6a14f6a381        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib71611afdd0381cc1884f5ddbbae1acc  <= 1'b0;
            sum0_00168                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ide3204bf317fdfb993410d338085b174        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I38fc49afce0298846ae8ed63ae715e81  <= 1'b0;
            sum0_00169                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic3a95140fc1029efa17a6557bc977719        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddc3e44d83e8253e5129b6cbf5082df7  <= 1'b0;
            sum0_00170                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I647d3a46bb2c7ed0f1ec08760b3858be        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I975a87bdda30c5b6be8d2f0e4b107450  <= 1'b0;
            sum0_00171                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4816747af9d9fc8dc85fd831336ec710        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I582bd96afa764ded148202f738b7a1df  <= 1'b0;
            sum0_00172                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I1f66c026a5437320bd1f4df2ff71663d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6fb88d97bc9ed37a06b729020a1df140  <= 1'b0;
            sum0_00173                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If347c58c328193f420286ea27a4afa20        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1500943c4a550e78fc169437b0a663b7  <= 1'b0;
            sum0_00174                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I7a126c8304be920f2a920315dc61ba7f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0b83f4ef8ba9badb27e81b32765ec5b6  <= 1'b0;
            sum0_00175                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I237327d6a74df1fb05537dc3691ebf11        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2c420acf428e44cdd9ca9998e276f258  <= 1'b0;
            sum0_00176                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I64a3e8bb4c87b066806d33a5306a2c53        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic7b6dae3017b55dd3cd27423d5f1b0ec  <= 1'b0;
            sum0_00177                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ibbca6ec39234473fb517447a8beacafc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4a91a7c9b2a0f3552b8f2ef4e2398be2  <= 1'b0;
            sum0_00178                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I78327356176a16fc996188b83b058cbc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I99ff29c7ba68b5d0819f1e1bead51287  <= 1'b0;
            sum0_00179                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ifec496c87a7a2474855067305ac8cba3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If06b00be0356a2be5074d958ddcdb2f9  <= 1'b0;
            sum0_00180                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I41584165a62caaa37ddebbf79bb8b617        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I604283449f13c7b225ea03f99f2e296a  <= 1'b0;
            sum0_00181                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Idf0916d6b025aad6eccb98ada5ba3aca        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2b600e5f5c146ee97c4044c08e1f5ad5  <= 1'b0;
            sum0_00182                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I00ef133d5a53f8f99f35b50327e5272b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9fe16403fc21bb1159a5e0305fd1ef69  <= 1'b0;
            sum0_00183                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6f0e302d38d75982d0761e306ce9f146        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iabdb9374e5caee281c25b003624b2c4e  <= 1'b0;
            sum0_00184                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I127eed5de00e10a020717e796de76c7d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibd12036702fe60b57354b3aac921559d  <= 1'b0;
            sum0_00185                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If9aad73aefb1b225f35e8c813b85fe87        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib1639811de6eb1c38257800c201fb704  <= 1'b0;
            sum0_00186                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I00a89ac37676521a081a21b1ec1a0798        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If926d98f659e8fe4bbf36ad2c5c852c5  <= 1'b0;
            sum0_00187                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I06f3a34f2b1770ef82ddc2a732b3d4fb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I211f8d7f97ebb8eb3e50313513abfb1b  <= 1'b0;
            sum0_00188                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4744d64a746f16004e3bedaaa41465f1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I304ac9f96945546cdf1b6f1fa7136731  <= 1'b0;
            sum0_00189                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ifae0cc6cc1c65d24bbe84c4ba938e2ea        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7a9800418bd5c195fc47a72370680b56  <= 1'b0;
            sum0_00190                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I1223c21129382d41e4f38ef4bbe60c2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5f6a61c9f0c67510e148e596f553a4d6  <= 1'b0;
            sum0_00191                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I14e36e16df00adcd7dc1973d3852d2d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8e313ceb21359bcc44114ab217b1c394  <= 1'b0;
            sum0_00192                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0d05ae27b53fb6939e4c2f862a8d20b2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4c9518755c33d725221ad79ee6badba9  <= 1'b0;
            sum0_00193                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I97a6fcc08929c3b7d15e36d7706ed13d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3c3cffec9f47c9979cb9503f222f370c  <= 1'b0;
            sum0_00194                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I1f04e86bf27596718836d0a09adbe120        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I68d6769541fdc3df321e192f645c667f  <= 1'b0;
            sum0_00195                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie40873cfd6d10a61a94a761becf588a8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ided55428cbb77f454c2607ac783d7548  <= 1'b0;
            sum0_00196                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I61960ed74fee948cc12bd1fd8384559a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifd3d4f3e2a388b3c70e7704d6351e0ba  <= 1'b0;
            sum0_00197                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8533a3ec4be4c49166184c94761eaebc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17d32f292758416fe02527dfd938fa0d  <= 1'b0;
            sum0_00198                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I00be319b5bdb85ffaf3bb0eca0b348b6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9ce3942aba354c1fd7d6b9a39c994d7b  <= 1'b0;
            sum0_00199                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie889c916b5af185b52ff5e2e3cc23045        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2c6c6041c9c69c84f4d64af6458955f5  <= 1'b0;
            sum0_00200                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I89697be6dcb2e7f972db498c1b1dea71        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I830a4fffe1244e071eb82c28ddc4a308  <= 1'b0;
            sum0_00201                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If13dfbfff7cd8e197bb44006a3db73bf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifad8e46fc3844bbfaf434a14f6b5869d  <= 1'b0;
            sum0_00202                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I87ed6c3e172c7a06bf6aefe7bf718d70        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I10a6c6a8fdb0003de1f360c148777d0f  <= 1'b0;
            sum0_00203                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0db87adc849839fab3a4c9884d5a4882        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4cde586fc28f8d03fc9934d56f7ff7b8  <= 1'b0;
            sum0_00204                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I535e01a6c35fd7b455e4b79b1d4bb414        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib83a067fb08e118dcf794902beef9405  <= 1'b0;
            sum0_00205                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia2d1c752cc4b405adb97a815e90a7b96        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I358cf9609272a4562423a85f9b2f56bf  <= 1'b0;
            sum0_00206                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9ac12eb3878f6fc7dc428fe5e7f35d97        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic1e9d9113150ad57954c0e369259dc62  <= 1'b0;
            sum0_00207                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If46fa11dfadb0691eaaa0a40836e08d8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If7fe3f5ccbb5b279e41fd183c8ff3974  <= 1'b0;
       end else begin
           if (start_dec || start_d6) begin //d7 for Id0cab90d8d20d57e2f2b9be52f7dd25d I37302ccecb8ae11c64170bc6bfa44eaa sum
               sum0_00000  <=
                      (Iea07d1adf9016a29cffd61d183e268d0) +
                      (If92db65b39a83e1c699e4cc6d7f9e57b) +
                      (I8f2986bc015fcc64ac5e5395ac6dd851) +
                      (I355725a804e0df68b4acf96ca98f2448) +
                      (I78212ae965ab2dcb2eed0b060d6b253f) +
                      (I0b56aa7a1b7549c91dddd3a06ecbaacf) +
                      (I71412803cc5229025487255aec62ec4f) +
                      (I32fcb28a27356bc6f403528836ea4c1f) +
                      (Iad354d876cb9fc72fc0143e6f7da9357) +
                      (If6e745bb85abba7282dae1f6f701225e) +
                      (I93bb43c1b89d4c70a57bdc019d64fd22) +
                      (I7a2e554d07bbea291f2cfc18694fca3a) +
                      (I3e59b2419c7dd1553b792d536208514e) +
                      (I46894c6526983bf1ce4b503159131b41) +
                      (I6404d0df952b5bf8292c753e4c6f35d8) +
                      (I8522c402e654d007abffcb0e904af5e6) +
                      (I5ed85845c39337c37791f16e718069b4) +
                      (I89013d61c1ea8da8b1c6071cc21c316f) +
                      (I4102100fa5f1dd299af0190862efcc42) +
                      (I4939f69abb1eac56d5021e06406a93b5) +
                      (Iadbd245bf842aebb456417579a3e6296) +
                      (Ifc8ece44a4e68c3117eda9e65f3084d2) +
                      (({q0_1[0],q0_0[0]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[0],q0_0[0]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00001  <=
                      (I91679dfab57a372eddc7f9b94a231edb) +
                      (I2213c1a2b831f421707a261f5a58b1b1) +
                      (Ic53b875b2ddcba11406eb2ca39354757) +
                      (I634484f00590216c0f74f975c9c83400) +
                      (Ib3b1db2d8b669988c887ed780e439b26) +
                      (I735db8b0ee0ec98e4cce0030b11508da) +
                      (If1607e907e626902ee26d15020a64c21) +
                      (I081b38dbb37d4c14a6a9fd3fefa13daa) +
                      (Ibac5e7b6d4bf5cd6926358318f0c418f) +
                      (Iadfc60386481092ae85cc148a2c40abb) +
                      (Ie0ee5445c56a5f9b41640b57422206de) +
                      (Ie5f8620371236cb11c9e88c16b509ee8) +
                      (I8d7c1fe2e33bbd45379b0325a3c5e989) +
                      (I4fbdc4ee57a3be42b62d9bd43078d6ef) +
                      (I5510b88bfd65811b3200adf4ef975b48) +
                      (Ib57ef2f577cca54713c16717cbbd1ce9) +
                      (I15943aa74e9fbbaebdc0d54eb6a3bffa) +
                      (I6ac24c46319a787daa5c545de8c6eeea) +
                      (I52403a0454e5fa002e79eaab7ea497bd) +
                      (I634f0ce28934600a1a31ab0d8e59b4a9) +
                      (I7103aa739616a39c03e675ea0efb0335) +
                      (I0296d01fd3f9a269a617efd4beea9b8b) +
                      (({q0_1[1],q0_0[1]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[1],q0_0[1]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00002  <=
                      (I065a81ba25962785215583e7ece27661) +
                      (I631a3300cb6685f47da7781940ec5d27) +
                      (I8bbe1a2ace8f51aa22cca5d9fc66f136) +
                      (I38c3e3e136acb79c8a0ff850bcc55f16) +
                      (I35b2c7e9cdc53a98913e1c16a3a47b37) +
                      (Ib1a2b31d49ae476e2f1fb9acba2d5af0) +
                      (Ic72f41f9bbf470aee3c9b9b8787b31c3) +
                      (I3ea4c33a9419820ed54460eb64134dff) +
                      (Ia0d940e16c8cbd4f7544f5a5cd7d83b2) +
                      (I4a8abfa0896ce414d9b98093ef84455f) +
                      (I680be647bf2a62e0ee9b5d379dc87b4f) +
                      (If4d75f83299a21802b6fbe136913489f) +
                      (Ibddfda6413e3dd2f483c3174ea836b6a) +
                      (I33bddb0adcc2af7b12a83bf843036385) +
                      (I529f92b82248efe2cf64f7da0ec8283c) +
                      (I2f34af0036985cd94ade9cc905bec065) +
                      (Ia1a0d8d7dfd6e877f15cce773f85f5b7) +
                      (I5dd29fd1a73df5662d2b636e7285bad9) +
                      (Ide530e6f4622c8a7b101b6dce9650e42) +
                      (Ibaf00a6780325882067a79f0c4d693d2) +
                      (I16e3559c63ebfed83d6698fc9a9cd93a) +
                      (I9747a02384abb1c2dd1f52b3a5a999cc) +
                      (({q0_1[2],q0_0[2]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[2],q0_0[2]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00003  <=
                      (Iceb7a1d4c23806b8f5824016779ad129) +
                      (I40ef50004a60ae58aedc49eb5e6797c9) +
                      (I753f92da60980736440aba814a156f1e) +
                      (I4ac79b67a8904b95f7912d24af420585) +
                      (Iad44c932cfa5c249c5e59f8c706173a8) +
                      (I10f14b6433498e3b9e9bf021b60115e8) +
                      (I96008f47b9f134c9c4274cfcfb28e550) +
                      (Id0344146d1a53d418add6d2b185377dd) +
                      (I1eede74f12d37331b399eb7136bc621f) +
                      (I3e4754acc31d99bc71525789bdee0c1a) +
                      (I11c1fc94a3bd6dffa17e1571cc6ae97c) +
                      (I5395ee57418c31e11cf847f0f514ec19) +
                      (Iff125392fa39afebae1637a19c4e23ec) +
                      (Ia6308e16fae5428f4ab6560f5b21479a) +
                      (I5ea02b5349cd4d99ccbcb6b26f0cfdd7) +
                      (I21de4f6194dec9e3c401934db92c25e7) +
                      (I57d0920119f8901bd4dea2d5f8fb5d90) +
                      (I89537301987d6da0dbe6cff3caab3ff4) +
                      (Iaf0bbbe791bb71d0f557dc71caa5fb87) +
                      (Ic7ff9cde71054c1ee9eef81eabdd7061) +
                      (I88c10c47ae424fbdcb852fbf1e94127c) +
                      (Icd2e75e47cab1d539ba9ff1b6e1d7155) +
                      (({q0_1[3],q0_0[3]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[3],q0_0[3]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00004  <=
                      (I37e6bc7aff363ed0ed1f84b23c5f3e34) +
                      (I733605337bf6972630c089d32fd7f98f) +
                      (Idcb1d8bbdeaed6768c2a418c3048e6ee) +
                      (Ia89da2f1890524ad3519ab403dd0686c) +
                      (Ie33a780b0221084898c9fc5b237b244a) +
                      (Iabbd1668e0014df518ede5216232834c) +
                      (Ibd89458312687610aa166a9538968851) +
                      (Icbaf92a8e9875bcb19a1d074779a9ea5) +
                      (I80f3c8559da8e97bc5397bb8b621a0bd) +
                      (I7a0eada108891aba06cecab5071232c9) +
                      (Ie21a2c9b22e7bf8425fb5c0f33e5f4f7) +
                      (Iaa5b2807e5cc2403c5787eeb3d10ca6b) +
                      (I6da2b3a481ee71b85f3087b36b399288) +
                      (I11094e852295755925c3c61f1df81643) +
                      (I9c633aa620cca127b0ff8cf882178e76) +
                      (I694d471fd353eb54aae08a2afa7b645a) +
                      (I816704585ad393f685731104ad3ec64f) +
                      (I85d95015a9ce27a18ccbf73bbbcdbd70) +
                      (I992e7c551b4aa818606c3465d33eb798) +
                      (I2ead0e9941e2280309ab53535b1e1ac1) +
                      (I56873feb8418005b5661c7382f2dbeec) +
                      (Ib6ea4a822da2ea32e0abf6cf8a33d295) +
                      (Id1659ccdeaea3e59eb2d3f65a65ebd05) +
                      (({q0_1[4],q0_0[4]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[4],q0_0[4]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00005  <=
                      (Ic2171967791a0329f3e39fc19d0a6bc8) +
                      (I7d5041a6796c00188f74936d283defe6) +
                      (Iba7608ee0a01af103e022bcaf564bf6b) +
                      (Iedbe9d0e48bd36064f59faea51afddb9) +
                      (Ic3871325d57b310c95ca02fcaca529eb) +
                      (I42f9b1f8ef24ad56c10086852678b456) +
                      (I3ed5d0fca86f35b3d4b4a89c6147d0cd) +
                      (Ib0126fb335e32793c400a97c5a4a337c) +
                      (I20590d8fb97ec0b2164ffe17826136a7) +
                      (I3c128efc9f80c9b8334bf7b61de71b43) +
                      (Ic7147944f8835e26b9838fdbdc18ca41) +
                      (I698b1dbc9d8664d1c86c7a763d97b3b7) +
                      (I508bbade361787127e1a2e8687ec884c) +
                      (I2afeb2a7b199c0c6738938f156ae4274) +
                      (I86255756ddd1f88b74e070b19f8c3bfa) +
                      (I7d4924388dc5373ad7936dca76797473) +
                      (Ie317e5ea2ca4ba2060d0f491290af96f) +
                      (I56ea52c50a188ec47e48740839a031c9) +
                      (Id9b9a8fe43992ec0793845715dd2226c) +
                      (I93b69bfb228db4b569a6772179d603be) +
                      (I71afab29cdb962e1f1ca21b61dfb50c6) +
                      (I9905e2686b350e8a6e7f790563a91294) +
                      (I524e78ae6a4204e17ba4532dba047d4b) +
                      (({q0_1[5],q0_0[5]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[5],q0_0[5]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00006  <=
                      (I71228fe4188ab1d9796081184a422094) +
                      (Ie19b39200436b0bfca13502ad36c21b9) +
                      (If6657f90c84ca5e2ba08ec705f34be03) +
                      (I60ec7459bbe99fce295406bee1f2af46) +
                      (I29ab844f80c105d247c5c15faa35863c) +
                      (I856fa68463aa5ef1ae53442699d38b33) +
                      (Ic3d00a27f15f8983a120395082854d6b) +
                      (I6b1d01c3cb8fb51e43cdb788b89816be) +
                      (Ib74a56900c1f8b159ad381f61acee801) +
                      (Ia5eba52d169755c507b9e0094e467fab) +
                      (I0899e8fec1a7209cd94757c0b2f87c9a) +
                      (I08ece7cd684e593e02321612b7a88cee) +
                      (I691c84d81c60a462e28e2b2bae3ea845) +
                      (I58dc9cce6384160c0a85c6efb3319cdb) +
                      (I56bf74b5890ec67090f499afdc0a9c88) +
                      (Ibaf2f1f8bda2f6b932dc30f8369c0e1f) +
                      (Id9364a29fd79b52d0442e18dc0227854) +
                      (Ica3a41ace27f7d94377981079952f4f7) +
                      (Ib57795a63d642a73456324bab41384b6) +
                      (Iabf572c97b48c6a7dcc19e56676e3a82) +
                      (Iefd370d0df1a93639af482f78a1e8706) +
                      (I995d2809ffaf0ecda6a004d01cb9c8c4) +
                      (I4e8ebc46bc068c3f9889d970db131112) +
                      (({q0_1[6],q0_0[6]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[6],q0_0[6]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00007  <=
                      (I7b561638da1b4a45ff59be81243e4471) +
                      (If0a3b88a66a816b25f17ced5d0e8f775) +
                      (I0374ada4fe50717f2158468b7ad205d4) +
                      (I357137b41bb91e0659b1ac6ead9b5c12) +
                      (I5d70bc64cf7b3d3ef4180e082e533237) +
                      (I7d9ad929660cd212387d893266b681da) +
                      (I34be4b353cf75603301372840c2f91c2) +
                      (I14834fc8e6489775359bcecf5a37ff4d) +
                      (I633a74e4dfa841c9fd13dbb6564c8493) +
                      (I157bd468200e63385583b9045758d81e) +
                      (I918c46173eebc5b2a95e041cfd91d958) +
                      (I4f8792c18bd07b23e82bbc44b4ca947f) +
                      (I8d0a1ae4c47edf1f2b99d1175aaa7197) +
                      (I734e601f5f9d568a44a48834559e04db) +
                      (Ie421da1dc5aaea57c50d0c7d9c5a2717) +
                      (Ief5cbddfbfb98fce4812a676849b9a98) +
                      (Id113cab2dd1949d32e3c1c15273185c8) +
                      (Icfe1a689e33b2b9aa9dba692d6d610b9) +
                      (Ia4b671f3360f3ce55db0dc0e4d78ddbe) +
                      (I60cbd4369e7ba9b6532f279e5c59084c) +
                      (Ifb6c65a00d9a2c31d8b1119b949828d8) +
                      (I4a777f0dd62b19dd340ad31517c4e789) +
                      (Ib75747cb32130d44b338ed8c8af8ca11) +
                      (({q0_1[7],q0_0[7]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[7],q0_0[7]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00008  <=
                      (Ic7e35cf8d5cd230b94c40714f16e2418) +
                      (Ic51bb9184dfd103703cd0c6ad6edff4b) +
                      (I103f1449c78c47396d6a54dc1c810934) +
                      (I56b3a97dc3037f0bb2eed93a9482c813) +
                      (I51e98035b35a35fdc52f5bab8f19c152) +
                      (Ia6a7f9beaceb08d81012f0e72171252f) +
                      (I21b062856ced09cb9131c01b5e166f32) +
                      (I4f1221ce7880729fe584b42ef3afe6b2) +
                      (Ie7f3f1d6cee7f02ae1b17740ed54c049) +
                      (Ib196f5bcf9152703dc32c5101076600a) +
                      (({q0_1[8],q0_0[8]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[8],q0_0[8]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00009  <=
                      (Ide9ef5a16d8fe32353c2c2a30e8ee3b0) +
                      (Iee6f2484a381bd42e441ff072ec582e4) +
                      (I53121a39de0bcba91a4d0438be2ae958) +
                      (Iff7950f24f0a6b0073942c37fff49d37) +
                      (Ide86f019e9573706c25bd8b4552396a8) +
                      (I2370042234b0e93bb66e44b97fca3e43) +
                      (If9efe7a1c359ec03014a52870ac13aec) +
                      (I6a6eb62960b616043415406ebfc21346) +
                      (I06c7728ef64be8311f48d10d766d0c44) +
                      (I9fe11f6c8147391aa4a5afd1a4e4f731) +
                      (({q0_1[9],q0_0[9]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[9],q0_0[9]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00010  <=
                      (Id50edc56fce48130247fdbc42eeff9ea) +
                      (If3e5161254eb9056914c46263b865c10) +
                      (I58703e8b6d04f8c69ac38f5fcfdc4efc) +
                      (Ie1f41720e296ced1b74cb325b666d88f) +
                      (I5d5701435c96f1078e741921b56e3c65) +
                      (Id96e744d9b10dcddd1ae0115ea57a76a) +
                      (I0c0060fe260afa3cdc72f35ffb6938ff) +
                      (Iaec1f186cb4a65da21d41e637fc628f7) +
                      (I9c15a6a5c0db11ede80ff6d04c9a56d8) +
                      (I8922487573e02d684a3d71448c3828f5) +
                      (({q0_1[10],q0_0[10]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[10],q0_0[10]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00011  <=
                      (I47f17afcd5871fc3ac378316fd3d7ae9) +
                      (Ia9642d79bb50567348083b4435c7d66d) +
                      (I2b2bd845428c49346ef8e94e95b618f8) +
                      (Ib730fdb59198f23d1e590f6d6039e96a) +
                      (I644e83f0a7d432fba38ffb2d99088eca) +
                      (I97f2b15ce0a74e68d5a4438111adcb0a) +
                      (I84c88b631bed5311cb6e99e58941149e) +
                      (I45c5e6710240685bf54b73b0d7a64271) +
                      (I5827bc87b5db1801b7db16e1e61515db) +
                      (I1c85c8f73ef80a6808c6aec0c8eca8ab) +
                      (({q0_1[11],q0_0[11]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[11],q0_0[11]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00012  <=
                      (Id13c99b7f7500c8195b54627efbc4232) +
                      (I4636821315d702a677dc93113872e647) +
                      (I9c981b0614a29386ca5e8ebc06a17f15) +
                      (I4df3d4dac24877b14e6d361bafc1a800) +
                      (I913d818403024510c55b65b56a38dd89) +
                      (({q0_1[12],q0_0[12]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[12],q0_0[12]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00013  <=
                      (I57015930f5b09a6c6b030ed01dad2177) +
                      (Ib54d55a70605119e37e9898b940ff636) +
                      (If7e146da4f3bd255b8457fd6902005f6) +
                      (Ied00d87af99ae55144fdde41ebfc1357) +
                      (I7774313f1ae5a2de98855aad572b3676) +
                      (({q0_1[13],q0_0[13]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[13],q0_0[13]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00014  <=
                      (I679baea452c3c6d04c53baa88edd8eb3) +
                      (If4132b39ddb92aa02d8d0346fb0e6691) +
                      (Iba70e737d52e6812a67c159520e5192f) +
                      (Ib9ceb8315f0cd848f861bab677c2c694) +
                      (I7846bc2cc11e08d05f7c853c4920d555) +
                      (({q0_1[14],q0_0[14]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[14],q0_0[14]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00015  <=
                      (I0865623d3350645e63fa6e6c9b78ac57) +
                      (I0262b30a4efa9f1cfb11d1c3940de9e7) +
                      (I7a2e79d42779ad235bca6ce3757cf588) +
                      (I09e9a3cd4c12d204f760758e873a177b) +
                      (I30b0b1d54912c1a41a02a25ab238bb54) +
                      (({q0_1[15],q0_0[15]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[15],q0_0[15]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00016  <=
                      (I49fb0909ddf66fc0073e6400f1a07844) +
                      (I9938397dc94002481984f5b560fadc58) +
                      (I4378d139db4b710e3587aa72df22b70d) +
                      (Ifa43d74fa91b7b9884969f575ef9ca8e) +
                      (I7c19a79f441ecbb73685db5a505e7479) +
                      (({q0_1[16],q0_0[16]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[16],q0_0[16]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00017  <=
                      (If2af8106efc1f7dd02c074af68278b3d) +
                      (I89a3f8d5f760d1a650f85814cbfdc017) +
                      (Ifae345c79662c3df3dff0fe68ad68746) +
                      (I88a61cf72347d695489909d0819332ab) +
                      (I9aaa036a6158d11c235bdc8406d79f4c) +
                      (({q0_1[17],q0_0[17]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[17],q0_0[17]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00018  <=
                      (Ie8df350430970b5f1229cda772440f85) +
                      (I7d77ac9b64b2e8cae21c6e36947e3ca2) +
                      (Ic1faed76fca5a9ceb7db26c2f43623d9) +
                      (I3ca2b9b77ed8d78a10aff42a07a53b07) +
                      (I1f00849ea055a7893df386aed162a7b6) +
                      (({q0_1[18],q0_0[18]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[18],q0_0[18]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00019  <=
                      (Iaf8a19fde3de660c3fa925593bebbe0c) +
                      (Icd1da43a4d95230e79dbd35a7ae41066) +
                      (Ice9079fb6e08d629f8c0c9ce332c8f11) +
                      (I15fafe2baba4d2f28037023a81ce0a81) +
                      (If4d5b48882e9e628cf51ad2ac2f38c22) +
                      (({q0_1[19],q0_0[19]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[19],q0_0[19]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00020  <=
                      (Id0eef1adba01447c14a6f005782dd9a2) +
                      (I1d1a7c5928982c278d068ebd262254da) +
                      (I6354a0e638340378124e4df7f3d145b8) +
                      (I0236c912c6d684bf4862b725be9d5951) +
                      (I6f3be51d69b2b64a04e55b8946d5dd56) +
                      (Icde3e6dbcf985682041f30903ad95572) +
                      (I46ee30b46020d91707689f3468f00e26) +
                      (I2605f078c1a9006c93855a9a2b0cf6b9) +
                      (I4d226dd2f0bfcdbea6a2e6a6613c1b64) +
                      (I5c942076b173cf527e1be2ddb8560e84) +
                      (Ic95191bccb18e26c10e56be395ca6b1a) +
                      (Ia284f974dd8a526f31eb81ed71a06e94) +
                      (Icc93450a007cee4c0a42717ed7600528) +
                      (I9ec9f389d0489908d497487e44c6edcd) +
                      (({q0_1[20],q0_0[20]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[20],q0_0[20]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00021  <=
                      (If8a527cc7f06a9963a80a880d225d34c) +
                      (I39ff4663007dbc89b403f3b08a69bb6c) +
                      (I9590eb28a81c730b83b92ef7653e71a1) +
                      (I2ba1acca919bddcc22a41a28d43a4e3e) +
                      (I62d8efd4227cb3dc88aa08b6585fafc8) +
                      (I749e987266a20840bb8a4b1a2a2fc5b0) +
                      (I7607af5d98e8070e3d15cee23cdf877e) +
                      (I2e11a697d7f17ac30302eadb500de72d) +
                      (Ia0886ce792e062e22d0c224158cdfb7d) +
                      (I6b3cd79aa87235ff174c0299b855dd3d) +
                      (Ie4ae993ddb776bdffec843db0def2f5c) +
                      (I3ed2da9b53daac0852a06ad1acfad21b) +
                      (Idefa29d4d4e2a6e9147f84893520096f) +
                      (Id1fbbe0594dae272856566522633bb3d) +
                      (({q0_1[21],q0_0[21]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[21],q0_0[21]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00022  <=
                      (I8070a3b7d8b1a7ae90c1a2d27aed09aa) +
                      (Ie88285ce2b9c71de02ebd62e8f44ca72) +
                      (Ica1997c6c569c1d1f45224fbaa4e6b59) +
                      (Iaf08bcaaeb15bb0c971432f7f8b16d0a) +
                      (Idcb37cfc357cc088c775409fb9225b51) +
                      (Ic419255414995e7168afb97b051fa64f) +
                      (Iee6da3120d73373627b25ab7c0dedd28) +
                      (I56fc99a22960232b305d6e683c66fcc7) +
                      (I0a9a09b0ab43d2a0f1d1d01e13f0333c) +
                      (Ibc73d07e0c97a6fcae791e04106cb082) +
                      (I224bbdf94ac86c5c376d1db4f4d4e060) +
                      (I43f2b69c6b427de3095c44d4166b77cd) +
                      (I1e50c90010a3df1a8ce1cff811cc7a0c) +
                      (Ie1817cbf3a80dae435a5571dfbd2f5ad) +
                      (({q0_1[22],q0_0[22]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[22],q0_0[22]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00023  <=
                      (I0052d562fb3182890c8828e52d437b11) +
                      (I1eedecb1d8ff505c75be7787199afada) +
                      (I7ef544597a185b1de63b4ffc4a1d44c2) +
                      (Iadeedf3870f0b1eae98d0f7dbbeff04a) +
                      (I70ae07db9b44d530be220f06401d3d3d) +
                      (I7992ea31927b4f0e268462a3b0f18c5d) +
                      (Iadf927d18644a232ad1f1eba7db82934) +
                      (I2a9c673cdd7ded79e09ada38c0f47e6f) +
                      (Ia86740e870d8063f0266b68ad6d7481d) +
                      (I6627bcdbaa8afb115123777abd45435b) +
                      (I96fe3eb633eff6958ac575b997460bb9) +
                      (Iefdcb71f2903b11f5cb0b8857f7a1727) +
                      (I2eb90278aaa54b9c8212b3b4af7c3617) +
                      (I43493f70f0336453d77caf7f27503daa) +
                      (({q0_1[23],q0_0[23]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[23],q0_0[23]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00024  <=
                      (I26a7fe395eb583258c1ac58aaaa3234a) +
                      (I21668ff77cf75570cae97f575cbcf644) +
                      (Ie48be9e6b6fd63baa104d0a6a4561a1a) +
                      (I05370777439b01811fe7f750d2f724f4) +
                      (Icdcd83341f6b5c404f91ec7e97d0550c) +
                      (Ibba4e82d1510ddc16eb4ef64893cec02) +
                      (Ifb00ae47340bc99669c71da34cccc59e) +
                      (({q0_1[24],q0_0[24]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[24],q0_0[24]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00025  <=
                      (I75a4cf2948bebc58e12bb039ed273ff2) +
                      (I5a9fdec7d7ff99fe33ad6cd8afd9e059) +
                      (I47b1695a74e4d27389b97543415dcc67) +
                      (Ieb38fa62119a5a77c060d6634e051298) +
                      (I3459d98131faef5a5040a03847890b55) +
                      (Ie9b9221b2122087cd5f309570b6d31ca) +
                      (Id4451722e8e2393d627dcd0175dc9903) +
                      (({q0_1[25],q0_0[25]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[25],q0_0[25]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00026  <=
                      (Ic10356f9069e3651b9c045c906e63512) +
                      (Ic3a431f39c678b7175ed30fde1fa6424) +
                      (Ib01cfd833a63500e03333f263805db3d) +
                      (I0b7b4c0a8503c751229edfe0237cc903) +
                      (Iace01234164c8a9f7c98eeb83268745b) +
                      (Iace8b3b3a4c16763132b5aaa6b24212d) +
                      (I80a89644e278e96b1cd1c4b7f764dc34) +
                      (({q0_1[26],q0_0[26]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[26],q0_0[26]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00027  <=
                      (Ia92d2276a8a23521ad1b88df7c27bc2e) +
                      (I39bbec42c442d1e8c818f46ad9c096a8) +
                      (I88f1b5c12759a5efb2d2ded8483c9ed2) +
                      (Iaf4ae293c576af16f5f43a8b86c1aa3d) +
                      (I68b575fcbc5321d4d26a22bcdbb506f6) +
                      (Idf600b93ee1018ecf969ed7944b6bc7b) +
                      (I1cd93172cf5996bc870063aa642188a2) +
                      (({q0_1[27],q0_0[27]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[27],q0_0[27]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00028  <=
                      (I4af080cb4e5cc525db95e5f401019e8c) +
                      (I6fc8044eb226a14ff1a786ddc96d2414) +
                      (I27fd0073dbcdee599fbe85cf48806efc) +
                      (Iaee6d725a8b2653eeac6d5acb91f8f36) +
                      (I4afdeba4fc2a12a6cbe3567a519367fc) +
                      (Ib42816335dd8475dcc78662c4c0786c1) +
                      (I343c9efe71164c01e9c7d599e032864a) +
                      (I108c269ceec4adcff9afeda01101b838) +
                      (I761983331fb6e3c6c437b3f1660f0b6b) +
                      (I70d32affde22f9dcb2d77430fca39069) +
                      (Ic08e85346f61da036a15345a13ac12f0) +
                      (If5dfdadb3868ed5a495007362f7db648) +
                      (Ia1ee5579358b564de06c08ca418a9bf4) +
                      (({q0_1[28],q0_0[28]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[28],q0_0[28]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00029  <=
                      (I9bb81dda8102b829441be46460eb8900) +
                      (I8eef6ca0a61a21882ea28b3d63735228) +
                      (I438522d92cce6f7010246424746ca255) +
                      (I92496f68b44a94565af28a2c28d6fbae) +
                      (I66528f43f614f0edb715564eba3c77c1) +
                      (I8cab9fba615b94fd4bb6934325be8ab8) +
                      (I92d9fec22d36b1baac8bd78abfc1bbd5) +
                      (I4eadce87f47df6d8f0e4acd057de5a09) +
                      (I73203143fe37933c16fff873c1abf512) +
                      (Ibed2a63af723a7abf96dacf1951e5266) +
                      (Id667c80003b5541de9f84d3b8709c828) +
                      (I02cbb4255db2b21ea32140f9e9ddb36b) +
                      (I65354f2069de0c25bbe7cd50fbe892aa) +
                      (({q0_1[29],q0_0[29]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[29],q0_0[29]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00030  <=
                      (Ic279867ebf3055980f3d813d5dc8dec6) +
                      (I5c05da8a222ad5effb9815cbf3ec25f3) +
                      (Ib8bf21f32c0e8b9cfa42a53807bfe3a3) +
                      (I7208256bb198bfce1be71390b01bc028) +
                      (I49f2a06ceb3a59773c65b19f54ff362b) +
                      (I86e495dc894d2aace15c1aff89798bf7) +
                      (I0d53bb5344cabe5fa5ce3ecf7122a260) +
                      (Ib2f5f5fc77ea8b529f2471c54388f2d1) +
                      (Idcada1bfb3c0d1f2a09aab58a2071a57) +
                      (I814b62120953991f9da055f118967e05) +
                      (I123a212546a8ac394051425db4924812) +
                      (Ie95f1a7e0effcec0aa423dc803056a13) +
                      (I106deaff50b8480eac31ddbae2ec7c61) +
                      (({q0_1[30],q0_0[30]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[30],q0_0[30]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00031  <=
                      (I68528be9951f5b8805411711cd11ea59) +
                      (I0f034a8f077b0ab231727b6298e366d8) +
                      (If9c12f8662333fb54a45cfa1bc5da487) +
                      (Ie1681d905517daafcc7584725cd6014c) +
                      (I2ff3edcdb6158f1e3c9a555aeefc0850) +
                      (I43b380be6df7df0d354223d0a0d6d6b6) +
                      (I23eb1dc4d1c992f804dd04a2d823c778) +
                      (I7f90f96c0260560ad5e6dc7448b2670a) +
                      (I07b417cdcc99eaea3413f563e26ddc73) +
                      (I2f3ab9654e515a54e22e73d6c130ccc3) +
                      (Iebdc41368d57498a04fa73e30b10a966) +
                      (I5b4305bef5b4350c1d7ae143667afddd) +
                      (I2795d21d343b83a69146314a2407cfa2) +
                      (({q0_1[31],q0_0[31]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[31],q0_0[31]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00032  <=
                      (Ic6386d7d8813731d612e24b715740275) +
                      (I4c366a57920ff090a98a2cb8b9caa00b) +
                      (I14cf5d43fc9864820a8a25efcc5c6d86) +
                      (I33b99994abbb5ecf8eed4de39033e4f8) +
                      (I7c3291f0250d13ca94802b0b071a95c6) +
                      (I2c926fd9d306e9ae13364e07c4b0395b) +
                      (({q0_1[32],q0_0[32]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[32],q0_0[32]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00033  <=
                      (Ib23edc35fa5bbfe0415fcf0861a22d9b) +
                      (I3e0e682047f7cc36142e668828cbff1e) +
                      (I99fb9030e8361e57818c07511479a9b8) +
                      (Ic87c3d7762a18772972552162e1d1a8c) +
                      (I7e393e6c1d1bc44daaab120d55f5dd59) +
                      (I448f126fd3932d5065abbe7bb2d92c56) +
                      (({q0_1[33],q0_0[33]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[33],q0_0[33]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00034  <=
                      (Ifc8c6df8904b97674f2970ebc95b523c) +
                      (Icd0622a90782b9c451950e7ab0399567) +
                      (I6493b3c087d4685a6b3f98c73dc2ff49) +
                      (I20c2057240417146df144b518b43d052) +
                      (Ied029d0bdea3bf134744c99426fa72dc) +
                      (Icb82c9ff4cb58159a1c3115c6fdd5f8c) +
                      (({q0_1[34],q0_0[34]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[34],q0_0[34]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00035  <=
                      (Ia3450e134e4086c35acbdee1e6042396) +
                      (I5a0f27df5158309f32f0df31e8ae3ae3) +
                      (I17d9e19854cef197fd3267618617efc3) +
                      (I2993acb61f1abe529f8a60c94a438550) +
                      (Ic8be2c94235fb40f78da33179ce4873a) +
                      (Ib3367565e4456da15e7c2315dccdb5e4) +
                      (({q0_1[35],q0_0[35]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[35],q0_0[35]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00036  <=
                      (I15a1671def323cd294591564ae6ef8b1) +
                      (Ic512effb493a06ece58a2af155135004) +
                      (I2c72248cbe49ec0a0febac2437b8a6dc) +
                      (I964e17c41a134c080e9c43412a514f3f) +
                      (I94f1724740defe5bb7e40041d0e266a0) +
                      (Ic19486b6ab0373b9c0ad8f7597782d8f) +
                      (I31243de90dc2a1656ca9d5e03bdd78da) +
                      (I242a30bdc8699d8ff550b25dd53d6c59) +
                      (({q0_1[36],q0_0[36]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[36],q0_0[36]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00037  <=
                      (I9d15f76bb68b214057566cba4b511214) +
                      (I9cc16a00912e7dfc05fb505a9db23cd8) +
                      (Iacf9640cbf486411d6ceb8fe1a2fd5c9) +
                      (I9015033ab0caf3fa41dae4de43f24a82) +
                      (Ia630e59cbce82a570ae3890a6c0221e5) +
                      (I4904ab14b19fa1b6befc218bc7be3842) +
                      (I282d2eb4e74e034694e33273b9cb19d5) +
                      (I3f33901c407a87e10d86c13c83dd52eb) +
                      (({q0_1[37],q0_0[37]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[37],q0_0[37]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00038  <=
                      (I43f41bf07836cee48069e9890c1de2a0) +
                      (Id88480a0a350bb5fcf01ed5fff0bbd4c) +
                      (I1d9b9ff357667a362f0442f19986f451) +
                      (Ice73589836da9028def6efb24a04dbbd) +
                      (Idb72c046c5996fbbd80b706666ffbd92) +
                      (Ie5757e7b1647ab7d43cdbcf98cbb77fc) +
                      (I6072331f838d82329a07a4ffa340c7b6) +
                      (Idf6875955525d80dc660ce956f4a84e7) +
                      (({q0_1[38],q0_0[38]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[38],q0_0[38]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00039  <=
                      (Ia96955d9c0a8a587e0afab37c8415d8c) +
                      (Ifec374bce7f5507438f550df22d61a01) +
                      (Ief67e897e57b96e2ec200e82bbc7caeb) +
                      (Ide604e9bbe35cb55892a4602e18b2527) +
                      (I262f2390e77ec486ccd3a6ed05816e2d) +
                      (I280e20c20c0b4f26278b3de9b2ff84e4) +
                      (Ib3a0307176d424a4733720416d71069d) +
                      (I76060709de3ea188748849f043c59ac0) +
                      (({q0_1[39],q0_0[39]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[39],q0_0[39]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00040  <=
                      (I8be20605d26d218911e80a883a90d085) +
                      (Ieafa9d74d4a61d28ac4a913db460bf33) +
                      (I6fd1b4395af175eff85b3bfeef4c329b) +
                      (I39e6d3fb468aa40ea73535e81556ea65) +
                      (Iae449b74e50e0907feae9e60f2329426) +
                      (Iebf769a6bdaf214c1006c55c608d4eda) +
                      (Ia030c08757123aae947f86ab8bfb6d94) +
                      (I8c35c5b343b552c22000e194c517ca12) +
                      (Ibf80bb564263ea85bd886a8617f09bb2) +
                      (({q0_1[40],q0_0[40]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[40],q0_0[40]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00041  <=
                      (Ib8dfd9b8badef282ca00a4f793c3c868) +
                      (I596ad7e132f272cb196b74faa8c75aa4) +
                      (Idc629414f6d0236ce0714cfaae23f065) +
                      (I157fdf8775206858c08682db3039b084) +
                      (Iacbb4daf5ce5c7eb1a2afe30d0cb5382) +
                      (I4e08021c0235fafb60200aab97827a8f) +
                      (I730634ea15ac94d241f3ad2d6393a227) +
                      (Iee367c535d9c39f872d2ec043e7e7b33) +
                      (I68bb1f26f878862f288c1f57049cf58b) +
                      (({q0_1[41],q0_0[41]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[41],q0_0[41]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00042  <=
                      (Ia9b5d9ede006c56a6d83905529c77b7b) +
                      (I1487170cb1f3370ad45efc801cefc8ab) +
                      (Id88568dd34fbee42c9cb8cc15ac5c31d) +
                      (Ia30539545e66c4cfc16828140149180a) +
                      (Icbfbb37bad6344005dd233b3605a784f) +
                      (I91a6408a11fab36a8ba3dbd3f895a803) +
                      (I47b878f27c30f79a37e97e022307e9e9) +
                      (Ie76b0739aec66f8860870e66e87a6445) +
                      (I50383e3d7c172eedfa00aa50a9faac4c) +
                      (({q0_1[42],q0_0[42]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[42],q0_0[42]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00043  <=
                      (Ifeaa99e03bda8ded058f98387de3d49d) +
                      (I4255ac1af4367c321567c4e46b06ab25) +
                      (Ia445bdc7def7d8c1eec31ab892c25c41) +
                      (Ic3b4752136ac08e343933ccc3a4ec47c) +
                      (Ica6707efd6d44ba6bbb87c0593a3d828) +
                      (I739267bcc50c54b8a685cb3c6afc5cc1) +
                      (I9160d11439c5140c0109b5190eb82e6b) +
                      (I6ff7b86cd7f63f9243646f1be10b2577) +
                      (I165653ab165cfafe2b74cd441331f9e1) +
                      (({q0_1[43],q0_0[43]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[43],q0_0[43]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00044  <=
                      (I08a8cd6965c23af6650568b654831b20) +
                      (I9b6a674dbcbfcf65f1ae0deb8fc3566d) +
                      (Ie3a336de822ac7baf8486b1618ef1126) +
                      (I5fc3c26d6c5aa893dfd5caa0f677233a) +
                      (Ie22b94121b58f17af14c75bfb27f96dd) +
                      (I0d9f8c99194d9d6e187b4ad02fcce8b4) +
                      (I71e101962e766a4d1484b3235359a4b5) +
                      (If2539da6722562bbf31786fd0036666a) +
                      (I22c8ccd4a9018ad1c129aa058bf579d8) +
                      (I83330fef69470d2f5def8e6d7d9c50d2) +
                      (I0539d598bbe3d50940329a282c801328) +
                      (I202f88fdc946494d55fc8831c2e8a34c) +
                      (I3ee10f6a7785a236db317515fdd23a2d) +
                      (I453fdf4fbb5af5bd28a20d7643da9eb2) +
                      (Ic4a6c02880a9aead7353332708e3f388) +
                      (I7fb3b66cb48521f8715f66bf5642cdb2) +
                      (({q0_1[44],q0_0[44]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[44],q0_0[44]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00045  <=
                      (I2fd872df07f50688486c0d602cfc5549) +
                      (Iccefa45795486757515d95e5908b306a) +
                      (Ib1357cb20f471f1670ac2448f964f8eb) +
                      (Iab953a8974a1eb619dc0f074c003b5f9) +
                      (I6e37582849c2c98fd15ad92d22c222da) +
                      (If004de0cac6e5f7701a1fce48c6936d5) +
                      (Ic1efa395cc1fd2c5a1d1559fb169a5a0) +
                      (I8e96c69e7d872be23229353808c34953) +
                      (Ib6aded6c73a8cc3cb964b0ae895b859e) +
                      (I939368b76d98b43826c68c7f468a5632) +
                      (I544f6263f16cd5e0b7cf28c511a8f6e3) +
                      (I484545c4d2c869d79eb17f51e11070a3) +
                      (I39289e6385a9bc378a9b8dd440249a7f) +
                      (Ie9cce5746a83479a567bbaeac6dbf497) +
                      (Ic044d7419cc43736d278c2df33b4a3cc) +
                      (I6714551e8885ef5e4490673fe1b2dad1) +
                      (({q0_1[45],q0_0[45]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[45],q0_0[45]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00046  <=
                      (Ie9ab3c88ac62369e3d92d110165a94a8) +
                      (If38feb4f76f761dce6145731ad235d7f) +
                      (I6359856a1843d8c8b65dc478bccb3acd) +
                      (If6f3d91c3c7a43622b9a522492cd83d3) +
                      (Id023a6298e65da1f4da3831f5136afc2) +
                      (I6b24690f394792edb0d82b3b9e110851) +
                      (I5b55c285f7e3e78447fee68532ab9f7f) +
                      (I32701d9e4b96853c53f0ab651a6a4ba2) +
                      (I82f266e5792cdb6e7ebd264e246161f5) +
                      (Ibfacfe5b83819afe7fbd4bffa2d6d4e2) +
                      (Ib8e68a77ad8b9e7cf415bee17645c3f9) +
                      (I644ee0055a55f54ab3544bb532e39c61) +
                      (Ic5467e42aa377c6ffd8f70673808774f) +
                      (Ic57eb4a034247a4c952d8224ea9f2bac) +
                      (Ia642db613c0ec1ca4e69afde7a14a839) +
                      (I432aa7cb844286c442356954f8814260) +
                      (({q0_1[46],q0_0[46]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[46],q0_0[46]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00047  <=
                      (If520c1cd27f9d4bc52d0d029f693b660) +
                      (Ie87075ac979410cc11099a356966b8a2) +
                      (I6fab46b1766878b26b53f352fee98223) +
                      (Ieaf14683f40374c4531326d228cb43c3) +
                      (I5149125aaaad943d891df6a3c2be93a0) +
                      (I770dff588ee1f52f58bea1921cb23383) +
                      (I8f0a90e761111a613d2488285534a500) +
                      (I765a8825e42180a6c63f7b33703bb483) +
                      (I512cc8f6519aa08aee18225b56d47c9f) +
                      (If08370fd0e8af818c6db20f43e74034d) +
                      (I0ff382edfc8051459657ffa3899f5f73) +
                      (I9d2864024148337277523ef7fa2e1600) +
                      (I1c85a2d1df6749a194072eb731506bfe) +
                      (I3e3ce8b4ead150a6eae2e5c701c7b598) +
                      (I45bc13ae0e0554a79c62cd9c6aa8f2a5) +
                      (I92678f5b52c9c55556ff7f17f0f607b7) +
                      (({q0_1[47],q0_0[47]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[47],q0_0[47]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00048  <=
                      (Ib4bdc9069d0c08655f5e87f705943eda) +
                      (Idbf9094c94c931f16fba468b9dd59a25) +
                      (I1c3c4ce44610e04c5eef2fcbc2ea5114) +
                      (Ie84be0ae8311d906eff08f7f5b214943) +
                      (Ic90b98708faa8c8b75d4bd9a52c292f7) +
                      (I8eba6f14f42701d22859fbea94bd1871) +
                      (I6d83efa9f988328f487e9232bf2633a2) +
                      (Ic23e01562c8a753fd70c343297be288a) +
                      (I5669856f88f5e2c98f64df696db76414) +
                      (({q0_1[48],q0_0[48]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[48],q0_0[48]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00049  <=
                      (Ic3a608b850709286ea0ad2f67425d9ac) +
                      (I5267fa34449e6eebe891017fc32d0749) +
                      (I599d01cfe6e54d8e45d64446c446818d) +
                      (I8f94dbafaac589ac9f14b56d4556ff96) +
                      (I754563caea429d3d0e22df5d193b84eb) +
                      (If7f373506cac70f8ba1222db135c27e8) +
                      (I69f563e7b7ad483893ac9c4684349769) +
                      (Ia0a02781c674fe5d769206448d475245) +
                      (I1b7a401bc11741e6f011fb9895b5c797) +
                      (({q0_1[49],q0_0[49]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[49],q0_0[49]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00050  <=
                      (Ieb528d666fdb708279184bb59eac25d9) +
                      (Ic3ff7ce12c836bf0693252b9a7a7cfe8) +
                      (I19bba6a58ad3ef959b33701f82761984) +
                      (I8acc93b34974c1e708b0e1591f7b2d3d) +
                      (Ib60d4ac0fcadcdfce5a14fb92f58423f) +
                      (I039f05d5be891a37e04556f1eae674d2) +
                      (Id0f75e19b94541ed5c5c352d13390d2d) +
                      (Ife1190f76c2e251704c2960c23330a48) +
                      (Id3e0c98bff2636e216b4d3a0ffd51054) +
                      (({q0_1[50],q0_0[50]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[50],q0_0[50]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00051  <=
                      (If4d3b31b87c0f723241d35ce7e854eba) +
                      (I72369dedfe36cb22269033cc305b730c) +
                      (Iec71fe7fcebccf1ae0d10a5d187fcc44) +
                      (Ie11da10808c4ca84f399535df6261307) +
                      (I280fa9d114e227cd649bf0e55e845651) +
                      (I94c4e11670b4233fa072517a8f19c901) +
                      (I4dca2dd40a7127ce44f83b430a34c738) +
                      (I1a24e98165afa62bd14986911a36fb6e) +
                      (Ife1164cad7cda4aa9a08d94dfe86add6) +
                      (({q0_1[51],q0_0[51]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[51],q0_0[51]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00052  <=
                      (I8d8d95ff26f33f69a182b32ccde23905) +
                      (I2508854bcbab37bd09c9465c377c06aa) +
                      (I140078292f7209eccacd53a8bab18016) +
                      (I141fb1cbe09f9abe282cffd4de815d25) +
                      (If79d1d378f7c6fd29fc3335ec5f5c51d) +
                      (I4a41999cea9357a85c73a0af509eeac9) +
                      (I8e517c401d62dbb10dcc96ab536f6afb) +
                      (I8ad3627f171eadcc960a688ac0afcbc0) +
                      (I85c4d3d6c8408c6f38741257ed177ca6) +
                      (Id66c47fd69c175a4393e975a269cf053) +
                      (I37dca40506d61bdeab1255ed4892ca20) +
                      (I340c98b886123c541a1b8d9fc8a6d48c) +
                      (({q0_1[52],q0_0[52]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[52],q0_0[52]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00053  <=
                      (I2dc64c3b06588542b027f997437bee63) +
                      (Id92a37c091100e9df08e24498ecb4022) +
                      (I74a4b9365391fd20c34588002ad40547) +
                      (I461195b7ae78743e09ee50486ad6ebe5) +
                      (I356d747600182675699a2d2634d4c5ce) +
                      (I87d6a5d30c3e4202cf51f33c7a770c51) +
                      (I960768a84aec9d5b8bc7c1c523024a25) +
                      (I09b5273bb15d48a7fd78559930fa6d1c) +
                      (I5814a85c45fd0f7be21ed325235fe4b7) +
                      (Ib06b60cf9933dd8952206c5f3ccced8e) +
                      (I67347c413b5efd8ff9e0d5bc7ab2a047) +
                      (I72b1bb104bf2843f161448baf7aab44b) +
                      (({q0_1[53],q0_0[53]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[53],q0_0[53]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00054  <=
                      (Ib23d889edb5a6d9f27de977d3b1a2616) +
                      (Ifaff9dd032cf96487be819c59b03000a) +
                      (I028ce03be0618b816e0ecdf43d4cd6e6) +
                      (I6ae2523095237282533e0b5f1c26b488) +
                      (I5aba6218461e8d571be03a3ef041ebaa) +
                      (I6ca8a1fa2c72b1c61d11dc7d1ba5f37b) +
                      (I3ec5819176ad4b0895a9118d90ab22b5) +
                      (I49b64469d298012dbb131d879bff38d6) +
                      (I95361d5f524ccb9feb42811af5c482e2) +
                      (I9c4b34b5fb1d59c132bcaeb6258675df) +
                      (I613d4b1e3b9e812b785c9cf14fefdfe6) +
                      (I848ed394bd4f0b199d11c0ff458394a7) +
                      (({q0_1[54],q0_0[54]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[54],q0_0[54]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00055  <=
                      (Ie65a0634454381e24bb3223a333e3ad0) +
                      (Iad166146f7df5e8068fc6efe4d3e4141) +
                      (I63e45abd4d27219bddcef06108b72021) +
                      (Id1bacd13718f7c29c26b63c239d04dd8) +
                      (Ia3104c69fb4f7abfb5efa3874169a7ad) +
                      (Ie1b7257c99831ec5864f65958ecf14fb) +
                      (I4accbad1b451ed2b622e15ef9ae16d13) +
                      (I5ce8b2f633011e89356243a1a71edeb6) +
                      (I3e5139f24e3d082eb31b0e61ea9fa1aa) +
                      (I61cc8a0f49e393721a62a776e4793deb) +
                      (Ie631e40caade823a196370fc3358f042) +
                      (I4c971e714427664c59c6371e14781bae) +
                      (({q0_1[55],q0_0[55]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[55],q0_0[55]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00056  <=
                      (I36ca732e811d67cd742d24fd4cae887b) +
                      (({q0_1[56],q0_0[56]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[56],q0_0[56]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00057  <=
                      (I354fdd241d5d07f0d8380fe8924e0a8c) +
                      (({q0_1[57],q0_0[57]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[57],q0_0[57]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00058  <=
                      (Id38b705f5d2863a020a475ffffc8afd6) +
                      (({q0_1[58],q0_0[58]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[58],q0_0[58]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00059  <=
                      (Id6e5d67e7bb7c4b999459374ea80459a) +
                      (({q0_1[59],q0_0[59]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[59],q0_0[59]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00060  <=
                      (I05341013abd4206eb66fcddfd63bfe26) +
                      (({q0_1[60],q0_0[60]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[60],q0_0[60]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00061  <=
                      (I15da71a21f5842cb65b543d9bc3e267b) +
                      (({q0_1[61],q0_0[61]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[61],q0_0[61]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00062  <=
                      (Iccf255fb3422c558465e45226068a16d) +
                      (({q0_1[62],q0_0[62]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[62],q0_0[62]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00063  <=
                      (I1c2674b2e6b269ed539827412c5199a5) +
                      (({q0_1[63],q0_0[63]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[63],q0_0[63]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00064  <=
                      (I6a3f405bb4a0c4448d9b9d3dd95d036c) +
                      (({q0_1[64],q0_0[64]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[64],q0_0[64]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00065  <=
                      (Ib528bb7a64cce4f694081d151fa6fa86) +
                      (({q0_1[65],q0_0[65]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[65],q0_0[65]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00066  <=
                      (Iaa40bd3abf668a21e0f87c7bda7b3f69) +
                      (({q0_1[66],q0_0[66]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[66],q0_0[66]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00067  <=
                      (I919d36a7f6ad42c4bbc23222beb73106) +
                      (({q0_1[67],q0_0[67]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[67],q0_0[67]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00068  <=
                      (I648d2a279dd1f587b1e45eeb35f2fa90) +
                      (({q0_1[68],q0_0[68]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[68],q0_0[68]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00069  <=
                      (I194a64bef92ecf6714141eaa5d41c9d4) +
                      (({q0_1[69],q0_0[69]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[69],q0_0[69]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00070  <=
                      (Id332e7f482524adeac7f7cdafcf5ca46) +
                      (({q0_1[70],q0_0[70]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[70],q0_0[70]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00071  <=
                      (I226383d68f89db716cfd8d08b837865a) +
                      (({q0_1[71],q0_0[71]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[71],q0_0[71]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00072  <=
                      (I2bdf5d319ba9089a4da34b108f5c5ae5) +
                      (({q0_1[72],q0_0[72]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[72],q0_0[72]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00073  <=
                      (Ia91800792941ec7cc60415c3f844e4ed) +
                      (({q0_1[73],q0_0[73]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[73],q0_0[73]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00074  <=
                      (Id7c507d96098ee7a955af8a48ee5d72a) +
                      (({q0_1[74],q0_0[74]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[74],q0_0[74]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00075  <=
                      (Ie15e4c1bcdb0e18085d4b320ac6a925c) +
                      (({q0_1[75],q0_0[75]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[75],q0_0[75]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00076  <=
                      (I5485d9edcafc6202f6e5f0969979802f) +
                      (({q0_1[76],q0_0[76]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[76],q0_0[76]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00077  <=
                      (I7fe364f9f537cbef782e7007848a1c10) +
                      (({q0_1[77],q0_0[77]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[77],q0_0[77]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00078  <=
                      (I52dcf5bace9cadcf8a895aaa6a8c1da8) +
                      (({q0_1[78],q0_0[78]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[78],q0_0[78]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00079  <=
                      (I13a9eec6175e695ab8bc4516cf57d6ec) +
                      (({q0_1[79],q0_0[79]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[79],q0_0[79]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00080  <=
                      (Iee73a7c685a4cee03f33d3ef379b1c8a) +
                      (({q0_1[80],q0_0[80]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[80],q0_0[80]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00081  <=
                      (I740dc91716e3906ad078e2c7cc3c925a) +
                      (({q0_1[81],q0_0[81]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[81],q0_0[81]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00082  <=
                      (I514d2dc697e9b39ba027c418a6df6cb9) +
                      (({q0_1[82],q0_0[82]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[82],q0_0[82]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00083  <=
                      (I782726e317a2aada9e755bcbc4b0d3fa) +
                      (({q0_1[83],q0_0[83]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[83],q0_0[83]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00084  <=
                      (I11eb26cf0f0b3a334e8f7317bf8d9eb0) +
                      (({q0_1[84],q0_0[84]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[84],q0_0[84]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00085  <=
                      (I26cb63ba20245b2c332b09e25c4409aa) +
                      (({q0_1[85],q0_0[85]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[85],q0_0[85]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00086  <=
                      (Idd7691d31f8d0c09ee988116d574ec59) +
                      (({q0_1[86],q0_0[86]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[86],q0_0[86]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00087  <=
                      (Iecc02842a2d2b9b9e8187f2d39e62e05) +
                      (({q0_1[87],q0_0[87]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[87],q0_0[87]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00088  <=
                      (I5551342f1751fc64f32744a46b9649be) +
                      (({q0_1[88],q0_0[88]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[88],q0_0[88]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00089  <=
                      (Iff7c29299f005c1cd5a16b64601e727e) +
                      (({q0_1[89],q0_0[89]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[89],q0_0[89]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00090  <=
                      (I17a5446e942bcc1dc2c96930e0a87a70) +
                      (({q0_1[90],q0_0[90]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[90],q0_0[90]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00091  <=
                      (I719b67f84e07e90dfd29a8cd5d94cf39) +
                      (({q0_1[91],q0_0[91]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[91],q0_0[91]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00092  <=
                      (I2c835dfb3596b8bf057a7cc21122c81f) +
                      (({q0_1[92],q0_0[92]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[92],q0_0[92]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00093  <=
                      (Ib71b3d357c98dcdfae5c777ca3082275) +
                      (({q0_1[93],q0_0[93]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[93],q0_0[93]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00094  <=
                      (I086bf19f620c8a8f6888e775cb1ed7f4) +
                      (({q0_1[94],q0_0[94]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[94],q0_0[94]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00095  <=
                      (I802c554d5b04af6b949677819a4966ed) +
                      (({q0_1[95],q0_0[95]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[95],q0_0[95]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00096  <=
                      (Iceefb06cb3715e1b41e6f7d89420e5ba) +
                      (({q0_1[96],q0_0[96]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[96],q0_0[96]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00097  <=
                      (I56948bc48c0220893d68004615a6ebaa) +
                      (({q0_1[97],q0_0[97]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[97],q0_0[97]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00098  <=
                      (Iec1368f034655d61354ab5b5e94d7d89) +
                      (({q0_1[98],q0_0[98]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[98],q0_0[98]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00099  <=
                      (I1e43c0aeeb8a2461d208eba24967af30) +
                      (({q0_1[99],q0_0[99]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[99],q0_0[99]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00100  <=
                      (Ia6eb85b127cf9c1a437611556296b967) +
                      (({q0_1[100],q0_0[100]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[100],q0_0[100]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00101  <=
                      (Ieba89aa901e61218074af53a2484a74b) +
                      (({q0_1[101],q0_0[101]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[101],q0_0[101]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00102  <=
                      (I8b3b875c6c07bd97ba598a5139156fa4) +
                      (({q0_1[102],q0_0[102]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[102],q0_0[102]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00103  <=
                      (I7b33ddad346077928620344542b9481e) +
                      (({q0_1[103],q0_0[103]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[103],q0_0[103]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00104  <=
                      (I11d967a5c5d14c88b5587d4cfed1d05f) +
                      (({q0_1[104],q0_0[104]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[104],q0_0[104]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00105  <=
                      (I27458d76b3ac6520fb379405c6b2956f) +
                      (({q0_1[105],q0_0[105]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[105],q0_0[105]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00106  <=
                      (I2525111a2fb5f10d64bbd16e148653b8) +
                      (({q0_1[106],q0_0[106]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[106],q0_0[106]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00107  <=
                      (I7b7cbcd1c6d2a2eeaaff474536a69eed) +
                      (({q0_1[107],q0_0[107]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[107],q0_0[107]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00108  <=
                      (Id2a7f0781d18dccc7c4e0b383b7cddfa) +
                      (({q0_1[108],q0_0[108]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[108],q0_0[108]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00109  <=
                      (If8bc141d98ebe1be7fa81cde5c65868e) +
                      (({q0_1[109],q0_0[109]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[109],q0_0[109]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00110  <=
                      (I8645e1326c66f5efef4b9c923599d1a3) +
                      (({q0_1[110],q0_0[110]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[110],q0_0[110]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00111  <=
                      (I0426ef66185128dd1ef4dbb68dcda585) +
                      (({q0_1[111],q0_0[111]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[111],q0_0[111]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00112  <=
                      (Iddd954df5bae9b4240e0512f746669a9) +
                      (({q0_1[112],q0_0[112]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[112],q0_0[112]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00113  <=
                      (I29e940970d87e8e09b26ab1b0b8f2286) +
                      (({q0_1[113],q0_0[113]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[113],q0_0[113]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00114  <=
                      (I488f6d9676aa85a55d030bf12e8997a7) +
                      (({q0_1[114],q0_0[114]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[114],q0_0[114]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00115  <=
                      (I99d761b75ade1fb2e8afbb1a77752609) +
                      (({q0_1[115],q0_0[115]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[115],q0_0[115]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00116  <=
                      (Iac4e3d20178049f9c59abf374752dccc) +
                      (({q0_1[116],q0_0[116]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[116],q0_0[116]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00117  <=
                      (I618d33f26badabfa578908903a613bce) +
                      (({q0_1[117],q0_0[117]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[117],q0_0[117]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00118  <=
                      (I822d7973afe090b2764335f1b72dfd0e) +
                      (({q0_1[118],q0_0[118]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[118],q0_0[118]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00119  <=
                      (I12c1035353e553b3b6a13bb174ce6020) +
                      (({q0_1[119],q0_0[119]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[119],q0_0[119]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00120  <=
                      (Ia6d61947d36fc128c689808c82db80f6) +
                      (({q0_1[120],q0_0[120]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[120],q0_0[120]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00121  <=
                      (Ie9b042f686381739b9ff219041f1e0ce) +
                      (({q0_1[121],q0_0[121]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[121],q0_0[121]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00122  <=
                      (I0c4268c01aed70ce4fc71531bf4bb862) +
                      (({q0_1[122],q0_0[122]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[122],q0_0[122]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00123  <=
                      (Ia34e42f8de91fa4861b0c6cac5dcfc29) +
                      (({q0_1[123],q0_0[123]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[123],q0_0[123]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00124  <=
                      (Ib7c5850b4f7cc77be2048d114a2128d9) +
                      (({q0_1[124],q0_0[124]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[124],q0_0[124]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00125  <=
                      (I32bb50faa2b246b2d3b462a79be597c5) +
                      (({q0_1[125],q0_0[125]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[125],q0_0[125]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00126  <=
                      (Idc6d40a49f05c5422758cee50f787eb1) +
                      (({q0_1[126],q0_0[126]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[126],q0_0[126]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00127  <=
                      (Ide1d7dc22a4b271ef764df14ac22366a) +
                      (({q0_1[127],q0_0[127]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[127],q0_0[127]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00128  <=
                      (I7ace6778ac86b3e05939a3fcc716136f) +
                      (({q0_1[128],q0_0[128]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[128],q0_0[128]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00129  <=
                      (I044e01e8d2df46e03f00a0af2beb0bf5) +
                      (({q0_1[129],q0_0[129]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[129],q0_0[129]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00130  <=
                      (I45a7ddcda2662e36b7617dfe64514346) +
                      (({q0_1[130],q0_0[130]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[130],q0_0[130]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00131  <=
                      (Idada779a1ac7b844867571d77054b657) +
                      (({q0_1[131],q0_0[131]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[131],q0_0[131]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00132  <=
                      (Ieeba01b18a244ab8c0ac263c138fabcc) +
                      (({q0_1[132],q0_0[132]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[132],q0_0[132]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00133  <=
                      (Ie4c9797a955778694dd8615219cb51e7) +
                      (({q0_1[133],q0_0[133]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[133],q0_0[133]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00134  <=
                      (I28a5ed4c239e64c76bb6e566b50cfd23) +
                      (({q0_1[134],q0_0[134]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[134],q0_0[134]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00135  <=
                      (I79a705ee1e414fe4a5fb14e9b3ce9597) +
                      (({q0_1[135],q0_0[135]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[135],q0_0[135]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00136  <=
                      (I04f90a907f10a7fa1ae3591b48094d5c) +
                      (({q0_1[136],q0_0[136]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[136],q0_0[136]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00137  <=
                      (I31d25b1b49e65216e90b39aa27acd6be) +
                      (({q0_1[137],q0_0[137]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[137],q0_0[137]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00138  <=
                      (I1f6540c5f037d861dee2c0091cba01ec) +
                      (({q0_1[138],q0_0[138]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[138],q0_0[138]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00139  <=
                      (I9632bb500b7faaaaeb649d74c21cbe8c) +
                      (({q0_1[139],q0_0[139]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[139],q0_0[139]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00140  <=
                      (Idd0217a35c3adc8abc7bb581a5df7a2d) +
                      (({q0_1[140],q0_0[140]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[140],q0_0[140]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00141  <=
                      (Ic05b46168884322644db4e331d37d759) +
                      (({q0_1[141],q0_0[141]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[141],q0_0[141]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00142  <=
                      (I53c88dc237bb2cd02d50fd7f0a168a48) +
                      (({q0_1[142],q0_0[142]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[142],q0_0[142]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00143  <=
                      (I7450d4ab3ef0227e93a02bfd620d047b) +
                      (({q0_1[143],q0_0[143]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[143],q0_0[143]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00144  <=
                      (I2b16e5b4e279bb29c3c675b72083e5fe) +
                      (({q0_1[144],q0_0[144]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[144],q0_0[144]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00145  <=
                      (I70c92e8ada46476d15ef4b3c620d2601) +
                      (({q0_1[145],q0_0[145]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[145],q0_0[145]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00146  <=
                      (Ib193b07804d6d5f111b06bda487bfa5f) +
                      (({q0_1[146],q0_0[146]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[146],q0_0[146]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00147  <=
                      (I885433b0ab16c6d87abe45af13c9e529) +
                      (({q0_1[147],q0_0[147]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[147],q0_0[147]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00148  <=
                      (I198c055930cb89d0390c336eda8fed4f) +
                      (({q0_1[148],q0_0[148]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[148],q0_0[148]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00149  <=
                      (I688a2c72e69b217d2673e8da75146a83) +
                      (({q0_1[149],q0_0[149]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[149],q0_0[149]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00150  <=
                      (I3b6fde4ed14cd68af1468ae1d4cc1a22) +
                      (({q0_1[150],q0_0[150]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[150],q0_0[150]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00151  <=
                      (I5d3df1e7563630311f56143ee6d97a8e) +
                      (({q0_1[151],q0_0[151]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[151],q0_0[151]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00152  <=
                      (I90a7ea789d3bf7f9126c786474a56da0) +
                      (({q0_1[152],q0_0[152]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[152],q0_0[152]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00153  <=
                      (I5029424c9d9fe923eeb858b1e62cd758) +
                      (({q0_1[153],q0_0[153]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[153],q0_0[153]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00154  <=
                      (I1e805c70d50c2765b4a03ad2982dc421) +
                      (({q0_1[154],q0_0[154]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[154],q0_0[154]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00155  <=
                      (Iba58175a7fd5c5da650222193caff0b3) +
                      (({q0_1[155],q0_0[155]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[155],q0_0[155]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00156  <=
                      (I7401a0501ba69c5559fbf00c77e58dc5) +
                      (({q0_1[156],q0_0[156]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[156],q0_0[156]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00157  <=
                      (Idd9f7ea657ea9cdcb45a7e4b573b9d50) +
                      (({q0_1[157],q0_0[157]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[157],q0_0[157]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00158  <=
                      (I53f275395dd6be17961a5edc3e8da7f2) +
                      (({q0_1[158],q0_0[158]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[158],q0_0[158]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00159  <=
                      (Icab010d78cd66b02e089c74f04bf4e75) +
                      (({q0_1[159],q0_0[159]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[159],q0_0[159]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00160  <=
                      (I376a48b7e0195a5aacc76a0ad8bd14b2) +
                      (({q0_1[160],q0_0[160]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[160],q0_0[160]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00161  <=
                      (I241622b0367dde514f96ece55c8c3964) +
                      (({q0_1[161],q0_0[161]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[161],q0_0[161]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00162  <=
                      (If94a1abfb972f63629d07e64dc23863c) +
                      (({q0_1[162],q0_0[162]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[162],q0_0[162]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00163  <=
                      (I07b9b1f4fa01b16cc69356057d3b6154) +
                      (({q0_1[163],q0_0[163]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[163],q0_0[163]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00164  <=
                      (I2288a6ad3b748b716249f4adc42d52c4) +
                      (({q0_1[164],q0_0[164]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[164],q0_0[164]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00165  <=
                      (I022df337bcc05ac5648b8ae2e42f3a76) +
                      (({q0_1[165],q0_0[165]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[165],q0_0[165]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00166  <=
                      (I60d9a7f95fb8623753002ecaf9a4efcc) +
                      (({q0_1[166],q0_0[166]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[166],q0_0[166]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00167  <=
                      (I23a74ea5e7174d95e6d16a5e85ac236b) +
                      (({q0_1[167],q0_0[167]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[167],q0_0[167]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00168  <=
                      (Ie697d28d757df82b3901564bda43251c) +
                      (({q0_1[168],q0_0[168]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[168],q0_0[168]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00169  <=
                      (I8572aedc94f7243ce5eacb332c81eae2) +
                      (({q0_1[169],q0_0[169]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[169],q0_0[169]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00170  <=
                      (I6734123aaf6320da75638b212812732f) +
                      (({q0_1[170],q0_0[170]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[170],q0_0[170]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00171  <=
                      (I7f6dc6f0f403c58f9aaaa70c2383a666) +
                      (({q0_1[171],q0_0[171]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[171],q0_0[171]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00172  <=
                      (I66391978843c39b6acbdb4847a01050a) +
                      (({q0_1[172],q0_0[172]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[172],q0_0[172]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00173  <=
                      (I4f756e4125c8af5c412944b273e01cb0) +
                      (({q0_1[173],q0_0[173]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[173],q0_0[173]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00174  <=
                      (Id2c9f7ac95de07148c54803f69347f56) +
                      (({q0_1[174],q0_0[174]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[174],q0_0[174]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00175  <=
                      (I5061e13a179d27e1ba5f89ce8ee0fd4a) +
                      (({q0_1[175],q0_0[175]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[175],q0_0[175]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00176  <=
                      (I0f7c32fc1548fb49b8041f55c157498a) +
                      (({q0_1[176],q0_0[176]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[176],q0_0[176]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00177  <=
                      (I89ffab735ee30423c82e079ed98216c5) +
                      (({q0_1[177],q0_0[177]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[177],q0_0[177]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00178  <=
                      (I9494921d8487ee0b314f75cf0380fd2f) +
                      (({q0_1[178],q0_0[178]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[178],q0_0[178]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00179  <=
                      (If2b3e7d1541cbd8ffc2b4cfc3ad13a57) +
                      (({q0_1[179],q0_0[179]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[179],q0_0[179]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00180  <=
                      (Idf3d79da44f2d686f5bd43c3c1427430) +
                      (({q0_1[180],q0_0[180]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[180],q0_0[180]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00181  <=
                      (If8125ad3c9e7f0a2b84106064d320996) +
                      (({q0_1[181],q0_0[181]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[181],q0_0[181]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00182  <=
                      (Ic9018b88fa91fb638bbab0613795ae13) +
                      (({q0_1[182],q0_0[182]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[182],q0_0[182]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00183  <=
                      (Iad4ea0196eb32f9a152c9e6fe5059e46) +
                      (({q0_1[183],q0_0[183]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[183],q0_0[183]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00184  <=
                      (Ia8ff29ed728e7f2ae4213f00328b495d) +
                      (({q0_1[184],q0_0[184]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[184],q0_0[184]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00185  <=
                      (I70717726200ec02929f679ef05496455) +
                      (({q0_1[185],q0_0[185]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[185],q0_0[185]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00186  <=
                      (Iaf1e4c7dae6ad89567836877c08f57d2) +
                      (({q0_1[186],q0_0[186]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[186],q0_0[186]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00187  <=
                      (Icd09aa81e9b43528af73e23b2f0f80cb) +
                      (({q0_1[187],q0_0[187]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[187],q0_0[187]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00188  <=
                      (I6ebb2b94f0f80425f8401ae823d92a1d) +
                      (({q0_1[188],q0_0[188]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[188],q0_0[188]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00189  <=
                      (I4a2c3204a6a9936d4a215b46c0ffd045) +
                      (({q0_1[189],q0_0[189]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[189],q0_0[189]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00190  <=
                      (Ib02c0694762c4815448b2c8d3df767c2) +
                      (({q0_1[190],q0_0[190]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[190],q0_0[190]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00191  <=
                      (I98cee6efbbe565d3a4de16703189782f) +
                      (({q0_1[191],q0_0[191]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[191],q0_0[191]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00192  <=
                      (Ibf981c01a9d44cbea3c6d8ead92bc2ab) +
                      (({q0_1[192],q0_0[192]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[192],q0_0[192]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00193  <=
                      (I864c33e8ea204d20a9baef4584f22d4e) +
                      (({q0_1[193],q0_0[193]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[193],q0_0[193]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00194  <=
                      (I6ad3228e0e2e1f19648d73e83ba5a229) +
                      (({q0_1[194],q0_0[194]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[194],q0_0[194]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00195  <=
                      (Ie099210a99a4899c53baf39559592690) +
                      (({q0_1[195],q0_0[195]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[195],q0_0[195]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00196  <=
                      (Ieeec71d9df4613555fade2ced7b3baf1) +
                      (({q0_1[196],q0_0[196]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[196],q0_0[196]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00197  <=
                      (I4931884e3544af182bcda9061091a42d) +
                      (({q0_1[197],q0_0[197]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[197],q0_0[197]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00198  <=
                      (Ib3fb10da528d450251764a9b9ede0dba) +
                      (({q0_1[198],q0_0[198]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[198],q0_0[198]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00199  <=
                      (Icdc9e676957b2223d60c413331fa982f) +
                      (({q0_1[199],q0_0[199]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[199],q0_0[199]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00200  <=
                      (I381f6051282c062ccf53866830344cd4) +
                      (({q0_1[200],q0_0[200]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[200],q0_0[200]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00201  <=
                      (Icfc21935c007fbbceb2a67ebe1a68a0b) +
                      (({q0_1[201],q0_0[201]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[201],q0_0[201]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00202  <=
                      (I120d597a80158374726e064fb0f099fb) +
                      (({q0_1[202],q0_0[202]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[202],q0_0[202]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00203  <=
                      (I2520aa556aadf851f58f0b1820498730) +
                      (({q0_1[203],q0_0[203]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[203],q0_0[203]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00204  <=
                      (I6203f49a08107f7185ebadeecf2c16b0) +
                      (({q0_1[204],q0_0[204]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[204],q0_0[204]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00205  <=
                      (Ia706fb593b63cebbee0321c154cb859b) +
                      (({q0_1[205],q0_0[205]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[205],q0_0[205]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00206  <=
                      (Ia4b5f2b07556629673fc6576bc49a5dc) +
                      (({q0_1[206],q0_0[206]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[206],q0_0[206]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               sum0_00207  <=
                      (Ic532c6b85b156f821e0742f47239a65c) +
                      (({q0_1[207],q0_0[207]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[207],q0_0[207]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"

                 if ({q0_1[0],q0_0[0]} != 1 ) begin
                 end
                 if ({q0_1[1],q0_0[1]} != 1 ) begin
                 end
                 if ({q0_1[2],q0_0[2]} != 0 ) begin
                 end
                 if ({q0_1[3],q0_0[3]} != 1 ) begin
                 end
                 if ({q0_1[4],q0_0[4]} != 0 ) begin
                 end
                 if ({q0_1[5],q0_0[5]} != 0 ) begin
                 end
                 if ({q0_1[6],q0_0[6]} != 0 ) begin
                 end
                 if ({q0_1[7],q0_0[7]} != 0 ) begin
                 end
                 if ({q0_1[8],q0_0[8]} != 0 ) begin
                 end
                 if ({q0_1[9],q0_0[9]} != 1 ) begin
                 end
                 if ({q0_1[10],q0_0[10]} != 1 ) begin
                 end
                 if ({q0_1[11],q0_0[11]} != 1 ) begin
                 end
                 if ({q0_1[12],q0_0[12]} != 1 ) begin
                 end
                 if ({q0_1[13],q0_0[13]} != 1 ) begin
                 end
                 if ({q0_1[14],q0_0[14]} != 0 ) begin
                 end
                 if ({q0_1[15],q0_0[15]} != 1 ) begin
                 end
                 if ({q0_1[16],q0_0[16]} != 0 ) begin
                 end
                 if ({q0_1[17],q0_0[17]} != 0 ) begin
                 end
                 if ({q0_1[18],q0_0[18]} != 1 ) begin
                 end
                 if ({q0_1[19],q0_0[19]} != 0 ) begin
                 end
                 if ({q0_1[20],q0_0[20]} != 1 ) begin
                 end
                 if ({q0_1[21],q0_0[21]} != 1 ) begin
                 end
                 if ({q0_1[22],q0_0[22]} != 0 ) begin
                 end
                 if ({q0_1[23],q0_0[23]} != 0 ) begin
                 end
                 if ({q0_1[24],q0_0[24]} != 0 ) begin
                 end
                 if ({q0_1[25],q0_0[25]} != 1 ) begin
                 end
                 if ({q0_1[26],q0_0[26]} != 1 ) begin
                 end
                 if ({q0_1[27],q0_0[27]} != 0 ) begin
                 end
                 if ({q0_1[28],q0_0[28]} != 0 ) begin
                 end
                 if ({q0_1[29],q0_0[29]} != 1 ) begin
                 end
                 if ({q0_1[30],q0_0[30]} != 1 ) begin
                 end
                 if ({q0_1[31],q0_0[31]} != 1 ) begin
                 end
                 if ({q0_1[32],q0_0[32]} != 0 ) begin
                 end
                 if ({q0_1[33],q0_0[33]} != 0 ) begin
                 end
                 if ({q0_1[34],q0_0[34]} != 1 ) begin
                 end
                 if ({q0_1[35],q0_0[35]} != 0 ) begin
                 end
                 if ({q0_1[36],q0_0[36]} != 0 ) begin
                 end
                 if ({q0_1[37],q0_0[37]} != 0 ) begin
                 end
                 if ({q0_1[38],q0_0[38]} != 0 ) begin
                 end
                 if ({q0_1[39],q0_0[39]} != 0 ) begin
                 end
                 if ({q0_1[40],q0_0[40]} != 1 ) begin
                 end
                 if ({q0_1[41],q0_0[41]} != 0 ) begin
                 end
                 if ({q0_1[42],q0_0[42]} != 0 ) begin
                 end
                 if ({q0_1[43],q0_0[43]} != 1 ) begin
                 end
                 if ({q0_1[44],q0_0[44]} != 1 ) begin
                 end
                 if ({q0_1[45],q0_0[45]} != 1 ) begin
                 end
                 if ({q0_1[46],q0_0[46]} != 1 ) begin
                 end
                 if ({q0_1[47],q0_0[47]} != 0 ) begin
                 end
                 if ({q0_1[48],q0_0[48]} != 0 ) begin
                 end
                 if ({q0_1[49],q0_0[49]} != 1 ) begin
                 end
                 if ({q0_1[50],q0_0[50]} != 1 ) begin
                 end
                 if ({q0_1[51],q0_0[51]} != 0 ) begin
                 end
                 if ({q0_1[52],q0_0[52]} != 1 ) begin
                 end
                 if ({q0_1[53],q0_0[53]} != 1 ) begin
                 end
                 if ({q0_1[54],q0_0[54]} != 0 ) begin
                 end
                 if ({q0_1[55],q0_0[55]} != 1 ) begin
                 end
                 if ({q0_1[56],q0_0[56]} != 1 ) begin
                 end
                 if ({q0_1[57],q0_0[57]} != 0 ) begin
                 end
                 if ({q0_1[58],q0_0[58]} != 0 ) begin
                 end
                 if ({q0_1[59],q0_0[59]} != 1 ) begin
                 end
                 if ({q0_1[60],q0_0[60]} != 0 ) begin
                 end
                 if ({q0_1[61],q0_0[61]} != 0 ) begin
                 end
                 if ({q0_1[62],q0_0[62]} != 0 ) begin
                 end
                 if ({q0_1[63],q0_0[63]} != 1 ) begin
                 end
                 if ({q0_1[64],q0_0[64]} != 0 ) begin
                 end
                 if ({q0_1[65],q0_0[65]} != 1 ) begin
                 end
                 if ({q0_1[66],q0_0[66]} != 1 ) begin
                 end
                 if ({q0_1[67],q0_0[67]} != 1 ) begin
                 end
                 if ({q0_1[68],q0_0[68]} != 1 ) begin
                 end
                 if ({q0_1[69],q0_0[69]} != 1 ) begin
                 end
                 if ({q0_1[70],q0_0[70]} != 1 ) begin
                 end
                 if ({q0_1[71],q0_0[71]} != 1 ) begin
                 end
                 if ({q0_1[72],q0_0[72]} != 0 ) begin
                 end
                 if ({q0_1[73],q0_0[73]} != 0 ) begin
                 end
                 if ({q0_1[74],q0_0[74]} != 1 ) begin
                 end
                 if ({q0_1[75],q0_0[75]} != 0 ) begin
                 end
                 if ({q0_1[76],q0_0[76]} != 0 ) begin
                 end
                 if ({q0_1[77],q0_0[77]} != 0 ) begin
                 end
                 if ({q0_1[78],q0_0[78]} != 0 ) begin
                 end
                 if ({q0_1[79],q0_0[79]} != 0 ) begin
                 end
                 if ({q0_1[80],q0_0[80]} != 0 ) begin
                 end
                 if ({q0_1[81],q0_0[81]} != 1 ) begin
                 end
                 if ({q0_1[82],q0_0[82]} != 1 ) begin
                 end
                 if ({q0_1[83],q0_0[83]} != 0 ) begin
                 end
                 if ({q0_1[84],q0_0[84]} != 0 ) begin
                 end
                 if ({q0_1[85],q0_0[85]} != 0 ) begin
                 end
                 if ({q0_1[86],q0_0[86]} != 0 ) begin
                 end
                 if ({q0_1[87],q0_0[87]} != 0 ) begin
                 end
                 if ({q0_1[88],q0_0[88]} != 0 ) begin
                 end
                 if ({q0_1[89],q0_0[89]} != 1 ) begin
                 end
                 if ({q0_1[90],q0_0[90]} != 0 ) begin
                 end
                 if ({q0_1[91],q0_0[91]} != 1 ) begin
                 end
                 if ({q0_1[92],q0_0[92]} != 0 ) begin
                 end
                 if ({q0_1[93],q0_0[93]} != 0 ) begin
                 end
                 if ({q0_1[94],q0_0[94]} != 0 ) begin
                 end
                 if ({q0_1[95],q0_0[95]} != 0 ) begin
                 end
                 if ({q0_1[96],q0_0[96]} != 0 ) begin
                 end
                 if ({q0_1[97],q0_0[97]} != 0 ) begin
                 end
                 if ({q0_1[98],q0_0[98]} != 0 ) begin
                 end
                 if ({q0_1[99],q0_0[99]} != 0 ) begin
                 end
                 if ({q0_1[100],q0_0[100]} != 1 ) begin
                 end
                 if ({q0_1[101],q0_0[101]} != 1 ) begin
                 end
                 if ({q0_1[102],q0_0[102]} != 1 ) begin
                 end
                 if ({q0_1[103],q0_0[103]} != 1 ) begin
                 end
                 if ({q0_1[104],q0_0[104]} != 0 ) begin
                 end
                 if ({q0_1[105],q0_0[105]} != 1 ) begin
                 end
                 if ({q0_1[106],q0_0[106]} != 1 ) begin
                 end
                 if ({q0_1[107],q0_0[107]} != 1 ) begin
                 end
                 if ({q0_1[108],q0_0[108]} != 0 ) begin
                 end
                 if ({q0_1[109],q0_0[109]} != 0 ) begin
                 end
                 if ({q0_1[110],q0_0[110]} != 0 ) begin
                 end
                 if ({q0_1[111],q0_0[111]} != 1 ) begin
                 end
                 if ({q0_1[112],q0_0[112]} != 1 ) begin
                 end
                 if ({q0_1[113],q0_0[113]} != 0 ) begin
                 end
                 if ({q0_1[114],q0_0[114]} != 0 ) begin
                 end
                 if ({q0_1[115],q0_0[115]} != 1 ) begin
                 end
                 if ({q0_1[116],q0_0[116]} != 1 ) begin
                 end
                 if ({q0_1[117],q0_0[117]} != 1 ) begin
                 end
                 if ({q0_1[118],q0_0[118]} != 1 ) begin
                 end
                 if ({q0_1[119],q0_0[119]} != 0 ) begin
                 end
                 if ({q0_1[120],q0_0[120]} != 1 ) begin
                 end
                 if ({q0_1[121],q0_0[121]} != 0 ) begin
                 end
                 if ({q0_1[122],q0_0[122]} != 0 ) begin
                 end
                 if ({q0_1[123],q0_0[123]} != 1 ) begin
                 end
                 if ({q0_1[124],q0_0[124]} != 0 ) begin
                 end
                 if ({q0_1[125],q0_0[125]} != 0 ) begin
                 end
                 if ({q0_1[126],q0_0[126]} != 1 ) begin
                 end
                 if ({q0_1[127],q0_0[127]} != 1 ) begin
                 end
                 if ({q0_1[128],q0_0[128]} != 1 ) begin
                 end
                 if ({q0_1[129],q0_0[129]} != 0 ) begin
                 end
                 if ({q0_1[130],q0_0[130]} != 1 ) begin
                 end
                 if ({q0_1[131],q0_0[131]} != 0 ) begin
                 end
                 if ({q0_1[132],q0_0[132]} != 0 ) begin
                 end
                 if ({q0_1[133],q0_0[133]} != 0 ) begin
                 end
                 if ({q0_1[134],q0_0[134]} != 1 ) begin
                 end
                 if ({q0_1[135],q0_0[135]} != 1 ) begin
                 end
                 if ({q0_1[136],q0_0[136]} != 1 ) begin
                 end
                 if ({q0_1[137],q0_0[137]} != 0 ) begin
                 end
                 if ({q0_1[138],q0_0[138]} != 1 ) begin
                 end
                 if ({q0_1[139],q0_0[139]} != 1 ) begin
                 end
                 if ({q0_1[140],q0_0[140]} != 1 ) begin
                 end
                 if ({q0_1[141],q0_0[141]} != 0 ) begin
                 end
                 if ({q0_1[142],q0_0[142]} != 0 ) begin
                 end
                 if ({q0_1[143],q0_0[143]} != 1 ) begin
                 end
                 if ({q0_1[144],q0_0[144]} != 0 ) begin
                 end
                 if ({q0_1[145],q0_0[145]} != 1 ) begin
                 end
                 if ({q0_1[146],q0_0[146]} != 0 ) begin
                 end
                 if ({q0_1[147],q0_0[147]} != 1 ) begin
                 end
                 if ({q0_1[148],q0_0[148]} != 1 ) begin
                 end
                 if ({q0_1[149],q0_0[149]} != 1 ) begin
                 end
                 if ({q0_1[150],q0_0[150]} != 1 ) begin
                 end
                 if ({q0_1[151],q0_0[151]} != 0 ) begin
                 end
                 if ({q0_1[152],q0_0[152]} != 1 ) begin
                 end
                 if ({q0_1[153],q0_0[153]} != 0 ) begin
                 end
                 if ({q0_1[154],q0_0[154]} != 0 ) begin
                 end
                 if ({q0_1[155],q0_0[155]} != 0 ) begin
                 end
                 if ({q0_1[156],q0_0[156]} != 0 ) begin
                 end
                 if ({q0_1[157],q0_0[157]} != 1 ) begin
                 end
                 if ({q0_1[158],q0_0[158]} != 0 ) begin
                 end
                 if ({q0_1[159],q0_0[159]} != 1 ) begin
                 end
                 if ({q0_1[160],q0_0[160]} != 1 ) begin
                 end
                 if ({q0_1[161],q0_0[161]} != 0 ) begin
                 end
                 if ({q0_1[162],q0_0[162]} != 0 ) begin
                 end
                 if ({q0_1[163],q0_0[163]} != 1 ) begin
                 end
                 if ({q0_1[164],q0_0[164]} != 0 ) begin
                 end
                 if ({q0_1[165],q0_0[165]} != 0 ) begin
                 end
                 if ({q0_1[166],q0_0[166]} != 1 ) begin
                 end
                 if ({q0_1[167],q0_0[167]} != 1 ) begin
                 end
                 if ({q0_1[168],q0_0[168]} != 0 ) begin
                 end
                 if ({q0_1[169],q0_0[169]} != 0 ) begin
                 end
                 if ({q0_1[170],q0_0[170]} != 1 ) begin
                 end
                 if ({q0_1[171],q0_0[171]} != 0 ) begin
                 end
                 if ({q0_1[172],q0_0[172]} != 1 ) begin
                 end
                 if ({q0_1[173],q0_0[173]} != 1 ) begin
                 end
                 if ({q0_1[174],q0_0[174]} != 0 ) begin
                 end
                 if ({q0_1[175],q0_0[175]} != 0 ) begin
                 end
                 if ({q0_1[176],q0_0[176]} != 1 ) begin
                 end
                 if ({q0_1[177],q0_0[177]} != 0 ) begin
                 end
                 if ({q0_1[178],q0_0[178]} != 1 ) begin
                 end
                 if ({q0_1[179],q0_0[179]} != 1 ) begin
                 end
                 if ({q0_1[180],q0_0[180]} != 1 ) begin
                 end
                 if ({q0_1[181],q0_0[181]} != 0 ) begin
                 end
                 if ({q0_1[182],q0_0[182]} != 1 ) begin
                 end
                 if ({q0_1[183],q0_0[183]} != 1 ) begin
                 end
                 if ({q0_1[184],q0_0[184]} != 1 ) begin
                 end
                 if ({q0_1[185],q0_0[185]} != 1 ) begin
                 end
                 if ({q0_1[186],q0_0[186]} != 0 ) begin
                 end
                 if ({q0_1[187],q0_0[187]} != 1 ) begin
                 end
                 if ({q0_1[188],q0_0[188]} != 0 ) begin
                 end
                 if ({q0_1[189],q0_0[189]} != 0 ) begin
                 end
                 if ({q0_1[190],q0_0[190]} != 0 ) begin
                 end
                 if ({q0_1[191],q0_0[191]} != 0 ) begin
                 end
                 if ({q0_1[192],q0_0[192]} != 1 ) begin
                 end
                 if ({q0_1[193],q0_0[193]} != 0 ) begin
                 end
                 if ({q0_1[194],q0_0[194]} != 0 ) begin
                 end
                 if ({q0_1[195],q0_0[195]} != 0 ) begin
                 end
                 if ({q0_1[196],q0_0[196]} != 0 ) begin
                 end
                 if ({q0_1[197],q0_0[197]} != 0 ) begin
                 end
                 if ({q0_1[198],q0_0[198]} != 0 ) begin
                 end
                 if ({q0_1[199],q0_0[199]} != 0 ) begin
                 end
                 if ({q0_1[200],q0_0[200]} != 0 ) begin
                 end
                 if ({q0_1[201],q0_0[201]} != 0 ) begin
                 end
                 if ({q0_1[202],q0_0[202]} != 1 ) begin
                 end
                 if ({q0_1[203],q0_0[203]} != 0 ) begin
                 end
                 if ({q0_1[204],q0_0[204]} != 0 ) begin
                 end
                 if ({q0_1[205],q0_0[205]} != 0 ) begin
                 end
                 if ({q0_1[206],q0_0[206]} != 1 ) begin
                 end
                 if ({q0_1[207],q0_0[207]} != 0 ) begin
                 end


           end

           if (start_d2) begin
            Ic93835a022c46b7aa00a465c407d7da2     <=
                                             wire_qout_00000_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00000 + 1 :
                                             wire_qout_00000_00000
                                             ;

            I92cb615e2c439914e72ce001256518e4  <=  wire_qout_00000_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2e30088bf29cedd7debc15b1e6ec4ada     <=
                                             wire_qout_00000_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00001 + 1 :
                                             wire_qout_00000_00001
                                             ;

            Iad799775eb657f8973e6dfcf70a9875c  <=  wire_qout_00000_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I38f512bfb84094d1e92a10a345d5505f     <=
                                             wire_qout_00000_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00002 + 1 :
                                             wire_qout_00000_00002
                                             ;

            Ifb064c69c7110c014593149ae69c75fb  <=  wire_qout_00000_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1e878f00f056f637625cb013a93325a8     <=
                                             wire_qout_00000_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00003 + 1 :
                                             wire_qout_00000_00003
                                             ;

            I7f7b30f2acbb8e31f50b58096b738254  <=  wire_qout_00000_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I25db27464b31fee41ccd7a3cfe4d403e     <=
                                             wire_qout_00000_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00004 + 1 :
                                             wire_qout_00000_00004
                                             ;

            Iefe4099ff7e457f6b9fefc83e176c1a0  <=  wire_qout_00000_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I19417a224c5cdf1211e9790aa29c4c5c     <=
                                             wire_qout_00000_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00005 + 1 :
                                             wire_qout_00000_00005
                                             ;

            Icddb43f9b760a4597a0bb637fb405616  <=  wire_qout_00000_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I16dcafa854ea9c67d8a080feb2ba9166     <=
                                             wire_qout_00000_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00006 + 1 :
                                             wire_qout_00000_00006
                                             ;

            Ic76e72b434b47c10ebac3fac4ea50bde  <=  wire_qout_00000_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7f63338eee2663fbe61fffd248433310     <=
                                             wire_qout_00000_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00007 + 1 :
                                             wire_qout_00000_00007
                                             ;

            I9eb87e62d23bc87d7cd82c0f329f247f  <=  wire_qout_00000_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icb1e3c56c8729c32d43c69710e345db2     <=
                                             wire_qout_00000_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00008 + 1 :
                                             wire_qout_00000_00008
                                             ;

            I2eac5b39c6f485c9ae0bd341f894633d  <=  wire_qout_00000_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6ece8e3c1e89613879336936f77d732f     <=
                                             wire_qout_00000_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00009 + 1 :
                                             wire_qout_00000_00009
                                             ;

            I76992221b1edff5684c482df7ac4693d  <=  wire_qout_00000_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I72a646ae7e32a16af0f5930a6e95b36a     <=
                                             wire_qout_00000_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00010 + 1 :
                                             wire_qout_00000_00010
                                             ;

            Iada5bc4a51dc1bf57bb9cca11326bdff  <=  wire_qout_00000_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7e72d119dd93a6ab05a23fde0a865866     <=
                                             wire_qout_00000_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00011 + 1 :
                                             wire_qout_00000_00011
                                             ;

            I364ed3f83c49626bc3b939e53524d9c7  <=  wire_qout_00000_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ied4fdf5805039cd2fcd042fd13755fdc     <=
                                             wire_qout_00000_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00012 + 1 :
                                             wire_qout_00000_00012
                                             ;

            Ic2b000c3b2ca3beff2d427caab04701a  <=  wire_qout_00000_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id44c2293b765cff450dd1d747c47c1f3     <=
                                             wire_qout_00000_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00013 + 1 :
                                             wire_qout_00000_00013
                                             ;

            I8e873fb2321eea82bb590a92411e2e2c  <=  wire_qout_00000_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8f4ed02f7aeb823b745040f7f3f43ac7     <=
                                             wire_qout_00000_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00014 + 1 :
                                             wire_qout_00000_00014
                                             ;

            If4cb744ee52b6ae793431cd038069b57  <=  wire_qout_00000_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6488b9b8f405d7d81a4874fab2678102     <=
                                             wire_qout_00000_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00015 + 1 :
                                             wire_qout_00000_00015
                                             ;

            I7741e239c16828889d488cc87647c154  <=  wire_qout_00000_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifff612d16828ec907a348479e19ddf31     <=
                                             wire_qout_00000_00016[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00016 + 1 :
                                             wire_qout_00000_00016
                                             ;

            I7979161aa1e2262ebea862004c387697  <=  wire_qout_00000_00016[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I268262076f22bc6b1507bc8f91b98a0a     <=
                                             wire_qout_00000_00017[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00017 + 1 :
                                             wire_qout_00000_00017
                                             ;

            Ic62fc602da3d16fe13d03a49a21269d0  <=  wire_qout_00000_00017[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If1f732841adb7c0cad1ba37c0f5fd517     <=
                                             wire_qout_00000_00018[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00018 + 1 :
                                             wire_qout_00000_00018
                                             ;

            I94009bb7239be96243902ab0f0abea7e  <=  wire_qout_00000_00018[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0df8a24f31c027756d248c3bd1b9bf7b     <=
                                             wire_qout_00000_00019[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00019 + 1 :
                                             wire_qout_00000_00019
                                             ;

            Iae7b72abf4d3c536330a229e3836b441  <=  wire_qout_00000_00019[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8ef901e733b12e76412eb36684e2b575     <=
                                             wire_qout_00000_00020[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00020 + 1 :
                                             wire_qout_00000_00020
                                             ;

            Ie5d9cc18b2dd300132470f206452ff17  <=  wire_qout_00000_00020[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia48916a02f68b1b8f5fc7fece04677bb     <=
                                             wire_qout_00000_00021[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00000_00021 + 1 :
                                             wire_qout_00000_00021
                                             ;

            I7c791c854d0bc28e8dd787545f8fbda0  <=  wire_qout_00000_00021[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia37409944d9fdd3b16e7007e13d82a79     <=
                                             wire_qout_00001_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00000 + 1 :
                                             wire_qout_00001_00000
                                             ;

            I5b177dd5c14ad082516b47f550875682  <=  wire_qout_00001_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idd65f149afe9d5f63ddaf34b82b11e95     <=
                                             wire_qout_00001_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00001 + 1 :
                                             wire_qout_00001_00001
                                             ;

            I55e4ad2d71a29ad63b4999d64ac0dc4f  <=  wire_qout_00001_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If2886d560854faed32ebd8e33d868973     <=
                                             wire_qout_00001_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00002 + 1 :
                                             wire_qout_00001_00002
                                             ;

            I59c5da6338f431a626c86a065a355c35  <=  wire_qout_00001_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I77778118bb3ea900c080754ff4c49c26     <=
                                             wire_qout_00001_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00003 + 1 :
                                             wire_qout_00001_00003
                                             ;

            Ia098bbeda8b755ece6b88eac83d03e55  <=  wire_qout_00001_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7292ed752d8741594d757730950feea4     <=
                                             wire_qout_00001_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00004 + 1 :
                                             wire_qout_00001_00004
                                             ;

            Ie7470dd75b54d14038de19e4d3043ba9  <=  wire_qout_00001_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I68cfd7868e061793ee8a41e69e80219b     <=
                                             wire_qout_00001_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00005 + 1 :
                                             wire_qout_00001_00005
                                             ;

            Ie95662d4faf6b5a4cd5ecfa41697b983  <=  wire_qout_00001_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I667ead814b303fca64ef047bb8246b19     <=
                                             wire_qout_00001_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00006 + 1 :
                                             wire_qout_00001_00006
                                             ;

            Ia1b617e3d141263b51e58c5ef0bd7a89  <=  wire_qout_00001_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4f25c7edb12e868cb5532e42b4ba5133     <=
                                             wire_qout_00001_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00007 + 1 :
                                             wire_qout_00001_00007
                                             ;

            If9a5d830e3ade0fd96b98f5949f165f0  <=  wire_qout_00001_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5aed2d82717f359bb5ac5a0ab91b7beb     <=
                                             wire_qout_00001_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00008 + 1 :
                                             wire_qout_00001_00008
                                             ;

            Id3de87169c440f95d406693ef77cacd6  <=  wire_qout_00001_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I92835fd54631deaefa7b214e2c4b9bff     <=
                                             wire_qout_00001_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00009 + 1 :
                                             wire_qout_00001_00009
                                             ;

            I3751f191f5009322acb7c9be4f8d7129  <=  wire_qout_00001_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I67e067da565635fcff166e3a7d0c446b     <=
                                             wire_qout_00001_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00010 + 1 :
                                             wire_qout_00001_00010
                                             ;

            Ic1927bb3335f6a28c0816eba12d3975e  <=  wire_qout_00001_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifdb0f307b1b9458c0487a1574ccc094b     <=
                                             wire_qout_00001_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00011 + 1 :
                                             wire_qout_00001_00011
                                             ;

            Ia659126b51468cfef48c97a135a71500  <=  wire_qout_00001_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5c6b7d143e42fd3b8bcdb7d7ed4da2c2     <=
                                             wire_qout_00001_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00012 + 1 :
                                             wire_qout_00001_00012
                                             ;

            I3c3c22bf63e55a81ae91b1dd1ef615a0  <=  wire_qout_00001_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie679a21d0136a08cc5e6526e9f8d1843     <=
                                             wire_qout_00001_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00013 + 1 :
                                             wire_qout_00001_00013
                                             ;

            Ia62832d325f86160285c4d1a790a32cb  <=  wire_qout_00001_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I611942a72a5e12f6afaea6bde6699ef6     <=
                                             wire_qout_00001_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00014 + 1 :
                                             wire_qout_00001_00014
                                             ;

            I83c7d177eec2dad0a924557cdc91ba77  <=  wire_qout_00001_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ica9883c97f823a4491cbee5b45c43590     <=
                                             wire_qout_00001_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00015 + 1 :
                                             wire_qout_00001_00015
                                             ;

            I7050adb9d06f767549b7f35c4679e391  <=  wire_qout_00001_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8e6addfc61f5bfb7af74fc2993639565     <=
                                             wire_qout_00001_00016[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00016 + 1 :
                                             wire_qout_00001_00016
                                             ;

            I04aacd95d9e44657f616e01c9053f0fb  <=  wire_qout_00001_00016[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9d53619f10e2a426f7297bbf7c81158a     <=
                                             wire_qout_00001_00017[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00017 + 1 :
                                             wire_qout_00001_00017
                                             ;

            I2ff317d57f59747c4524ef4278d51092  <=  wire_qout_00001_00017[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8a055c27778913287ad951183fa0d4d6     <=
                                             wire_qout_00001_00018[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00018 + 1 :
                                             wire_qout_00001_00018
                                             ;

            I8bd2a9d90074500698b302cb8db7f03a  <=  wire_qout_00001_00018[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8f6ae5c80bb2f50084b5f5ee5ab0ffc3     <=
                                             wire_qout_00001_00019[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00019 + 1 :
                                             wire_qout_00001_00019
                                             ;

            I3b8cdfb1440732ce98cd1676e05a2af1  <=  wire_qout_00001_00019[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3db8b3a342e8e2f13a448246aa001c2f     <=
                                             wire_qout_00001_00020[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00020 + 1 :
                                             wire_qout_00001_00020
                                             ;

            I671de3d408b5b783541663c7f1e3a6fa  <=  wire_qout_00001_00020[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibbee0996ea0f5e16b1f711345be7f2ae     <=
                                             wire_qout_00001_00021[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00001_00021 + 1 :
                                             wire_qout_00001_00021
                                             ;

            I446857735e680cae93a24dccb59b1924  <=  wire_qout_00001_00021[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idb777f1eb4c3cbba103b9b43f948ccf9     <=
                                             wire_qout_00002_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00000 + 1 :
                                             wire_qout_00002_00000
                                             ;

            I77b05a8aa92c66a235195a66dc13c0cc  <=  wire_qout_00002_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id5e46b1f8844c7587f99d22170581a24     <=
                                             wire_qout_00002_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00001 + 1 :
                                             wire_qout_00002_00001
                                             ;

            Ie92110d19f4886cdfcfacd0920c06a4e  <=  wire_qout_00002_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I67aadabd3cf49456cace7392a1e7a35a     <=
                                             wire_qout_00002_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00002 + 1 :
                                             wire_qout_00002_00002
                                             ;

            I36ba87b69b5b9dd919319230f697dfad  <=  wire_qout_00002_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id5635595d6b7b6dd7e6d510a27ad6702     <=
                                             wire_qout_00002_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00003 + 1 :
                                             wire_qout_00002_00003
                                             ;

            Id20e72ac258d1d1b6cdca1e6c9e3596d  <=  wire_qout_00002_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ice783314a4868f0bba8bc3c5e3b65ae4     <=
                                             wire_qout_00002_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00004 + 1 :
                                             wire_qout_00002_00004
                                             ;

            Ifc34f5d6b7a7d0533439794958959856  <=  wire_qout_00002_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib2d9b7f58cf571b904be02e6073f9b94     <=
                                             wire_qout_00002_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00005 + 1 :
                                             wire_qout_00002_00005
                                             ;

            I849ee5d34760be03d4285185136aa52e  <=  wire_qout_00002_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I61b6effae91ae4bdcce4550eb5cf0796     <=
                                             wire_qout_00002_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00006 + 1 :
                                             wire_qout_00002_00006
                                             ;

            Ia3559d98eb372b7307f30ad1f7c4c7cd  <=  wire_qout_00002_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If5cf6e81b0e3b77f6a45f2555201acc2     <=
                                             wire_qout_00002_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00007 + 1 :
                                             wire_qout_00002_00007
                                             ;

            I7332e088bbff69db19c62685e033d26a  <=  wire_qout_00002_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I62fae5bf51588f28c3521715b834909d     <=
                                             wire_qout_00002_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00008 + 1 :
                                             wire_qout_00002_00008
                                             ;

            I44daa5992b00e7af19adbee70bf01f2b  <=  wire_qout_00002_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If5cbdab78a4cf86b6285a400d0e0ac90     <=
                                             wire_qout_00002_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00009 + 1 :
                                             wire_qout_00002_00009
                                             ;

            Ie517386cb5832e406fefc5e85eb2e7d1  <=  wire_qout_00002_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6e481cc49441c08bcd9fdcabbe90a000     <=
                                             wire_qout_00002_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00010 + 1 :
                                             wire_qout_00002_00010
                                             ;

            I9b096ce09467c10f448496fda13987d2  <=  wire_qout_00002_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3aa663be3dd604564ef68b9a2b9d7319     <=
                                             wire_qout_00002_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00011 + 1 :
                                             wire_qout_00002_00011
                                             ;

            If1c0a3726041f70e508d68cbf6e40e04  <=  wire_qout_00002_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8031632ee8700c63c207e2d6a6bdb630     <=
                                             wire_qout_00002_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00012 + 1 :
                                             wire_qout_00002_00012
                                             ;

            Iaf36ce8598a29573979c683a5e2cf9fd  <=  wire_qout_00002_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If9be2701858da0bdffbf2dff7bcfd7e1     <=
                                             wire_qout_00002_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00013 + 1 :
                                             wire_qout_00002_00013
                                             ;

            Ice82cfe55a5f226746e59e5c8beb46be  <=  wire_qout_00002_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ief209532f4cbf1c6a41bea414577f825     <=
                                             wire_qout_00002_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00014 + 1 :
                                             wire_qout_00002_00014
                                             ;

            Iea1297491d1dfe98f395d8c73808a893  <=  wire_qout_00002_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1c8953ad3f64f3c3cc506808aad29dab     <=
                                             wire_qout_00002_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00015 + 1 :
                                             wire_qout_00002_00015
                                             ;

            If43dd31198c8a0da6fabd194cf13bb70  <=  wire_qout_00002_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1b519d88bbf86cfb080a50ea0480a128     <=
                                             wire_qout_00002_00016[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00016 + 1 :
                                             wire_qout_00002_00016
                                             ;

            Ibeb8c72b90b50c6897224ca1a792fa56  <=  wire_qout_00002_00016[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5b8258f35d889071109216b464abb2a4     <=
                                             wire_qout_00002_00017[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00017 + 1 :
                                             wire_qout_00002_00017
                                             ;

            I8e87530a131b5a73cad6df68b9e4967f  <=  wire_qout_00002_00017[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id9681d4e0e4d375f9279de115a4337a3     <=
                                             wire_qout_00002_00018[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00018 + 1 :
                                             wire_qout_00002_00018
                                             ;

            Idf8d15c7bd7705b9aafbda09c3a5b46c  <=  wire_qout_00002_00018[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib42144ece00b82debd70011724a29c91     <=
                                             wire_qout_00002_00019[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00019 + 1 :
                                             wire_qout_00002_00019
                                             ;

            I2aea17846a53e2eb2968581ee2c48226  <=  wire_qout_00002_00019[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic5717058a1815f63f164de1b1defe8cb     <=
                                             wire_qout_00002_00020[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00020 + 1 :
                                             wire_qout_00002_00020
                                             ;

            I169d8f2bb5fde5b202b4239b7a7f1ed5  <=  wire_qout_00002_00020[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iea41672f012f225d64d9c75b198c812f     <=
                                             wire_qout_00002_00021[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00002_00021 + 1 :
                                             wire_qout_00002_00021
                                             ;

            I40a223380fb4414a3f26a08cb90025ec  <=  wire_qout_00002_00021[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7a070bd014e1d2c5e55e5fcba88a5664     <=
                                             wire_qout_00003_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00000 + 1 :
                                             wire_qout_00003_00000
                                             ;

            Ie117f6ec475f5d6444998af151ce4e69  <=  wire_qout_00003_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4a0a8b28429b708363458c74230b0fc2     <=
                                             wire_qout_00003_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00001 + 1 :
                                             wire_qout_00003_00001
                                             ;

            If7f3174da35dd39af7f4792aaa649bf1  <=  wire_qout_00003_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If585e4075ac1740f3b141ae6a50200f7     <=
                                             wire_qout_00003_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00002 + 1 :
                                             wire_qout_00003_00002
                                             ;

            I719a892ad54e63b217c7271741b29cc5  <=  wire_qout_00003_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie1a68cf09bb21a1629369fde87f51bea     <=
                                             wire_qout_00003_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00003 + 1 :
                                             wire_qout_00003_00003
                                             ;

            I4acf6d84471cd237f65c9b2391b7a20c  <=  wire_qout_00003_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I72b8547125d0ad6c1ad39a68b55c818c     <=
                                             wire_qout_00003_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00004 + 1 :
                                             wire_qout_00003_00004
                                             ;

            I7a387a1f887c32e9d0f8e89912a8618c  <=  wire_qout_00003_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie14ba4a8657740f9a8d057258db2cb09     <=
                                             wire_qout_00003_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00005 + 1 :
                                             wire_qout_00003_00005
                                             ;

            Ib862ac63c230ccde7fae0e62f9d047fe  <=  wire_qout_00003_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I27490a69fb2a1f6f298639254c37cf9e     <=
                                             wire_qout_00003_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00006 + 1 :
                                             wire_qout_00003_00006
                                             ;

            I8f1a8a22637d37c3692e808d5eb3d543  <=  wire_qout_00003_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I49b9c212fbe74a5dd8b087e417296186     <=
                                             wire_qout_00003_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00007 + 1 :
                                             wire_qout_00003_00007
                                             ;

            I6f420c64640dfb0c001f57df7e3b4504  <=  wire_qout_00003_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0a8e6f5cc8b6ea599b7605abe6479bec     <=
                                             wire_qout_00003_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00008 + 1 :
                                             wire_qout_00003_00008
                                             ;

            I3600031716c2b4e21c9f577d34e033dc  <=  wire_qout_00003_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib6d94b34d3886717e4016fec196f277f     <=
                                             wire_qout_00003_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00009 + 1 :
                                             wire_qout_00003_00009
                                             ;

            I002820a37fa7c6c504c487df4368e2cf  <=  wire_qout_00003_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id7e53d36da7171e036ebfc984dbcea6e     <=
                                             wire_qout_00003_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00010 + 1 :
                                             wire_qout_00003_00010
                                             ;

            I8a4c1f23212ff846400651b100add502  <=  wire_qout_00003_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2ec254d80fd0683d782302cf3839559b     <=
                                             wire_qout_00003_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00011 + 1 :
                                             wire_qout_00003_00011
                                             ;

            Ice1ce5b4c30841dd92268559ebadafcf  <=  wire_qout_00003_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibbedaef61051d5df82cd6d55e05c80da     <=
                                             wire_qout_00003_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00012 + 1 :
                                             wire_qout_00003_00012
                                             ;

            I3eeeb1949945032d6c1759875426b733  <=  wire_qout_00003_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I501336bb7ba172c05dd5840036e6228c     <=
                                             wire_qout_00003_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00013 + 1 :
                                             wire_qout_00003_00013
                                             ;

            I384d5377ee6b8f7eb2db23a2e444ddbc  <=  wire_qout_00003_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8e5c4c6c63e42054359cee697cc0d026     <=
                                             wire_qout_00003_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00014 + 1 :
                                             wire_qout_00003_00014
                                             ;

            I30d615203b697787ead37394953925cc  <=  wire_qout_00003_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id3daa6db921871b752bf92366446afcc     <=
                                             wire_qout_00003_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00015 + 1 :
                                             wire_qout_00003_00015
                                             ;

            Ib16548d471f0a4f4625852ea04335dcc  <=  wire_qout_00003_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id8367ec60787bfad0da8aa76c6ed8ddb     <=
                                             wire_qout_00003_00016[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00016 + 1 :
                                             wire_qout_00003_00016
                                             ;

            I0987c561670b7b2b6683303c1be39561  <=  wire_qout_00003_00016[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I533649312ec995f1f9e514c59a8675b1     <=
                                             wire_qout_00003_00017[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00017 + 1 :
                                             wire_qout_00003_00017
                                             ;

            I2bdf4736022e5da7294a0e851006a124  <=  wire_qout_00003_00017[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0621d0b2c83e70b4afd65eb9dca4b514     <=
                                             wire_qout_00003_00018[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00018 + 1 :
                                             wire_qout_00003_00018
                                             ;

            Ic6fd9592d2ffcb8f4ca83c6f0bd19975  <=  wire_qout_00003_00018[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2ae01892a3cd0432618d7280b31daddb     <=
                                             wire_qout_00003_00019[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00019 + 1 :
                                             wire_qout_00003_00019
                                             ;

            I14bf11ad80890227e47fda26ae1b9c24  <=  wire_qout_00003_00019[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5ed8a2f30bd2ea269341c2267ae3fe83     <=
                                             wire_qout_00003_00020[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00020 + 1 :
                                             wire_qout_00003_00020
                                             ;

            I8ca17b6cf35e1b1f8f601604575d3f27  <=  wire_qout_00003_00020[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2c819e7f62c0dc0aac650074b203163b     <=
                                             wire_qout_00003_00021[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00003_00021 + 1 :
                                             wire_qout_00003_00021
                                             ;

            I275cd09649a750edb8ae8313e4e1e279  <=  wire_qout_00003_00021[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I30e20b58913d6fbe5817e1956ba8e570     <=
                                             wire_qout_00004_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00000 + 1 :
                                             wire_qout_00004_00000
                                             ;

            I7d6a6026eb3c4d06e682523424f9628f  <=  wire_qout_00004_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1b922bed7f3c4a6705f3ce7a885a68cd     <=
                                             wire_qout_00004_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00001 + 1 :
                                             wire_qout_00004_00001
                                             ;

            Ia0c192e590d8c914555b434ce5a634a8  <=  wire_qout_00004_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2f65f0917713ecc8585392d3b557c1bf     <=
                                             wire_qout_00004_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00002 + 1 :
                                             wire_qout_00004_00002
                                             ;

            Ic98c8641d2022080297c54ff2539e75d  <=  wire_qout_00004_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3301533e7d9e527118a67c462f1b4357     <=
                                             wire_qout_00004_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00003 + 1 :
                                             wire_qout_00004_00003
                                             ;

            I87f34821cd0b58f8855b25c75f2dd32d  <=  wire_qout_00004_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I52a88bdb1f03da82730f7579b7b5305d     <=
                                             wire_qout_00004_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00004 + 1 :
                                             wire_qout_00004_00004
                                             ;

            I87211ac14d832ad3205d47fb83cf256a  <=  wire_qout_00004_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I644c730662b3725d26cd46fb46106104     <=
                                             wire_qout_00004_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00005 + 1 :
                                             wire_qout_00004_00005
                                             ;

            Ib81431cfb3b281555fa7e5b4582a2524  <=  wire_qout_00004_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3da3e36c76c4123bec6879bccb39e933     <=
                                             wire_qout_00004_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00006 + 1 :
                                             wire_qout_00004_00006
                                             ;

            I835b902949c2c4c09b757d4d35574a76  <=  wire_qout_00004_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iebde55cddc8170f7dd8855ea55eff0ce     <=
                                             wire_qout_00004_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00007 + 1 :
                                             wire_qout_00004_00007
                                             ;

            I8510240df7dc41f85ad58a39868a1fd7  <=  wire_qout_00004_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie673e2d92a7090b2fa1c5e14a2e03be3     <=
                                             wire_qout_00004_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00008 + 1 :
                                             wire_qout_00004_00008
                                             ;

            I1b6abc8fbab3849b285e9f88a4fe867b  <=  wire_qout_00004_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If90afe75714f8660ad0eb9f9ea06cd6b     <=
                                             wire_qout_00004_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00009 + 1 :
                                             wire_qout_00004_00009
                                             ;

            Ied638fee34f8baed4154b0b72e43a21e  <=  wire_qout_00004_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifd96e3a6e0050c30a4308328cfecb21f     <=
                                             wire_qout_00004_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00010 + 1 :
                                             wire_qout_00004_00010
                                             ;

            I14fa7aebb608d4a3d67176ba27d34d9a  <=  wire_qout_00004_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I68b92cc2d83e9a718edd2aea82314016     <=
                                             wire_qout_00004_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00011 + 1 :
                                             wire_qout_00004_00011
                                             ;

            Iad90879acba3fc2101829549264960f3  <=  wire_qout_00004_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6bdbb92363f0e072ed04654e9aad17a5     <=
                                             wire_qout_00004_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00012 + 1 :
                                             wire_qout_00004_00012
                                             ;

            Ife0952b85f14a960007b67646b0cd969  <=  wire_qout_00004_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I87a4267db59b97ef1b9bca8743cb0322     <=
                                             wire_qout_00004_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00013 + 1 :
                                             wire_qout_00004_00013
                                             ;

            If876ca6a14ffb4323503ed46666bc25f  <=  wire_qout_00004_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I44eacb2bea725efab7c0dd560279f0f8     <=
                                             wire_qout_00004_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00014 + 1 :
                                             wire_qout_00004_00014
                                             ;

            If2dfcbf493b761fb5d7c622e739b23f3  <=  wire_qout_00004_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I87a2736466c5ee62b7cc55f17e715ffa     <=
                                             wire_qout_00004_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00015 + 1 :
                                             wire_qout_00004_00015
                                             ;

            I2c8f4a147b363d9c5ef0e080d9a9ed40  <=  wire_qout_00004_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7a66c7713ba126fdc24940cd92f7e10b     <=
                                             wire_qout_00004_00016[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00016 + 1 :
                                             wire_qout_00004_00016
                                             ;

            I485f9d1104a965d5d035feef912a2ca8  <=  wire_qout_00004_00016[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1f11c579f34c41aade41c53f53468057     <=
                                             wire_qout_00004_00017[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00017 + 1 :
                                             wire_qout_00004_00017
                                             ;

            I10fca5f2cbf5e2bc3433c0dda579a051  <=  wire_qout_00004_00017[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I651a438f70583d476ae10f066e035435     <=
                                             wire_qout_00004_00018[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00018 + 1 :
                                             wire_qout_00004_00018
                                             ;

            If8572800d5d80cc92dd917b60447b63b  <=  wire_qout_00004_00018[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibdf17fa73794c846e15fe0a915b071e5     <=
                                             wire_qout_00004_00019[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00019 + 1 :
                                             wire_qout_00004_00019
                                             ;

            I24645082ef16129eed1c574f5fc601ca  <=  wire_qout_00004_00019[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I76d3221fbcefc0ee08655f7ba4919f3c     <=
                                             wire_qout_00004_00020[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00020 + 1 :
                                             wire_qout_00004_00020
                                             ;

            I207a0f6184a0b3be71766a8b47ea5535  <=  wire_qout_00004_00020[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3458f69c90ea8b20b3d1f67e9a13ec2e     <=
                                             wire_qout_00004_00021[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00021 + 1 :
                                             wire_qout_00004_00021
                                             ;

            I5cac08dabbb6de3b01c821d4db93a8e3  <=  wire_qout_00004_00021[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia2d6e9e1e92a30c7028af50ddfbb9bf9     <=
                                             wire_qout_00004_00022[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00004_00022 + 1 :
                                             wire_qout_00004_00022
                                             ;

            Ibe6b8c57d7ff47b6fdad5fadf1f6b841  <=  wire_qout_00004_00022[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I66c91b5133d9812a03daecc0b14211f8     <=
                                             wire_qout_00005_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00000 + 1 :
                                             wire_qout_00005_00000
                                             ;

            I477326720157df2503149125a43ee987  <=  wire_qout_00005_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifb5986949e88167526d9fcfe07b417ca     <=
                                             wire_qout_00005_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00001 + 1 :
                                             wire_qout_00005_00001
                                             ;

            I2c741a5fed7d88e9bdd6b7459feac649  <=  wire_qout_00005_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iedada801ca6cd173ee523ef335e91ff6     <=
                                             wire_qout_00005_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00002 + 1 :
                                             wire_qout_00005_00002
                                             ;

            I17a6511072c7fb4846be5844decf17d6  <=  wire_qout_00005_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4e2722e547586da7565b2d91a7fc91e7     <=
                                             wire_qout_00005_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00003 + 1 :
                                             wire_qout_00005_00003
                                             ;

            I5ebc3047985651f4b9a957d502a97e95  <=  wire_qout_00005_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib321a8ceda62c64ab25dc1c718301bda     <=
                                             wire_qout_00005_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00004 + 1 :
                                             wire_qout_00005_00004
                                             ;

            Ifa09fc1b009d073d5a9973b430c63469  <=  wire_qout_00005_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I58daeebec4873e6c1c07c090ff81235c     <=
                                             wire_qout_00005_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00005 + 1 :
                                             wire_qout_00005_00005
                                             ;

            Ie6212a29c7c6b035cfff4c869f945b68  <=  wire_qout_00005_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3f103fbbe49c86c9db46129bd4632cab     <=
                                             wire_qout_00005_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00006 + 1 :
                                             wire_qout_00005_00006
                                             ;

            If343015b4815b01dae88bbb6f2017b3d  <=  wire_qout_00005_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id6697ca17f1bd6ddd112951b9d89a8ea     <=
                                             wire_qout_00005_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00007 + 1 :
                                             wire_qout_00005_00007
                                             ;

            Ia0116a3cebf94318ed5b287960957ad6  <=  wire_qout_00005_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I445ede2983c7470b4418a2ec0cbbd5e1     <=
                                             wire_qout_00005_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00008 + 1 :
                                             wire_qout_00005_00008
                                             ;

            Id75c23e80cdf25d883806ed20d4ae783  <=  wire_qout_00005_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I034e56cd77ee400ed81b78177b202930     <=
                                             wire_qout_00005_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00009 + 1 :
                                             wire_qout_00005_00009
                                             ;

            I1b43f29e0ddb72467befd6f3a9c1c829  <=  wire_qout_00005_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I08edadbd9366786f96b44268d096b4aa     <=
                                             wire_qout_00005_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00010 + 1 :
                                             wire_qout_00005_00010
                                             ;

            I3fd0fa3b774d30a267d61e9427d09f3f  <=  wire_qout_00005_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8f86a7af86eb04c5df18e09888cdce7b     <=
                                             wire_qout_00005_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00011 + 1 :
                                             wire_qout_00005_00011
                                             ;

            I2eb08ebaa07a1004638cdd61a7209b7d  <=  wire_qout_00005_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic00d037a11f8a27ab34e4daab8c9c2e6     <=
                                             wire_qout_00005_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00012 + 1 :
                                             wire_qout_00005_00012
                                             ;

            I258c45897919cec5c6acaddee7f3a41b  <=  wire_qout_00005_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4d95ceccc6c3ad37f13c98339c59e5c4     <=
                                             wire_qout_00005_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00013 + 1 :
                                             wire_qout_00005_00013
                                             ;

            Ib42d37576e3aff3d205f1f8822cc58b5  <=  wire_qout_00005_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1ea967d377f462a0e06d7d0d4d95b342     <=
                                             wire_qout_00005_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00014 + 1 :
                                             wire_qout_00005_00014
                                             ;

            I1c2ee281cd47a8414851c5e1c758ea65  <=  wire_qout_00005_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib0feec63123e66bd6ad6935e9b7fa6bf     <=
                                             wire_qout_00005_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00015 + 1 :
                                             wire_qout_00005_00015
                                             ;

            Ie644d131c4f2c603e8e64c5581fdf822  <=  wire_qout_00005_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7d120060ddae9ff8f7206b3ef63eda50     <=
                                             wire_qout_00005_00016[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00016 + 1 :
                                             wire_qout_00005_00016
                                             ;

            I9b76f0121a3f7e887e7121db50024ab4  <=  wire_qout_00005_00016[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib47f8f72386e2e65a88fbadd3a705225     <=
                                             wire_qout_00005_00017[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00017 + 1 :
                                             wire_qout_00005_00017
                                             ;

            I9eaf4e9ebe07717503ff69b51f0e1905  <=  wire_qout_00005_00017[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4e0efc35346e2934f5bb4c34a4bc5f90     <=
                                             wire_qout_00005_00018[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00018 + 1 :
                                             wire_qout_00005_00018
                                             ;

            Icb0841ecf142687c3aa23e68f01c927c  <=  wire_qout_00005_00018[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3ca1014802f58087e3434a1e0df19c01     <=
                                             wire_qout_00005_00019[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00019 + 1 :
                                             wire_qout_00005_00019
                                             ;

            Ie8c0fac00a9de74870e59cbf9e87a39b  <=  wire_qout_00005_00019[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I688a3879b7be1544e6f94b4221c03213     <=
                                             wire_qout_00005_00020[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00020 + 1 :
                                             wire_qout_00005_00020
                                             ;

            Iae5d6faac1f5685cb1d400ee2b1d85e0  <=  wire_qout_00005_00020[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic22988138610c8671ec342f65f34c7ae     <=
                                             wire_qout_00005_00021[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00021 + 1 :
                                             wire_qout_00005_00021
                                             ;

            Ib62b02ddf0f57bee49838d19783ef6c3  <=  wire_qout_00005_00021[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0b85fdd83569e5cbb7d71eed50cb32fd     <=
                                             wire_qout_00005_00022[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00005_00022 + 1 :
                                             wire_qout_00005_00022
                                             ;

            Ibd59d0e5a062f149bd0e91ba76985a13  <=  wire_qout_00005_00022[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idf55390c11e5b41ebc2a28e0af109913     <=
                                             wire_qout_00006_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00000 + 1 :
                                             wire_qout_00006_00000
                                             ;

            I876fdba97e755b74532f7ab191fbac14  <=  wire_qout_00006_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6b48935ea25672ee9a42f49eae9e519f     <=
                                             wire_qout_00006_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00001 + 1 :
                                             wire_qout_00006_00001
                                             ;

            I8edf1a08ef943f06ee28771c6e140e28  <=  wire_qout_00006_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6a9e6c39c20e45773dab7823a7ff9486     <=
                                             wire_qout_00006_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00002 + 1 :
                                             wire_qout_00006_00002
                                             ;

            I7e12ad8a8ef857e02f4563b2f3a7f0ca  <=  wire_qout_00006_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I42907182010c5889ddb7a700ead16525     <=
                                             wire_qout_00006_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00003 + 1 :
                                             wire_qout_00006_00003
                                             ;

            I17b3a9df6752da6cc987e902e6bbad48  <=  wire_qout_00006_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib6c26f3e3358cc2ed6fbda83eabd4bd3     <=
                                             wire_qout_00006_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00004 + 1 :
                                             wire_qout_00006_00004
                                             ;

            I487496233a32f657171b3789590d0522  <=  wire_qout_00006_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia50d85808790790450f87a5246874b3f     <=
                                             wire_qout_00006_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00005 + 1 :
                                             wire_qout_00006_00005
                                             ;

            Ie34534dfd435b3d1cf35e82ca71e83ba  <=  wire_qout_00006_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id4a1744702d7808a80bc40697c864765     <=
                                             wire_qout_00006_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00006 + 1 :
                                             wire_qout_00006_00006
                                             ;

            I0e8679271ba733bb87c44b6b9f0b6ed2  <=  wire_qout_00006_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0cf3d2f3e6793a2dcf15949da16ad28d     <=
                                             wire_qout_00006_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00007 + 1 :
                                             wire_qout_00006_00007
                                             ;

            Ic14760b65c6fe150c3c48e64389a41d8  <=  wire_qout_00006_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I90bd9107f4c931fa1ccb92998ea8cdeb     <=
                                             wire_qout_00006_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00008 + 1 :
                                             wire_qout_00006_00008
                                             ;

            Ied6c684cdd280b41ffab93a026d27282  <=  wire_qout_00006_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ida1c729e6bfcec2c31a92aa9002f2c68     <=
                                             wire_qout_00006_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00009 + 1 :
                                             wire_qout_00006_00009
                                             ;

            Id0f4dbb72da33748d8baf723c5a32567  <=  wire_qout_00006_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib848feeccd0ea78ebc8ba8368534c3d1     <=
                                             wire_qout_00006_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00010 + 1 :
                                             wire_qout_00006_00010
                                             ;

            Ib0bb71b1f8829347b3a9a7543f9dd964  <=  wire_qout_00006_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icc11970bbae3adcfa33a0e5dba3e78f4     <=
                                             wire_qout_00006_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00011 + 1 :
                                             wire_qout_00006_00011
                                             ;

            I47cbb92d2284aef7b9e56e88f0ba6f7e  <=  wire_qout_00006_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I86bb4ef4bdd7af8861280ef30fbeeeea     <=
                                             wire_qout_00006_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00012 + 1 :
                                             wire_qout_00006_00012
                                             ;

            Ic69094123b75ae36e3e54f179a9f2cb5  <=  wire_qout_00006_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7e0c259c6c7bacdff5edc44a22e005ba     <=
                                             wire_qout_00006_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00013 + 1 :
                                             wire_qout_00006_00013
                                             ;

            I07abbbd75d91018ac53f53e64cffafb9  <=  wire_qout_00006_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I897ddba059b27f7ed009b0cb70cfb46f     <=
                                             wire_qout_00006_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00014 + 1 :
                                             wire_qout_00006_00014
                                             ;

            Ib02268d5048c7c8e83118070e927453f  <=  wire_qout_00006_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4496243eb0542a514b551b4d09bffd7d     <=
                                             wire_qout_00006_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00015 + 1 :
                                             wire_qout_00006_00015
                                             ;

            Idc2a9c6dd8d2aa912548c918c8a488f4  <=  wire_qout_00006_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic931fb08b2e8441321ebdeed84576a0d     <=
                                             wire_qout_00006_00016[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00016 + 1 :
                                             wire_qout_00006_00016
                                             ;

            I5ad7eb9d3ce7c712515254f892d1670d  <=  wire_qout_00006_00016[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ieb6af5390b98e893ee05a939c16d2ffd     <=
                                             wire_qout_00006_00017[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00017 + 1 :
                                             wire_qout_00006_00017
                                             ;

            Ife25829fb3c5023b7d69bbaadf9cf77e  <=  wire_qout_00006_00017[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic2a54bad4c5a8885dd24b8687c6db0de     <=
                                             wire_qout_00006_00018[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00018 + 1 :
                                             wire_qout_00006_00018
                                             ;

            I8b2a79aa4ac88e6b4ca8188a7852022e  <=  wire_qout_00006_00018[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6ecbad763d2b48b78a0584beaefc78ee     <=
                                             wire_qout_00006_00019[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00019 + 1 :
                                             wire_qout_00006_00019
                                             ;

            I081e2595b18f306a74d070203447ecf6  <=  wire_qout_00006_00019[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I20556d23c873c71c7ebc8a961bf40251     <=
                                             wire_qout_00006_00020[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00020 + 1 :
                                             wire_qout_00006_00020
                                             ;

            I68b152a599887c0039dd9d45c528c219  <=  wire_qout_00006_00020[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I79012e6351e6320c22437aa216ea4df1     <=
                                             wire_qout_00006_00021[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00021 + 1 :
                                             wire_qout_00006_00021
                                             ;

            Id051f1d5454802e0eb37e22248efe8ca  <=  wire_qout_00006_00021[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibf74ab9af877d27c3a6f3881f00ddaf1     <=
                                             wire_qout_00006_00022[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00006_00022 + 1 :
                                             wire_qout_00006_00022
                                             ;

            Ic4c6f707f461cebbc4c93f2ba664ae7b  <=  wire_qout_00006_00022[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I843d35db35d7b42a87ce78d3772cec2f     <=
                                             wire_qout_00007_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00000 + 1 :
                                             wire_qout_00007_00000
                                             ;

            Ia538dadbd6ae3711740595a18c89b65d  <=  wire_qout_00007_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2b1398b4bfd374d7221b0a68da28e979     <=
                                             wire_qout_00007_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00001 + 1 :
                                             wire_qout_00007_00001
                                             ;

            Ie7d9730b191781c78391141d95d4f8bd  <=  wire_qout_00007_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6f615d6e74b0c02f8e4265523ad16404     <=
                                             wire_qout_00007_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00002 + 1 :
                                             wire_qout_00007_00002
                                             ;

            I12f2f886517647044cc251861721bbb9  <=  wire_qout_00007_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iae8a98dd4a7cbfbc56c1404b6a2020af     <=
                                             wire_qout_00007_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00003 + 1 :
                                             wire_qout_00007_00003
                                             ;

            I615053b36a1851a06125e2ed5ec7f880  <=  wire_qout_00007_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iad53375a54d01c559c74981bf279dfb5     <=
                                             wire_qout_00007_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00004 + 1 :
                                             wire_qout_00007_00004
                                             ;

            Ifbc6aa14cd448bbe416897a3671ba857  <=  wire_qout_00007_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5db1307f922e0c742d7d9f3a79a4a4f3     <=
                                             wire_qout_00007_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00005 + 1 :
                                             wire_qout_00007_00005
                                             ;

            Ie596289582a73e37f78f4ca4cab21e3c  <=  wire_qout_00007_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9f78172ed5bf73752196f9a8810005f3     <=
                                             wire_qout_00007_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00006 + 1 :
                                             wire_qout_00007_00006
                                             ;

            Ifad8c7bacf72583f91be27fbe5b7a1e1  <=  wire_qout_00007_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If85a22d670d47f491dd7568d0453ba1d     <=
                                             wire_qout_00007_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00007 + 1 :
                                             wire_qout_00007_00007
                                             ;

            Ie74c72742807ae4243748fd27d80d626  <=  wire_qout_00007_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib9e529170b2896e930a839295796fd31     <=
                                             wire_qout_00007_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00008 + 1 :
                                             wire_qout_00007_00008
                                             ;

            Ie7a68c2b368a295f95571bc4a109b9f1  <=  wire_qout_00007_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib7af536846bac40c1f221d1f72c6c25c     <=
                                             wire_qout_00007_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00009 + 1 :
                                             wire_qout_00007_00009
                                             ;

            Id88a7edf897eea1b4a137141789a04f5  <=  wire_qout_00007_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib0eb61a2cb831dd35ce9850994e7c2da     <=
                                             wire_qout_00007_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00010 + 1 :
                                             wire_qout_00007_00010
                                             ;

            Ib13436ad16a37d656d6b1ee95b9aee20  <=  wire_qout_00007_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I89d338f59960af7a47595d6afa206abc     <=
                                             wire_qout_00007_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00011 + 1 :
                                             wire_qout_00007_00011
                                             ;

            Idc07dc30c0a957e474546ac7a60df38f  <=  wire_qout_00007_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib3c1176eb8991e3e85855a9fe845c303     <=
                                             wire_qout_00007_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00012 + 1 :
                                             wire_qout_00007_00012
                                             ;

            I595665d8128bb87ab62741d7ac520a4b  <=  wire_qout_00007_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I93073d05d509b821a743998cf32c58ee     <=
                                             wire_qout_00007_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00013 + 1 :
                                             wire_qout_00007_00013
                                             ;

            I256050251d23250854ff337bef28e460  <=  wire_qout_00007_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iab6dac1909c1564c3890ffecc13418df     <=
                                             wire_qout_00007_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00014 + 1 :
                                             wire_qout_00007_00014
                                             ;

            I82f0e5a32d1bcd761a74f1f9ce8c88ba  <=  wire_qout_00007_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1b75eeb29167a171d89f6e67039436d5     <=
                                             wire_qout_00007_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00015 + 1 :
                                             wire_qout_00007_00015
                                             ;

            I98febac90cccb5fc1f3d966b6e38c4d3  <=  wire_qout_00007_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3a31adc52a1405555017b2ddf219b407     <=
                                             wire_qout_00007_00016[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00016 + 1 :
                                             wire_qout_00007_00016
                                             ;

            Ib534288c2cf976b6ec85db743bc2a823  <=  wire_qout_00007_00016[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iaadba89c6a370240fc0758029f7d8db0     <=
                                             wire_qout_00007_00017[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00017 + 1 :
                                             wire_qout_00007_00017
                                             ;

            If988b82b86db1f4ff6d3695f7b0197e4  <=  wire_qout_00007_00017[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4f4a64fb3ced7d9f7ee4513178e9655a     <=
                                             wire_qout_00007_00018[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00018 + 1 :
                                             wire_qout_00007_00018
                                             ;

            I6ef260ef75e47b011a46ba2080ac3684  <=  wire_qout_00007_00018[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0c76ca58f69c91758e755cd581241284     <=
                                             wire_qout_00007_00019[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00019 + 1 :
                                             wire_qout_00007_00019
                                             ;

            Ifc1da524e7670772834d521a6fc4c96f  <=  wire_qout_00007_00019[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2312bce18958346149c868846e04643b     <=
                                             wire_qout_00007_00020[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00020 + 1 :
                                             wire_qout_00007_00020
                                             ;

            I852d5295a32984af00c95f6d9389555e  <=  wire_qout_00007_00020[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3e154098cb0a48f1c23234f46613f406     <=
                                             wire_qout_00007_00021[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00021 + 1 :
                                             wire_qout_00007_00021
                                             ;

            I3c0a621dbef864fd1f566bc2e47f32c6  <=  wire_qout_00007_00021[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1645c1c588bcbf15dd62d47e08b8e139     <=
                                             wire_qout_00007_00022[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00007_00022 + 1 :
                                             wire_qout_00007_00022
                                             ;

            Ic04828ba2db8239b093043c27476d345  <=  wire_qout_00007_00022[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4c25de66590e1745d37112e08d8c8e2c     <=
                                             wire_qout_00008_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00008_00000 + 1 :
                                             wire_qout_00008_00000
                                             ;

            I319012bc6fe93d78de57bcace0caaef5  <=  wire_qout_00008_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia03092ac621b8dd1c206fea1e8b0215f     <=
                                             wire_qout_00008_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00008_00001 + 1 :
                                             wire_qout_00008_00001
                                             ;

            Ibb35bace971548c9fc98d773d1aff712  <=  wire_qout_00008_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5c9bdb033436dc9f6069baca31f24c2d     <=
                                             wire_qout_00008_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00008_00002 + 1 :
                                             wire_qout_00008_00002
                                             ;

            I90023493600924a76d2192080cf6194e  <=  wire_qout_00008_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8f07cf4865480f18ad6945974ec2231c     <=
                                             wire_qout_00008_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00008_00003 + 1 :
                                             wire_qout_00008_00003
                                             ;

            Ia9f5ce4603af279bbd9b486b67016482  <=  wire_qout_00008_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4a7119e8862fe4a6a4100dd9ac67dd24     <=
                                             wire_qout_00008_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00008_00004 + 1 :
                                             wire_qout_00008_00004
                                             ;

            I05721e06a1acdcc0571907c7d853f18c  <=  wire_qout_00008_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id78fcfc6724a05f46d44d7c3e7d0c756     <=
                                             wire_qout_00008_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00008_00005 + 1 :
                                             wire_qout_00008_00005
                                             ;

            Ibfcfd3151af0d82bfce293ada44059b3  <=  wire_qout_00008_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7cbd9d619623cbabf8ed6b1fece8f012     <=
                                             wire_qout_00008_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00008_00006 + 1 :
                                             wire_qout_00008_00006
                                             ;

            I9539fcc40d26b13015a864718b116d5b  <=  wire_qout_00008_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I58951165d251e370b0f3b3fb537aed18     <=
                                             wire_qout_00008_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00008_00007 + 1 :
                                             wire_qout_00008_00007
                                             ;

            I5490039998187a1a2efc3549e3dee7d6  <=  wire_qout_00008_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I21daac106f526d84cb8fa5239c19499d     <=
                                             wire_qout_00008_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00008_00008 + 1 :
                                             wire_qout_00008_00008
                                             ;

            I2b97a79c90f6578c8b2f321f8d598cc8  <=  wire_qout_00008_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I178029cec3a5d6141abdfa91b91fdbf4     <=
                                             wire_qout_00008_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00008_00009 + 1 :
                                             wire_qout_00008_00009
                                             ;

            I0c616f736879c28a5222de3d6f49a587  <=  wire_qout_00008_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I96dfb2efbb55a644616e3474ed07c364     <=
                                             wire_qout_00009_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00009_00000 + 1 :
                                             wire_qout_00009_00000
                                             ;

            I5590d801fd7fb496019d4c31b7c6d898  <=  wire_qout_00009_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7a17d8f0e2d16c441044db68ee037731     <=
                                             wire_qout_00009_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00009_00001 + 1 :
                                             wire_qout_00009_00001
                                             ;

            I27e1d2e0e980216b27b90ea48c061025  <=  wire_qout_00009_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2ced9bb3ae6bdc5b5ef2865fb46abf07     <=
                                             wire_qout_00009_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00009_00002 + 1 :
                                             wire_qout_00009_00002
                                             ;

            I474f6bd977f4197742d0bddb3bece684  <=  wire_qout_00009_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I89a93384020d93cf4d26b3902e06cd9e     <=
                                             wire_qout_00009_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00009_00003 + 1 :
                                             wire_qout_00009_00003
                                             ;

            Iaa1e981134f5a5c02983c49562683bc5  <=  wire_qout_00009_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibbb47d29b9a45559c13ffa3b046c66f5     <=
                                             wire_qout_00009_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00009_00004 + 1 :
                                             wire_qout_00009_00004
                                             ;

            Ib051eb1091a85f85a1e50007f1b27cab  <=  wire_qout_00009_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0034177eb1049577a3578b371527f34b     <=
                                             wire_qout_00009_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00009_00005 + 1 :
                                             wire_qout_00009_00005
                                             ;

            I6b5645cdde4b35a16fe3e91d90caaa4e  <=  wire_qout_00009_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I22d9ea7bb5a1a3405bcd04b9af40fa62     <=
                                             wire_qout_00009_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00009_00006 + 1 :
                                             wire_qout_00009_00006
                                             ;

            I8850ab26807dcd55fefadf6310729ca7  <=  wire_qout_00009_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8a632e7a911bf5726fee587189cb6f16     <=
                                             wire_qout_00009_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00009_00007 + 1 :
                                             wire_qout_00009_00007
                                             ;

            Ic5cb81c821716a8aabf8cc2283ff73ba  <=  wire_qout_00009_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3765afc490b34e8a310998a4ebcff8cb     <=
                                             wire_qout_00009_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00009_00008 + 1 :
                                             wire_qout_00009_00008
                                             ;

            I9a6923c6368526a53ef70e16471386ef  <=  wire_qout_00009_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7607e800ae46a96e016b303120da4247     <=
                                             wire_qout_00009_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00009_00009 + 1 :
                                             wire_qout_00009_00009
                                             ;

            I620b8ecdcaccc1ec80ebcf9fa6af0017  <=  wire_qout_00009_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I29b2f1fddee5e32f217d25410bcfce4f     <=
                                             wire_qout_00010_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00010_00000 + 1 :
                                             wire_qout_00010_00000
                                             ;

            I141cda06bae0c5666e3bc61c6fe5ad66  <=  wire_qout_00010_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iba5f8a31a81f6aa06f5e38c03dc6db54     <=
                                             wire_qout_00010_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00010_00001 + 1 :
                                             wire_qout_00010_00001
                                             ;

            Ia9c273b32d0701c7f185ab2de9e57829  <=  wire_qout_00010_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifcb5c907ad503331317599e4e0ce7be8     <=
                                             wire_qout_00010_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00010_00002 + 1 :
                                             wire_qout_00010_00002
                                             ;

            Ic3fb524ab434e80b3289c9241b65d224  <=  wire_qout_00010_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I62d6f2ab4ec8b6ecfa544ad4d90eb30b     <=
                                             wire_qout_00010_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00010_00003 + 1 :
                                             wire_qout_00010_00003
                                             ;

            I23c8b64e433af0bd00cef44e38df99f8  <=  wire_qout_00010_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ide65414c51b3cb182c0f2f238903d60a     <=
                                             wire_qout_00010_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00010_00004 + 1 :
                                             wire_qout_00010_00004
                                             ;

            If6a5dc79c0f6ce348956286737a369d8  <=  wire_qout_00010_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I03a8dc2288eaeb619e746990e20cc868     <=
                                             wire_qout_00010_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00010_00005 + 1 :
                                             wire_qout_00010_00005
                                             ;

            I34e6e9d2153e4a70ee36ab85e72d5318  <=  wire_qout_00010_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id81c1b44d16ddbcd466382c60fe84986     <=
                                             wire_qout_00010_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00010_00006 + 1 :
                                             wire_qout_00010_00006
                                             ;

            Ifdabf743a8cb46b7053000ff48ea0c60  <=  wire_qout_00010_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I503d72f4a2fd20dbf35aa27321d2ede7     <=
                                             wire_qout_00010_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00010_00007 + 1 :
                                             wire_qout_00010_00007
                                             ;

            I22f5bb821a2571d1764978fd76c8f1d0  <=  wire_qout_00010_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id6595a4cf33062d1f05cbcee2d0685f1     <=
                                             wire_qout_00010_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00010_00008 + 1 :
                                             wire_qout_00010_00008
                                             ;

            I1b695aa715615662eff7065c742b0859  <=  wire_qout_00010_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I83ebdd7331ca8fbcf5250851b346c0b0     <=
                                             wire_qout_00010_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00010_00009 + 1 :
                                             wire_qout_00010_00009
                                             ;

            Iec91b3ca3b54010755d57f8b8ea4a544  <=  wire_qout_00010_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7f6ea26cdfe5986065e7b5aa6842cc1c     <=
                                             wire_qout_00011_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00011_00000 + 1 :
                                             wire_qout_00011_00000
                                             ;

            I06ad520cb02e46d34c45f207d42a9243  <=  wire_qout_00011_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idab1ec32c20f93c4cc1acb38158f92d5     <=
                                             wire_qout_00011_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00011_00001 + 1 :
                                             wire_qout_00011_00001
                                             ;

            I9d18ff3465afd8cae63abba68487542e  <=  wire_qout_00011_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0738add83419502e73674ded2f1ad6c7     <=
                                             wire_qout_00011_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00011_00002 + 1 :
                                             wire_qout_00011_00002
                                             ;

            I914dedc1d5e5e21c9b8d07ec0ecc01f9  <=  wire_qout_00011_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6c93e63a8e5a2dbd598f1565c7323b39     <=
                                             wire_qout_00011_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00011_00003 + 1 :
                                             wire_qout_00011_00003
                                             ;

            I3375fff5ee0d4b4b12c5a70fbdee59fe  <=  wire_qout_00011_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4aa57a9d46371f1680d5f95596f60b5d     <=
                                             wire_qout_00011_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00011_00004 + 1 :
                                             wire_qout_00011_00004
                                             ;

            Ia8e304ca12c82e41cb8e4de7be199394  <=  wire_qout_00011_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5369a7203b78951a3c006c2d3b22507c     <=
                                             wire_qout_00011_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00011_00005 + 1 :
                                             wire_qout_00011_00005
                                             ;

            I3566f2779e860008b1a5d305366a07c9  <=  wire_qout_00011_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie72a79a6966cf198687b7c8a8bcdeb13     <=
                                             wire_qout_00011_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00011_00006 + 1 :
                                             wire_qout_00011_00006
                                             ;

            Ie68b31360c12a83c6095254b6f14603c  <=  wire_qout_00011_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie917ae4c44ab0f9c2f1747ff0d2a754e     <=
                                             wire_qout_00011_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00011_00007 + 1 :
                                             wire_qout_00011_00007
                                             ;

            I42ae0c42360c977b35429ce290516a6f  <=  wire_qout_00011_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0b1a31ccb34a742552c11b1945e23dd8     <=
                                             wire_qout_00011_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00011_00008 + 1 :
                                             wire_qout_00011_00008
                                             ;

            Ibe01835305315fab50269c72ef849b61  <=  wire_qout_00011_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9a65a845cf2eced39050e8481665f557     <=
                                             wire_qout_00011_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00011_00009 + 1 :
                                             wire_qout_00011_00009
                                             ;

            Id806a2df1c4519bbbe811791cb4072f9  <=  wire_qout_00011_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3b402b35d38a9fde312c89b82297c1a5     <=
                                             wire_qout_00012_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00012_00000 + 1 :
                                             wire_qout_00012_00000
                                             ;

            Ifb70a30f8bade95f402e71f95fe6644b  <=  wire_qout_00012_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I309fa33562370e339c19e2377e6a6a7a     <=
                                             wire_qout_00012_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00012_00001 + 1 :
                                             wire_qout_00012_00001
                                             ;

            I592a495aecc800236c3470ff8e6adbb5  <=  wire_qout_00012_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7d06aed81222a030837cad2074c68e19     <=
                                             wire_qout_00012_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00012_00002 + 1 :
                                             wire_qout_00012_00002
                                             ;

            I1c8024aa9d81704d2dcf63e34853f8cf  <=  wire_qout_00012_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I835cc6af0cd8189035f2441c2e0d3100     <=
                                             wire_qout_00012_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00012_00003 + 1 :
                                             wire_qout_00012_00003
                                             ;

            Ief03713f5cf37200373a20d42c7fc9eb  <=  wire_qout_00012_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If6f768d12f04087246a0d65de1aef99b     <=
                                             wire_qout_00012_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00012_00004 + 1 :
                                             wire_qout_00012_00004
                                             ;

            Ic3cb34aae74c5f1a870b3635f8a40764  <=  wire_qout_00012_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie4b180e1e2cadb865b0eaf6509f99dbb     <=
                                             wire_qout_00013_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00013_00000 + 1 :
                                             wire_qout_00013_00000
                                             ;

            Ifa3df8b249467cc1e827c69925ef415f  <=  wire_qout_00013_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie329a11fc3f6f59f6f1790612fde3250     <=
                                             wire_qout_00013_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00013_00001 + 1 :
                                             wire_qout_00013_00001
                                             ;

            Icf3ad912aaeaa0c5cd1ab0edb898d6e8  <=  wire_qout_00013_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idb7ddbee4076f7bf49177e69f5e4d112     <=
                                             wire_qout_00013_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00013_00002 + 1 :
                                             wire_qout_00013_00002
                                             ;

            Ib774f380e3d7cfd1f5f064e93d8134b4  <=  wire_qout_00013_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I614d66a7dca2d08efdfdc157ca803d5c     <=
                                             wire_qout_00013_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00013_00003 + 1 :
                                             wire_qout_00013_00003
                                             ;

            Ic07c650e6e49892a41cfaf3a37471426  <=  wire_qout_00013_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iea16eb0ab70ebb1bc47ae55e11ced62d     <=
                                             wire_qout_00013_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00013_00004 + 1 :
                                             wire_qout_00013_00004
                                             ;

            Ib1073489d63ea33d7f3892f4ff875358  <=  wire_qout_00013_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifa8db43284d5bbebaed4f72d65cf9f92     <=
                                             wire_qout_00014_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00014_00000 + 1 :
                                             wire_qout_00014_00000
                                             ;

            I174b6c36f2af82f8047cc76543a3b4ee  <=  wire_qout_00014_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I365d9f3e8b2a9890427f07386deeb093     <=
                                             wire_qout_00014_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00014_00001 + 1 :
                                             wire_qout_00014_00001
                                             ;

            I953b975a89adcc88039284970e9b3404  <=  wire_qout_00014_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I466aaa0b6cde2ade1901797b8c11e32c     <=
                                             wire_qout_00014_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00014_00002 + 1 :
                                             wire_qout_00014_00002
                                             ;

            If2b40d249c531e10cc22d1335f350441  <=  wire_qout_00014_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7057e329a65ab240ed6cfa824307af65     <=
                                             wire_qout_00014_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00014_00003 + 1 :
                                             wire_qout_00014_00003
                                             ;

            I44ccc3ae897109dd51f9afeef93daca4  <=  wire_qout_00014_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I624e50e3457d33d12680eaf8e7c34aa3     <=
                                             wire_qout_00014_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00014_00004 + 1 :
                                             wire_qout_00014_00004
                                             ;

            Ie9236599cea94cfb603c6b977fdbb44a  <=  wire_qout_00014_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9f356fd6820c33fdb5baff05a781e192     <=
                                             wire_qout_00015_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00015_00000 + 1 :
                                             wire_qout_00015_00000
                                             ;

            I25f1ee9cee4d04bd8fec1fe601d016d7  <=  wire_qout_00015_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I39b9c7c664fe7017731877d145d55b44     <=
                                             wire_qout_00015_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00015_00001 + 1 :
                                             wire_qout_00015_00001
                                             ;

            I5ec1e530b9007a75a778af4d82ab427b  <=  wire_qout_00015_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic62ffbb9e58e0d08b0dec24bba1dc6f2     <=
                                             wire_qout_00015_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00015_00002 + 1 :
                                             wire_qout_00015_00002
                                             ;

            I8a9e516aa824260998d10db758642bb0  <=  wire_qout_00015_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8da2a532288fb817e7dc0cb7b4e3761c     <=
                                             wire_qout_00015_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00015_00003 + 1 :
                                             wire_qout_00015_00003
                                             ;

            I70dd1350d65155ee7b562f4c79024a3d  <=  wire_qout_00015_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6a6e559f5c98f846014e8107fea5a5d9     <=
                                             wire_qout_00015_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00015_00004 + 1 :
                                             wire_qout_00015_00004
                                             ;

            Ic9146d8b3dd0c612073b70b8a8791e8c  <=  wire_qout_00015_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibef9219f577b1a62dfdd77296fbfb24d     <=
                                             wire_qout_00016_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00016_00000 + 1 :
                                             wire_qout_00016_00000
                                             ;

            I857d3155df0b6dd704514b039c66fa97  <=  wire_qout_00016_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I52e6688b5bfff75529d18e20b22832ce     <=
                                             wire_qout_00016_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00016_00001 + 1 :
                                             wire_qout_00016_00001
                                             ;

            Idc1b8aa2f81a7fbd87e4f5821d14bf01  <=  wire_qout_00016_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iff22c49354eefca0ea3c5959c14b782c     <=
                                             wire_qout_00016_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00016_00002 + 1 :
                                             wire_qout_00016_00002
                                             ;

            I68b585571699a57bc6ba5e8955467119  <=  wire_qout_00016_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie5377bbdb4111ed00356d5b7737102f3     <=
                                             wire_qout_00016_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00016_00003 + 1 :
                                             wire_qout_00016_00003
                                             ;

            Ib70e99c3acc76286a6811bcacc9284de  <=  wire_qout_00016_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I55bf0f3379a8c44634b8f0a3d06c049e     <=
                                             wire_qout_00016_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00016_00004 + 1 :
                                             wire_qout_00016_00004
                                             ;

            Iee17ece482d04964d3c21a092ec955a4  <=  wire_qout_00016_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9bc9541607f4f6aedb686cdde297bcda     <=
                                             wire_qout_00017_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00017_00000 + 1 :
                                             wire_qout_00017_00000
                                             ;

            I5a247475beb737d470f03507e55f5b24  <=  wire_qout_00017_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia4620554fbb1d81a71a15a846e4be2f5     <=
                                             wire_qout_00017_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00017_00001 + 1 :
                                             wire_qout_00017_00001
                                             ;

            I13b0c9578f7b6b3b7e6704d7b44079c4  <=  wire_qout_00017_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibb31b35388ba8ba2ecf98449308ee67d     <=
                                             wire_qout_00017_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00017_00002 + 1 :
                                             wire_qout_00017_00002
                                             ;

            I41eff06fe1dea8be4613945de596d3ca  <=  wire_qout_00017_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia20410fb3d56587f89a54c00b943b305     <=
                                             wire_qout_00017_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00017_00003 + 1 :
                                             wire_qout_00017_00003
                                             ;

            I08f22261d5713c0636d77c7938f592d6  <=  wire_qout_00017_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9d268f3da12e35b9a4229b7340c0f018     <=
                                             wire_qout_00017_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00017_00004 + 1 :
                                             wire_qout_00017_00004
                                             ;

            I1c7e41b9cb1bdb6f649c88c0ed3f4100  <=  wire_qout_00017_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2fce29bd666082eedb2fb3ec8b5ae4dd     <=
                                             wire_qout_00018_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00018_00000 + 1 :
                                             wire_qout_00018_00000
                                             ;

            Idd59a5357d4c835379ed180ac0924bf1  <=  wire_qout_00018_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia1e8b61e2579a90f5c88ded11c7322c2     <=
                                             wire_qout_00018_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00018_00001 + 1 :
                                             wire_qout_00018_00001
                                             ;

            Ibe7e5c2cb9c50eca34a3859d13e83a92  <=  wire_qout_00018_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8cf3718ba65b7fed72e3955f190e34d1     <=
                                             wire_qout_00018_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00018_00002 + 1 :
                                             wire_qout_00018_00002
                                             ;

            Ibf5c141c5cc0a6a20c05b52bf8282476  <=  wire_qout_00018_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7e802d300af54d394b4ee041798c0513     <=
                                             wire_qout_00018_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00018_00003 + 1 :
                                             wire_qout_00018_00003
                                             ;

            I0038305f94aaefe2cd1a243580d95932  <=  wire_qout_00018_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id4fd5a4b97cfa1e176a26f3a823c5516     <=
                                             wire_qout_00018_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00018_00004 + 1 :
                                             wire_qout_00018_00004
                                             ;

            I5364deb983adc2ae505ed2b8c57f876d  <=  wire_qout_00018_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icbf8d4e75fc66c05eb49c5075696fb07     <=
                                             wire_qout_00019_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00019_00000 + 1 :
                                             wire_qout_00019_00000
                                             ;

            Ifdb5589982db805a0416e1c01276249a  <=  wire_qout_00019_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I746a7e90adb2f213b75ae12a161aca0d     <=
                                             wire_qout_00019_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00019_00001 + 1 :
                                             wire_qout_00019_00001
                                             ;

            I8bb5522183b65583fda83067990b3e94  <=  wire_qout_00019_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icb1029aaaaed8c698862ea9c5e22132c     <=
                                             wire_qout_00019_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00019_00002 + 1 :
                                             wire_qout_00019_00002
                                             ;

            I1e77fe6aeaba852aba34ed37dd53add6  <=  wire_qout_00019_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib93ea7028c172373b53cdafecae32a67     <=
                                             wire_qout_00019_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00019_00003 + 1 :
                                             wire_qout_00019_00003
                                             ;

            I9171019227f35760d02d0c8ce786f4d3  <=  wire_qout_00019_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If9628275b000e418f3903daebfdace92     <=
                                             wire_qout_00019_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00019_00004 + 1 :
                                             wire_qout_00019_00004
                                             ;

            I6e92a48aaab94074a555efa9bd1e7243  <=  wire_qout_00019_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I830202fb6f08f98c7f71893a881bd555     <=
                                             wire_qout_00020_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00000 + 1 :
                                             wire_qout_00020_00000
                                             ;

            I3bc094d67805664859fdcb66f1360e64  <=  wire_qout_00020_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6f38bc9359562f57c1603355e9ee312b     <=
                                             wire_qout_00020_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00001 + 1 :
                                             wire_qout_00020_00001
                                             ;

            I2518ccf385b3b677d95983bc550282e8  <=  wire_qout_00020_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4701b732d59c26e3790a63c1936f9a24     <=
                                             wire_qout_00020_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00002 + 1 :
                                             wire_qout_00020_00002
                                             ;

            I7547c56b32513ad45d775b4502596d9d  <=  wire_qout_00020_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib5d28d8f73d17ab6df6a1291e50c04ab     <=
                                             wire_qout_00020_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00003 + 1 :
                                             wire_qout_00020_00003
                                             ;

            I013d84bfd582acc7accf07ec522961fa  <=  wire_qout_00020_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I81259f391db792339824ad5dd1a0057b     <=
                                             wire_qout_00020_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00004 + 1 :
                                             wire_qout_00020_00004
                                             ;

            I0ec27b590ee6dcdd9c1086105e3b6c23  <=  wire_qout_00020_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6f09ac63effe67a86798b9b4e1690664     <=
                                             wire_qout_00020_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00005 + 1 :
                                             wire_qout_00020_00005
                                             ;

            I4cdc955fa9afc75c2c977de4ec540e1e  <=  wire_qout_00020_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I370b4b3a0048a93ba374a40e170c75a3     <=
                                             wire_qout_00020_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00006 + 1 :
                                             wire_qout_00020_00006
                                             ;

            Ieefbb5d6f4ac1e586832c5c0f513c5a2  <=  wire_qout_00020_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3f8476d0aa0ea2439b67ea1a4adf36c5     <=
                                             wire_qout_00020_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00007 + 1 :
                                             wire_qout_00020_00007
                                             ;

            Ic828cdd5dfde844df4c150921af2a443  <=  wire_qout_00020_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I35b52dba10a8a5b22b518388fecac82d     <=
                                             wire_qout_00020_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00008 + 1 :
                                             wire_qout_00020_00008
                                             ;

            Idf1ecab26889c4adcb835fda6b1cb368  <=  wire_qout_00020_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic7db274ed18e6fdecf30381a31238777     <=
                                             wire_qout_00020_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00009 + 1 :
                                             wire_qout_00020_00009
                                             ;

            I00d3f14b20e1ea7d726533386e0eba27  <=  wire_qout_00020_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2c4e538a8db759e9799541d9178ec61e     <=
                                             wire_qout_00020_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00010 + 1 :
                                             wire_qout_00020_00010
                                             ;

            I7f720a18542528f0c9bfb14f699ff4da  <=  wire_qout_00020_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ief6d4c3f5ef8663e111ef99347b023f5     <=
                                             wire_qout_00020_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00011 + 1 :
                                             wire_qout_00020_00011
                                             ;

            Ia98a6f01e4eb5bc74d50d350e79be426  <=  wire_qout_00020_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id95e964e5faecb52c72669b0d28a4bf5     <=
                                             wire_qout_00020_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00012 + 1 :
                                             wire_qout_00020_00012
                                             ;

            I182b43872d50de6f7afb700f178b160e  <=  wire_qout_00020_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0fcef4538102ac6d24aa7090d5405afa     <=
                                             wire_qout_00020_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00020_00013 + 1 :
                                             wire_qout_00020_00013
                                             ;

            Ic9b72b2a91d951cf08cf54ed215ecaa8  <=  wire_qout_00020_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I055019e38eec6badd1739033d43d7d97     <=
                                             wire_qout_00021_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00000 + 1 :
                                             wire_qout_00021_00000
                                             ;

            I93084ccf5b5e4efaee968b497bb2a775  <=  wire_qout_00021_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I35c20a6e823da77a870b421eef2e0a95     <=
                                             wire_qout_00021_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00001 + 1 :
                                             wire_qout_00021_00001
                                             ;

            Id38852415486e6989b89a0d85ad6771b  <=  wire_qout_00021_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I32cc12cdacef1a4ef64577e0fa977f46     <=
                                             wire_qout_00021_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00002 + 1 :
                                             wire_qout_00021_00002
                                             ;

            I17cf58ef5326978c62c03c56090a299f  <=  wire_qout_00021_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I26b3f2360ca4a8caee61b2f3a3a08267     <=
                                             wire_qout_00021_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00003 + 1 :
                                             wire_qout_00021_00003
                                             ;

            Ie41ca18c7d11a47e274f9c33f75393ec  <=  wire_qout_00021_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5ef9b7dc0c63e9ca6a5fb5f7ffa06041     <=
                                             wire_qout_00021_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00004 + 1 :
                                             wire_qout_00021_00004
                                             ;

            I7b80b4902fe98c10dd72c9eb082346e5  <=  wire_qout_00021_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If881473b05090f40a027d7eeee7f7ed9     <=
                                             wire_qout_00021_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00005 + 1 :
                                             wire_qout_00021_00005
                                             ;

            I20ffba20af04b99954bf719589e90d1a  <=  wire_qout_00021_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I23bd59ab5b038935301396aaf2acefc1     <=
                                             wire_qout_00021_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00006 + 1 :
                                             wire_qout_00021_00006
                                             ;

            If8fe5af7e5c3c97b5a713f6bcf919f1f  <=  wire_qout_00021_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I874386d94dacf84e699d159af1a49836     <=
                                             wire_qout_00021_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00007 + 1 :
                                             wire_qout_00021_00007
                                             ;

            Idc5fb0f3a04ab32948e249e088a11b11  <=  wire_qout_00021_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I95bfe51a759bf4165168e5e3b99d6b34     <=
                                             wire_qout_00021_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00008 + 1 :
                                             wire_qout_00021_00008
                                             ;

            Ia9f1e580e8f441394d719d52a7bad688  <=  wire_qout_00021_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4ba5b2f9b7ec0937ecd2c9945cf6de87     <=
                                             wire_qout_00021_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00009 + 1 :
                                             wire_qout_00021_00009
                                             ;

            I02849282dd1bd663fd39baccf41762f9  <=  wire_qout_00021_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0b08fb8db0e8a1de3d416907c87fe700     <=
                                             wire_qout_00021_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00010 + 1 :
                                             wire_qout_00021_00010
                                             ;

            Ie4cda4648f6ceb76b8fb74f290ab6439  <=  wire_qout_00021_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie030d12e5acf9ef4975a17c83b2481c1     <=
                                             wire_qout_00021_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00011 + 1 :
                                             wire_qout_00021_00011
                                             ;

            I24135210c23b2422a42c90ee25594191  <=  wire_qout_00021_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia7a0e852d3dfcef950804ea0ebb0c80a     <=
                                             wire_qout_00021_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00012 + 1 :
                                             wire_qout_00021_00012
                                             ;

            Ib08897f9216599042f7b97b137e07fe1  <=  wire_qout_00021_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iaa4c38d030eab2b7899399aa0d7886d9     <=
                                             wire_qout_00021_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00021_00013 + 1 :
                                             wire_qout_00021_00013
                                             ;

            I51e14ece9ab6607f83e6ba27f3f046a9  <=  wire_qout_00021_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icce7ff1d652d4d9c2be5ecf679059bbe     <=
                                             wire_qout_00022_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00000 + 1 :
                                             wire_qout_00022_00000
                                             ;

            I7a626ec321bf963a5401892a7e3891c7  <=  wire_qout_00022_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If816bc5eacaea23443602e575ddf60b8     <=
                                             wire_qout_00022_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00001 + 1 :
                                             wire_qout_00022_00001
                                             ;

            If76f04fe0baf171d7df2c0cd849aea2b  <=  wire_qout_00022_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3b224a4ded05446cc5300d430bdd1947     <=
                                             wire_qout_00022_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00002 + 1 :
                                             wire_qout_00022_00002
                                             ;

            Ia9c8cc5e3becf3d48feedec8fa2c93a4  <=  wire_qout_00022_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia5fc5cfb0e52237b407b37a3858fccb5     <=
                                             wire_qout_00022_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00003 + 1 :
                                             wire_qout_00022_00003
                                             ;

            If3b77c41fabcdb283f2c6fdacaa5e9a4  <=  wire_qout_00022_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I92f8ba6e7f8e9b30fb5b6973eb8fd03e     <=
                                             wire_qout_00022_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00004 + 1 :
                                             wire_qout_00022_00004
                                             ;

            Ie5373b01a92f2ff85be8077cfef2175a  <=  wire_qout_00022_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icdfa60d2a024dd934f7e6639c6cb2c28     <=
                                             wire_qout_00022_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00005 + 1 :
                                             wire_qout_00022_00005
                                             ;

            I5109afc4dc91780e05704ea5e1399e3e  <=  wire_qout_00022_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifff70b976513eaa42b6bd4b80c98611e     <=
                                             wire_qout_00022_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00006 + 1 :
                                             wire_qout_00022_00006
                                             ;

            I3e0b41bee4c76eb5f3340ad23bfa01ad  <=  wire_qout_00022_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ica12fa8b631b70a6bbe9f6e92bf73ea0     <=
                                             wire_qout_00022_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00007 + 1 :
                                             wire_qout_00022_00007
                                             ;

            Ic0732810fd355d59a3168be896a0f9ac  <=  wire_qout_00022_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie69c255335760f706c644b115887269b     <=
                                             wire_qout_00022_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00008 + 1 :
                                             wire_qout_00022_00008
                                             ;

            I220e32641265b46527ca61111f7ebf1b  <=  wire_qout_00022_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idb06676b41de19bc86eae34c292183d9     <=
                                             wire_qout_00022_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00009 + 1 :
                                             wire_qout_00022_00009
                                             ;

            Ice59d2af73d0b0f2ae91a2ef0c2b7f04  <=  wire_qout_00022_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib21d2306d5ded3406fac754e69a10d20     <=
                                             wire_qout_00022_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00010 + 1 :
                                             wire_qout_00022_00010
                                             ;

            Ic308610ea8bb62ecb6094192e02dbdba  <=  wire_qout_00022_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib41d1aa2dcf81879976fb8964cbf6f79     <=
                                             wire_qout_00022_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00011 + 1 :
                                             wire_qout_00022_00011
                                             ;

            I33ee415d85e2bcd8f975d34b880f6ea7  <=  wire_qout_00022_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5f8f5e246f008b8d8c75f72828337bab     <=
                                             wire_qout_00022_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00012 + 1 :
                                             wire_qout_00022_00012
                                             ;

            Ie61f299252b8fecfd3e8634b64df5a90  <=  wire_qout_00022_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id6625e78da0e14d2eeb19cc8ac6520e0     <=
                                             wire_qout_00022_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00022_00013 + 1 :
                                             wire_qout_00022_00013
                                             ;

            Icc67656ad2dd3fffae4e5abe02f8fff9  <=  wire_qout_00022_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6d9ddc6afa559ac35c042df1a9390ce9     <=
                                             wire_qout_00023_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00000 + 1 :
                                             wire_qout_00023_00000
                                             ;

            I0c47ccef4b55410286248884a7249703  <=  wire_qout_00023_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9334055c7833676469670372d3c5cc31     <=
                                             wire_qout_00023_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00001 + 1 :
                                             wire_qout_00023_00001
                                             ;

            I94e4041b482064334fd0ed92b91bde89  <=  wire_qout_00023_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0c97d772c737c6ff85b584bf69ccaf93     <=
                                             wire_qout_00023_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00002 + 1 :
                                             wire_qout_00023_00002
                                             ;

            I39d3bce4060032a81e6b6a1c1805cfe8  <=  wire_qout_00023_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic6ce97ae85d91dd8a79f3f9d0da375a2     <=
                                             wire_qout_00023_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00003 + 1 :
                                             wire_qout_00023_00003
                                             ;

            Ifb422c30663eb4824caa72326b238df6  <=  wire_qout_00023_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I83ff9a2750b298b0f7c9b6ce13f574af     <=
                                             wire_qout_00023_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00004 + 1 :
                                             wire_qout_00023_00004
                                             ;

            I41ab6fb6ec6ef7ffff70e50f25f217b6  <=  wire_qout_00023_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I85699a2a05c343a6a9e828af6d445e9e     <=
                                             wire_qout_00023_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00005 + 1 :
                                             wire_qout_00023_00005
                                             ;

            I3ce10718a2211184999663c3c2493cc1  <=  wire_qout_00023_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I51f6e39b24b2554884e381be79f47ff2     <=
                                             wire_qout_00023_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00006 + 1 :
                                             wire_qout_00023_00006
                                             ;

            I877e8d94236c3d8b0a31858a98fba5d6  <=  wire_qout_00023_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9f65fd05c6929300860c8cbbde5607f2     <=
                                             wire_qout_00023_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00007 + 1 :
                                             wire_qout_00023_00007
                                             ;

            Iff2f1716cbd73b406d8f07c22dc79fc8  <=  wire_qout_00023_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If09761d8f06051d4287ee29ac9c9fa19     <=
                                             wire_qout_00023_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00008 + 1 :
                                             wire_qout_00023_00008
                                             ;

            Ibc48fabc172f27ebce18d0a9b5120dc5  <=  wire_qout_00023_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I33bfbe0bcca6d32c86b9576577e3f265     <=
                                             wire_qout_00023_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00009 + 1 :
                                             wire_qout_00023_00009
                                             ;

            Ie562ebb336e476a81f20a652d4cb20f1  <=  wire_qout_00023_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If2921210b1c05ecbf00af3a2bcb96ef4     <=
                                             wire_qout_00023_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00010 + 1 :
                                             wire_qout_00023_00010
                                             ;

            Ib5ee5a6ffc45ed1fece0822dc4619b57  <=  wire_qout_00023_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib074e38e280474a782da831a3e0028b4     <=
                                             wire_qout_00023_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00011 + 1 :
                                             wire_qout_00023_00011
                                             ;

            I86ba73ee348f80e2f9891d2ebc8a02ed  <=  wire_qout_00023_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I507449dde0bc0c8f53a10759436ec731     <=
                                             wire_qout_00023_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00012 + 1 :
                                             wire_qout_00023_00012
                                             ;

            I1e96d5af3d0e3fdce39530dfd0131a7d  <=  wire_qout_00023_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id55a3e3f2d75baeba71a345fad695c69     <=
                                             wire_qout_00023_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00023_00013 + 1 :
                                             wire_qout_00023_00013
                                             ;

            I38352b363fa37f6f822fbc1a39100968  <=  wire_qout_00023_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I20984f43d22671639a7a178ad15aec04     <=
                                             wire_qout_00024_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00024_00000 + 1 :
                                             wire_qout_00024_00000
                                             ;

            I4ba41864bb1d2130c6971e0b2903027a  <=  wire_qout_00024_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I59f88336d6bdd50ded87d353fb5ce3e9     <=
                                             wire_qout_00024_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00024_00001 + 1 :
                                             wire_qout_00024_00001
                                             ;

            Ib68deeb7bec4ca3585d1a4dcbf8793f1  <=  wire_qout_00024_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I488635e3f7ed77ea88199f5bffd4b1d6     <=
                                             wire_qout_00024_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00024_00002 + 1 :
                                             wire_qout_00024_00002
                                             ;

            Ida3d808d100e0bba290f96ed9e744e65  <=  wire_qout_00024_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie6893017d21c050ba10d206854f4a9f4     <=
                                             wire_qout_00024_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00024_00003 + 1 :
                                             wire_qout_00024_00003
                                             ;

            I4d4901ff372f6820ca9c8c29cefa664a  <=  wire_qout_00024_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id3f68b4dc0ab60673208b7d2081f3533     <=
                                             wire_qout_00024_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00024_00004 + 1 :
                                             wire_qout_00024_00004
                                             ;

            Ib99e1b93fb7fbda260d93eea3d24c3e9  <=  wire_qout_00024_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I433756b944e061a824a89bda241e879f     <=
                                             wire_qout_00024_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00024_00005 + 1 :
                                             wire_qout_00024_00005
                                             ;

            I019e399a1cef87745e025a7d74e94db0  <=  wire_qout_00024_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2eb60a922aa4f7482dd92b9351d53a2d     <=
                                             wire_qout_00024_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00024_00006 + 1 :
                                             wire_qout_00024_00006
                                             ;

            Ia8974083bfd064f2c27dcd421490fcfd  <=  wire_qout_00024_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0867979e1b159c8ceae548930376f482     <=
                                             wire_qout_00025_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00025_00000 + 1 :
                                             wire_qout_00025_00000
                                             ;

            I8fd5787ebf758919e7cb75d7419441e8  <=  wire_qout_00025_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4accfbeae8a5ee0dbeab23ef3a116145     <=
                                             wire_qout_00025_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00025_00001 + 1 :
                                             wire_qout_00025_00001
                                             ;

            Id14074d5230885c38b89b09b130ecf68  <=  wire_qout_00025_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic7570b0b7c5bef5758f68562ae4c90f6     <=
                                             wire_qout_00025_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00025_00002 + 1 :
                                             wire_qout_00025_00002
                                             ;

            I86fefad34d3c864dd0e725133f303b4f  <=  wire_qout_00025_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iceadadc4456881fdeea85934a9bf4d6c     <=
                                             wire_qout_00025_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00025_00003 + 1 :
                                             wire_qout_00025_00003
                                             ;

            I1ca188bcdebbf41d84f7a5220bd1d195  <=  wire_qout_00025_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7b2b617ae67424f54961eebce42de77e     <=
                                             wire_qout_00025_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00025_00004 + 1 :
                                             wire_qout_00025_00004
                                             ;

            Ifc640243288c9b37b7eb9e00351b23f0  <=  wire_qout_00025_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I953f0f8af76f89b2d9ab4abf19fb411d     <=
                                             wire_qout_00025_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00025_00005 + 1 :
                                             wire_qout_00025_00005
                                             ;

            I3d149293f106ae8680c7f4702daa0bd6  <=  wire_qout_00025_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I915b4736dcb20f831d02e48f4e79f008     <=
                                             wire_qout_00025_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00025_00006 + 1 :
                                             wire_qout_00025_00006
                                             ;

            Ie232799bd6c4ec99e24c78f3ad798265  <=  wire_qout_00025_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib7eec587348ae1ca1f00c0a3ad10ad27     <=
                                             wire_qout_00026_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00026_00000 + 1 :
                                             wire_qout_00026_00000
                                             ;

            Ifebcf64858d5e2d07ad7894d6182eb11  <=  wire_qout_00026_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I001a212686304248c8359e5fc01227c0     <=
                                             wire_qout_00026_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00026_00001 + 1 :
                                             wire_qout_00026_00001
                                             ;

            Ibab55499323660588ec82ebd07ab0572  <=  wire_qout_00026_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibb7554e012c0fc1223c29b759c900666     <=
                                             wire_qout_00026_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00026_00002 + 1 :
                                             wire_qout_00026_00002
                                             ;

            I89af7644c48a80d7d22f50b008d35841  <=  wire_qout_00026_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9aeb9c42b54a05be6bf9b7b88b6860ba     <=
                                             wire_qout_00026_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00026_00003 + 1 :
                                             wire_qout_00026_00003
                                             ;

            I0152dc6e6a7acd72a2144623e63998ef  <=  wire_qout_00026_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6a5a5966965b0790b906c6fda71aef80     <=
                                             wire_qout_00026_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00026_00004 + 1 :
                                             wire_qout_00026_00004
                                             ;

            I951dedd7af44c3865a8f36888432d0c9  <=  wire_qout_00026_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic943083ca65ace6c42d73f4234739a06     <=
                                             wire_qout_00026_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00026_00005 + 1 :
                                             wire_qout_00026_00005
                                             ;

            I8188dd7cb03854c6f709de06ff785d91  <=  wire_qout_00026_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id0b321686d4c39621024cf0dd99822dc     <=
                                             wire_qout_00026_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00026_00006 + 1 :
                                             wire_qout_00026_00006
                                             ;

            I3b30b4ab00a49e10a75587aa324d6132  <=  wire_qout_00026_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0839dd3787442f1b79b87e02436bfdce     <=
                                             wire_qout_00027_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00027_00000 + 1 :
                                             wire_qout_00027_00000
                                             ;

            Ie50aca688b3433fad7565998cb900155  <=  wire_qout_00027_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I89e6a9fd97d8aa4dd3b832c3be4697b2     <=
                                             wire_qout_00027_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00027_00001 + 1 :
                                             wire_qout_00027_00001
                                             ;

            I3342fe0c5d3ee5021892d53eb45bde21  <=  wire_qout_00027_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I93d4157f48b132642752220059861e98     <=
                                             wire_qout_00027_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00027_00002 + 1 :
                                             wire_qout_00027_00002
                                             ;

            I5134b762ac428bed07ce102d8927a418  <=  wire_qout_00027_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8fc4faa2891d7fd3479ac1f788f481dc     <=
                                             wire_qout_00027_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00027_00003 + 1 :
                                             wire_qout_00027_00003
                                             ;

            Ic14f948884da19a272a4760ffaab9ea9  <=  wire_qout_00027_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I440f30e9cb4bc89233b46ea00b4cbeb4     <=
                                             wire_qout_00027_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00027_00004 + 1 :
                                             wire_qout_00027_00004
                                             ;

            I46e1047bca2b38e62b4de80d1d2249de  <=  wire_qout_00027_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6568bfd8780c11e0b1b049a01f92abd8     <=
                                             wire_qout_00027_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00027_00005 + 1 :
                                             wire_qout_00027_00005
                                             ;

            I866b30a63b3b5fb708934a1cbb0e1d9a  <=  wire_qout_00027_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibf7dc4da07f9955d5d4c7e1f63f1ad68     <=
                                             wire_qout_00027_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00027_00006 + 1 :
                                             wire_qout_00027_00006
                                             ;

            Iaddc1f2e822fd2fe9d9046d759a82cb4  <=  wire_qout_00027_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7ec1a328587b72a39c462083efea0ee0     <=
                                             wire_qout_00028_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00000 + 1 :
                                             wire_qout_00028_00000
                                             ;

            If9285bf7611bcc5ea6432215c349e021  <=  wire_qout_00028_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iaf028e7ab4dc77a7649f15d603834b5f     <=
                                             wire_qout_00028_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00001 + 1 :
                                             wire_qout_00028_00001
                                             ;

            Id277f5f05551eeb5dec1701056330da1  <=  wire_qout_00028_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I58db79a8e9f0cd1ded379897ba2f27ae     <=
                                             wire_qout_00028_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00002 + 1 :
                                             wire_qout_00028_00002
                                             ;

            I9963d0b24763ed8038b1f3922b8f9548  <=  wire_qout_00028_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6d3cb4ccb4e51c7e6603d0abd1a082c4     <=
                                             wire_qout_00028_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00003 + 1 :
                                             wire_qout_00028_00003
                                             ;

            Ia98de3691917dfb63bebdc3f8655c8be  <=  wire_qout_00028_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I79f75f49ea8a29d684af396014b2f3ab     <=
                                             wire_qout_00028_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00004 + 1 :
                                             wire_qout_00028_00004
                                             ;

            I0bce960fcc58938e6a1e01b912eabbf2  <=  wire_qout_00028_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9c5ecd86bedb189fada40fae9d751a68     <=
                                             wire_qout_00028_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00005 + 1 :
                                             wire_qout_00028_00005
                                             ;

            Ice5f7168aeb940d48093cc9df7cba36b  <=  wire_qout_00028_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iad5f06e1989ead7d306c70a3b02cb8f4     <=
                                             wire_qout_00028_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00006 + 1 :
                                             wire_qout_00028_00006
                                             ;

            I859d795a7d141eb777c1f3c038203794  <=  wire_qout_00028_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If6d1a410df5a4aea6a01337a6074fbd9     <=
                                             wire_qout_00028_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00007 + 1 :
                                             wire_qout_00028_00007
                                             ;

            I0dccb8eaad52ce4d780696a8485420f1  <=  wire_qout_00028_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3bc40a4db14566b5099b14cee5f61135     <=
                                             wire_qout_00028_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00008 + 1 :
                                             wire_qout_00028_00008
                                             ;

            I6d4fc81ced37c159303c243af04d345e  <=  wire_qout_00028_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7e683fd8235d7cfbf4ff407a286f07de     <=
                                             wire_qout_00028_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00009 + 1 :
                                             wire_qout_00028_00009
                                             ;

            Iefdb8bd28839af9413a3906cbfe715e6  <=  wire_qout_00028_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I97afcedf05e588b7976d6005191dc916     <=
                                             wire_qout_00028_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00010 + 1 :
                                             wire_qout_00028_00010
                                             ;

            I0615acb0f7cf79b5f6ae8e91cb525dc9  <=  wire_qout_00028_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib8d8eec0aaa662adf2837c9b705fce7e     <=
                                             wire_qout_00028_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00011 + 1 :
                                             wire_qout_00028_00011
                                             ;

            Ieed4c810a5bb69de112522dcf00b16ed  <=  wire_qout_00028_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icbd765be950123705955e2c5d7ace84b     <=
                                             wire_qout_00028_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00028_00012 + 1 :
                                             wire_qout_00028_00012
                                             ;

            If533578cacb685a95afbb8e1c05d3c07  <=  wire_qout_00028_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I706e8f5617cfae1e6fc83db18c8b5fe3     <=
                                             wire_qout_00029_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00000 + 1 :
                                             wire_qout_00029_00000
                                             ;

            Ia858ff5551286beffd4cf82f876d30ac  <=  wire_qout_00029_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1dd8f8c7f1b673898096b1f3ae383197     <=
                                             wire_qout_00029_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00001 + 1 :
                                             wire_qout_00029_00001
                                             ;

            I4c66570630a650fa7b9bec543f685487  <=  wire_qout_00029_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I10ca8978cf4659265ed25a27d09acc1c     <=
                                             wire_qout_00029_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00002 + 1 :
                                             wire_qout_00029_00002
                                             ;

            If10f33385e236eaba56cbab8c2883399  <=  wire_qout_00029_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iec4656b32460def4a608b6b0f6486af9     <=
                                             wire_qout_00029_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00003 + 1 :
                                             wire_qout_00029_00003
                                             ;

            I7cb58e4c486e683faa4acad4756815d5  <=  wire_qout_00029_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5f4475897d1d58965da1b35fe0ef8c01     <=
                                             wire_qout_00029_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00004 + 1 :
                                             wire_qout_00029_00004
                                             ;

            I452e51cca9acec44e36e4efd21b43034  <=  wire_qout_00029_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ife61469306df3cf220666b187f1496a9     <=
                                             wire_qout_00029_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00005 + 1 :
                                             wire_qout_00029_00005
                                             ;

            Ice0234f25de4ab1f03a3cb01a2d61dbf  <=  wire_qout_00029_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib49319b9dfa4914f92f423ceaf840014     <=
                                             wire_qout_00029_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00006 + 1 :
                                             wire_qout_00029_00006
                                             ;

            I12a18a1f8d4416e9bc8abee6ac3dacfc  <=  wire_qout_00029_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I93ff2f879233cac9b9f0dd2f4c082c09     <=
                                             wire_qout_00029_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00007 + 1 :
                                             wire_qout_00029_00007
                                             ;

            Id17ada8dae3f9810d1892d34f2288859  <=  wire_qout_00029_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I44597d694e9c5d29280e503d72a27c8d     <=
                                             wire_qout_00029_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00008 + 1 :
                                             wire_qout_00029_00008
                                             ;

            Ia2c5fe53cb5b318fa63d09881609655f  <=  wire_qout_00029_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I04a19448c5e75af8021ad02d1a708bb0     <=
                                             wire_qout_00029_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00009 + 1 :
                                             wire_qout_00029_00009
                                             ;

            I579c7926e7b78f4ffc606adc10522f53  <=  wire_qout_00029_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I71a3093121c2f19dcd1412b468652fa8     <=
                                             wire_qout_00029_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00010 + 1 :
                                             wire_qout_00029_00010
                                             ;

            Iffa06a336949f56f4e5a88a06d8b7e60  <=  wire_qout_00029_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3ae09c82029c617034fe6aacbe9e94e6     <=
                                             wire_qout_00029_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00011 + 1 :
                                             wire_qout_00029_00011
                                             ;

            Iaf82668eb49248709540f2f529f1b3e4  <=  wire_qout_00029_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie7af6b3b441f910b000a333afad6c76f     <=
                                             wire_qout_00029_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00029_00012 + 1 :
                                             wire_qout_00029_00012
                                             ;

            I90b3708abdf742370f06cc513ee307e1  <=  wire_qout_00029_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4d71dfea8407aa5b5cbb991bc4fea963     <=
                                             wire_qout_00030_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00000 + 1 :
                                             wire_qout_00030_00000
                                             ;

            Ia17906696bd0e095d7a5297da2e049ea  <=  wire_qout_00030_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1a082caecc831a90e74674ba35da4183     <=
                                             wire_qout_00030_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00001 + 1 :
                                             wire_qout_00030_00001
                                             ;

            I180d4f3b23b518271d7cb8189fbeadc5  <=  wire_qout_00030_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iec1de44616a2354a56ab1f681059d4c5     <=
                                             wire_qout_00030_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00002 + 1 :
                                             wire_qout_00030_00002
                                             ;

            Id79636d195efff260c430978f0bcee9c  <=  wire_qout_00030_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie3c2318e64d0e218c3db557404c4aac8     <=
                                             wire_qout_00030_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00003 + 1 :
                                             wire_qout_00030_00003
                                             ;

            Idbf4ad11ab2a27044193448c8739fec6  <=  wire_qout_00030_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9a251d50f41e51b1a5cc2475f267e8a0     <=
                                             wire_qout_00030_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00004 + 1 :
                                             wire_qout_00030_00004
                                             ;

            I3051f561a5e1131ebf167cb6ccb5adf4  <=  wire_qout_00030_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9b5767a49f7b9dcb8fdaea924835033c     <=
                                             wire_qout_00030_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00005 + 1 :
                                             wire_qout_00030_00005
                                             ;

            I9322a2a61900943075bbc23c72a3f65d  <=  wire_qout_00030_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6ca1e6700a19d03621a193c7240bff54     <=
                                             wire_qout_00030_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00006 + 1 :
                                             wire_qout_00030_00006
                                             ;

            Iedc463e359dd3003d9f7e50f3e858e93  <=  wire_qout_00030_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I931c597ff12bffce581f653346202f83     <=
                                             wire_qout_00030_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00007 + 1 :
                                             wire_qout_00030_00007
                                             ;

            Ie7cfdd25541414ff3f8d6e5d7677fbe5  <=  wire_qout_00030_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia3a2c5d59f6340917ca3933c05ba4678     <=
                                             wire_qout_00030_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00008 + 1 :
                                             wire_qout_00030_00008
                                             ;

            I1e93f0470d2818249f1c28ef2a399a0e  <=  wire_qout_00030_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie83d0a8ee5ed214bc7577467748aaa04     <=
                                             wire_qout_00030_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00009 + 1 :
                                             wire_qout_00030_00009
                                             ;

            I5d6e576b0fa7e3219aaf9ccc345085b8  <=  wire_qout_00030_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iaac29552e5fc65aaf4f0116f917b707c     <=
                                             wire_qout_00030_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00010 + 1 :
                                             wire_qout_00030_00010
                                             ;

            Id962beade26396738ba0e97f67d5e261  <=  wire_qout_00030_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie2c8eac7204b98139c03b6fbfff9af36     <=
                                             wire_qout_00030_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00011 + 1 :
                                             wire_qout_00030_00011
                                             ;

            Id0ab747d92288f23cef793567b2363d1  <=  wire_qout_00030_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ied7fcdaec662cb3c2f89f131986fa102     <=
                                             wire_qout_00030_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00030_00012 + 1 :
                                             wire_qout_00030_00012
                                             ;

            Ie536879e6fa9be65376d7f00e0fc40d0  <=  wire_qout_00030_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib16a17d6430570b45a304d847ee2b11c     <=
                                             wire_qout_00031_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00000 + 1 :
                                             wire_qout_00031_00000
                                             ;

            Ibf312ae4f51fbc44b43848f9df62a45f  <=  wire_qout_00031_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I42169e454756fe4d1c5f17f2eeb2e091     <=
                                             wire_qout_00031_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00001 + 1 :
                                             wire_qout_00031_00001
                                             ;

            Icfc03646b36b971b9fa57d04a26dbfc4  <=  wire_qout_00031_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6fde38a3a92e06fa77123e3279813c41     <=
                                             wire_qout_00031_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00002 + 1 :
                                             wire_qout_00031_00002
                                             ;

            I4f134c0669b5a6a8c7e03be7eee30c6c  <=  wire_qout_00031_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id8ee16437e8d6d6da6d37440e04097b6     <=
                                             wire_qout_00031_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00003 + 1 :
                                             wire_qout_00031_00003
                                             ;

            I6c765e677f42fe600b848698c8a78349  <=  wire_qout_00031_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibf249d8e5acced9b064132575f40e001     <=
                                             wire_qout_00031_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00004 + 1 :
                                             wire_qout_00031_00004
                                             ;

            I284b23051c85300c2a1e3afe8f25e99e  <=  wire_qout_00031_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I580659084e3d17b48de6b1c66154fcf5     <=
                                             wire_qout_00031_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00005 + 1 :
                                             wire_qout_00031_00005
                                             ;

            I9b560d9baf8a7422b0dd84720e924ced  <=  wire_qout_00031_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7a14e45d43ab77b265501902152c8616     <=
                                             wire_qout_00031_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00006 + 1 :
                                             wire_qout_00031_00006
                                             ;

            I457ae11ad90c8478751eb4b42764e158  <=  wire_qout_00031_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I81ba868784103e0eb05a44d981d4d666     <=
                                             wire_qout_00031_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00007 + 1 :
                                             wire_qout_00031_00007
                                             ;

            I2b7822d5d77aaed61eee87570564df76  <=  wire_qout_00031_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic6b88783957cbaf253648a30b22f6b1c     <=
                                             wire_qout_00031_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00008 + 1 :
                                             wire_qout_00031_00008
                                             ;

            Ibdad0ab78e4404c852e60a2b04c3a5f6  <=  wire_qout_00031_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4103c218a85a1d08db5c4f4b5686b2e5     <=
                                             wire_qout_00031_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00009 + 1 :
                                             wire_qout_00031_00009
                                             ;

            Ic4efba3932e598784f5b9ad6ad04772d  <=  wire_qout_00031_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0e6c0958af503e4a120a49d02a432863     <=
                                             wire_qout_00031_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00010 + 1 :
                                             wire_qout_00031_00010
                                             ;

            Ia03836a4e93d2f36513227d1dfaea0fa  <=  wire_qout_00031_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8f76b31e8f15c0e5fe24dcb723418111     <=
                                             wire_qout_00031_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00011 + 1 :
                                             wire_qout_00031_00011
                                             ;

            I138fb0c48f2d27e3315e237d9e61d653  <=  wire_qout_00031_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id1457221b58344b60070aa026436df2c     <=
                                             wire_qout_00031_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00031_00012 + 1 :
                                             wire_qout_00031_00012
                                             ;

            Id0b1c46fa4caa63a4c63a44ba3c5ef8a  <=  wire_qout_00031_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icc31966508e03d8869e81d8aeb243705     <=
                                             wire_qout_00032_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00032_00000 + 1 :
                                             wire_qout_00032_00000
                                             ;

            I3566033cf5c9a06977c9182925750707  <=  wire_qout_00032_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9dcccf542ba434b6e0fde6f012f98f92     <=
                                             wire_qout_00032_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00032_00001 + 1 :
                                             wire_qout_00032_00001
                                             ;

            I02812a8a833bb69eb168a1004b6fafdf  <=  wire_qout_00032_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I51ccbb824a5e1e340eefd173c4491728     <=
                                             wire_qout_00032_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00032_00002 + 1 :
                                             wire_qout_00032_00002
                                             ;

            Ie886c5effc85f1fe0b6411db4a2cde77  <=  wire_qout_00032_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib7ae1730dcd8bc708bbfcc6a9f97ac66     <=
                                             wire_qout_00032_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00032_00003 + 1 :
                                             wire_qout_00032_00003
                                             ;

            Ibab1d13cd6a4f7b0c79c9f845339e53f  <=  wire_qout_00032_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4714f5c91203fcfa552f0fcf71b87442     <=
                                             wire_qout_00032_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00032_00004 + 1 :
                                             wire_qout_00032_00004
                                             ;

            I7b813d83b13bb7bc13940cf5714c06ba  <=  wire_qout_00032_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3b6d1e84fdd1019249886fa5fe65895b     <=
                                             wire_qout_00032_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00032_00005 + 1 :
                                             wire_qout_00032_00005
                                             ;

            I09031235f61238b0e32ff52641aab70e  <=  wire_qout_00032_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia8a7d4207dbabc7970bf36f3fe74f72d     <=
                                             wire_qout_00033_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00033_00000 + 1 :
                                             wire_qout_00033_00000
                                             ;

            I5402fd208dc7ca81dfd2920a9cfa2715  <=  wire_qout_00033_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I84047457b43ef33874f4550c3b773460     <=
                                             wire_qout_00033_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00033_00001 + 1 :
                                             wire_qout_00033_00001
                                             ;

            Ia01c82761aeb124cd92fb15ee367ee8b  <=  wire_qout_00033_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5e51563c3e69beca0b463742e6e5f9ee     <=
                                             wire_qout_00033_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00033_00002 + 1 :
                                             wire_qout_00033_00002
                                             ;

            Ib1a40247057324b0bd810c844bf11f51  <=  wire_qout_00033_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6c8d14e31c80811ccab1b6ab09d28089     <=
                                             wire_qout_00033_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00033_00003 + 1 :
                                             wire_qout_00033_00003
                                             ;

            Ied8bd4b6fd0e4fbcced6d20eb7435f55  <=  wire_qout_00033_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I50b3b7490c9b65b6e662cc86b163a2df     <=
                                             wire_qout_00033_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00033_00004 + 1 :
                                             wire_qout_00033_00004
                                             ;

            I4ee312036de8c08300c358edcff1e1e9  <=  wire_qout_00033_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8351a2110a3d73ad8803cf17e3317017     <=
                                             wire_qout_00033_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00033_00005 + 1 :
                                             wire_qout_00033_00005
                                             ;

            I477a920e2326828bf026b0a6b6a18e2b  <=  wire_qout_00033_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1e6c696951688d581f21ab2302593335     <=
                                             wire_qout_00034_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00034_00000 + 1 :
                                             wire_qout_00034_00000
                                             ;

            Ic11a6b77b84c44180eb99220a0c4c9f6  <=  wire_qout_00034_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie9840e28133eebdca0be313552195c7b     <=
                                             wire_qout_00034_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00034_00001 + 1 :
                                             wire_qout_00034_00001
                                             ;

            If0970d9f7b053fce3ced3521b4885588  <=  wire_qout_00034_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I82812258a8032e273cab7139266be1b6     <=
                                             wire_qout_00034_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00034_00002 + 1 :
                                             wire_qout_00034_00002
                                             ;

            Ic7ebdc317c978eb275eca41d5b9106a5  <=  wire_qout_00034_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I27ab6fd9927518e29ed36d7a7a241498     <=
                                             wire_qout_00034_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00034_00003 + 1 :
                                             wire_qout_00034_00003
                                             ;

            Ibe3d3e6bc58efc2e9d9eb1f96cdfe424  <=  wire_qout_00034_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I05b0f33a3808ac53b29d8d8309447650     <=
                                             wire_qout_00034_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00034_00004 + 1 :
                                             wire_qout_00034_00004
                                             ;

            I1dd4671765f8826c2fe20c592c5e32c8  <=  wire_qout_00034_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If150ebf242231f0d22c996a71552f6eb     <=
                                             wire_qout_00034_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00034_00005 + 1 :
                                             wire_qout_00034_00005
                                             ;

            I6cde57127c5bd2732e71ecb7738fad6d  <=  wire_qout_00034_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If2d0a2b58510715e74787cb60719cb5b     <=
                                             wire_qout_00035_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00035_00000 + 1 :
                                             wire_qout_00035_00000
                                             ;

            If6ce2fa9f0b8bc74442ed8262b5089cf  <=  wire_qout_00035_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib6745a6d17034a29501e022bd846bf2f     <=
                                             wire_qout_00035_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00035_00001 + 1 :
                                             wire_qout_00035_00001
                                             ;

            Ib0001d7298ad1f3b1c7603173a70d8b5  <=  wire_qout_00035_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iae09c127dfe86c9f7bdbeff447c777f5     <=
                                             wire_qout_00035_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00035_00002 + 1 :
                                             wire_qout_00035_00002
                                             ;

            I05e739fc87e962848f265e2c73338cac  <=  wire_qout_00035_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I742128de6b237ed48e3a7ccd3788f0d7     <=
                                             wire_qout_00035_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00035_00003 + 1 :
                                             wire_qout_00035_00003
                                             ;

            Iaaaf373f7e6f55214915b93da9bd71d3  <=  wire_qout_00035_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id5e8fda13ba8f6d95d694d0f30da75bb     <=
                                             wire_qout_00035_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00035_00004 + 1 :
                                             wire_qout_00035_00004
                                             ;

            I47b0847946b0e00961233ac0101fa2a7  <=  wire_qout_00035_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1aa5a04e40f9b1685c77e4d101c3ccf4     <=
                                             wire_qout_00035_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00035_00005 + 1 :
                                             wire_qout_00035_00005
                                             ;

            I2f23d4cdb6f5f827513aa60266936e4f  <=  wire_qout_00035_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ife1adea26d13bc299bb2de241ad4a6ea     <=
                                             wire_qout_00036_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00036_00000 + 1 :
                                             wire_qout_00036_00000
                                             ;

            Ia67f9b902a21de0414eb8dda52171991  <=  wire_qout_00036_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifcf6c761f0f253921710af87ab1d2247     <=
                                             wire_qout_00036_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00036_00001 + 1 :
                                             wire_qout_00036_00001
                                             ;

            I87b10521099179c18652c86d5887c908  <=  wire_qout_00036_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1478e6a9113c124bdc4361908af6643f     <=
                                             wire_qout_00036_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00036_00002 + 1 :
                                             wire_qout_00036_00002
                                             ;

            I84057a3b319ab3d6a2ed8f2310f970fc  <=  wire_qout_00036_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0afd42151925883835844cf5deef6156     <=
                                             wire_qout_00036_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00036_00003 + 1 :
                                             wire_qout_00036_00003
                                             ;

            I67d57e38df8cb35ca686ac2eb44e233e  <=  wire_qout_00036_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2b4ab0aadffb3a1bb86f45ebc8acf085     <=
                                             wire_qout_00036_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00036_00004 + 1 :
                                             wire_qout_00036_00004
                                             ;

            I23955b54e486f0f0d21a2809a9472b86  <=  wire_qout_00036_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iffa867719ba9c31a8756cc5e6bf81147     <=
                                             wire_qout_00036_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00036_00005 + 1 :
                                             wire_qout_00036_00005
                                             ;

            I1e11f0088959aa40b4ad1a047b59caf4  <=  wire_qout_00036_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibb62b6cb003f0d5549c864075f23d19b     <=
                                             wire_qout_00036_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00036_00006 + 1 :
                                             wire_qout_00036_00006
                                             ;

            I68c35d63dc95baff41b4dc27a86d2342  <=  wire_qout_00036_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3690d101ae99f258cc58b4482cc378c8     <=
                                             wire_qout_00036_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00036_00007 + 1 :
                                             wire_qout_00036_00007
                                             ;

            I837183265ee22d080e81fea468ab0887  <=  wire_qout_00036_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id597e95ce8a168ab67890085a26870d0     <=
                                             wire_qout_00037_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00037_00000 + 1 :
                                             wire_qout_00037_00000
                                             ;

            I413b1c1985a6c9c6f202e85ff901e3a8  <=  wire_qout_00037_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I98df60eb8f65641f9cccce4023be905c     <=
                                             wire_qout_00037_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00037_00001 + 1 :
                                             wire_qout_00037_00001
                                             ;

            Ic32c6734132776c290155a80025fe366  <=  wire_qout_00037_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibcb4fbdee372353b79c460cdeafdfe4e     <=
                                             wire_qout_00037_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00037_00002 + 1 :
                                             wire_qout_00037_00002
                                             ;

            I624958486d181501c7a8ec2642cb503c  <=  wire_qout_00037_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I74dbf75966d047a4a9e91c1bc793666f     <=
                                             wire_qout_00037_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00037_00003 + 1 :
                                             wire_qout_00037_00003
                                             ;

            I04864c28351edb33b61a103add6fb875  <=  wire_qout_00037_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I79b8d9f9447c4c1b551ec6c1e8903040     <=
                                             wire_qout_00037_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00037_00004 + 1 :
                                             wire_qout_00037_00004
                                             ;

            Ida3dd5e990ce3c237e9628a9a090901e  <=  wire_qout_00037_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib34b66548621fabe0753223712b1369f     <=
                                             wire_qout_00037_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00037_00005 + 1 :
                                             wire_qout_00037_00005
                                             ;

            Id182a776b03f48fb139c28194ae7ab6b  <=  wire_qout_00037_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie5b3eb4c00bedfaecc3215d43ff28362     <=
                                             wire_qout_00037_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00037_00006 + 1 :
                                             wire_qout_00037_00006
                                             ;

            I0c5539373b3868d0664a92157b4b4226  <=  wire_qout_00037_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icf3a1b0b6dbcf959b44379024f3c4169     <=
                                             wire_qout_00037_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00037_00007 + 1 :
                                             wire_qout_00037_00007
                                             ;

            Ic0191941cb968bbd7644c21767423d2e  <=  wire_qout_00037_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I918c2bbe7c71f8c6a07b0bad8811f4e7     <=
                                             wire_qout_00038_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00038_00000 + 1 :
                                             wire_qout_00038_00000
                                             ;

            I163cf58b9a308e0439a8dc7c1526e6b5  <=  wire_qout_00038_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iedd960a21b1c08b4a5293cff200218b3     <=
                                             wire_qout_00038_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00038_00001 + 1 :
                                             wire_qout_00038_00001
                                             ;

            Ie08ad9bd71329858c1742c8f571a1c36  <=  wire_qout_00038_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If9722c28747df3a59b0ecf8200907e98     <=
                                             wire_qout_00038_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00038_00002 + 1 :
                                             wire_qout_00038_00002
                                             ;

            I3c10d579f80bd0106506ad047d75f188  <=  wire_qout_00038_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib83df72c8b73a333d0699a8bbbec16be     <=
                                             wire_qout_00038_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00038_00003 + 1 :
                                             wire_qout_00038_00003
                                             ;

            Ieca2767ac27170058499d83016447aa7  <=  wire_qout_00038_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ide3798a77f709a9f694523338b081f70     <=
                                             wire_qout_00038_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00038_00004 + 1 :
                                             wire_qout_00038_00004
                                             ;

            Ib9c194ec16f435a9357cb344cf25bdcc  <=  wire_qout_00038_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0a9722a805604433562f85c62b168b96     <=
                                             wire_qout_00038_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00038_00005 + 1 :
                                             wire_qout_00038_00005
                                             ;

            Ic920452d5997a8477724fa78c86c0fba  <=  wire_qout_00038_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If9480ec13cd538ed03a43e56bd6264a6     <=
                                             wire_qout_00038_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00038_00006 + 1 :
                                             wire_qout_00038_00006
                                             ;

            I6eea5fde8e2517554ad6ba25018572dc  <=  wire_qout_00038_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I433ecf86b7704c5552e5fb5cafe0d529     <=
                                             wire_qout_00038_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00038_00007 + 1 :
                                             wire_qout_00038_00007
                                             ;

            I9ad2f6fd2d7f68011fc926ec9abd5c34  <=  wire_qout_00038_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8326f0b2d25139609e2c5e466724f224     <=
                                             wire_qout_00039_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00039_00000 + 1 :
                                             wire_qout_00039_00000
                                             ;

            Ied33f18cbb778d5ba744d249f91c950b  <=  wire_qout_00039_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibbe211d9955cdf2810c9003d1fb78074     <=
                                             wire_qout_00039_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00039_00001 + 1 :
                                             wire_qout_00039_00001
                                             ;

            Ibabf61085ca7af8dfc7927b3656a76f7  <=  wire_qout_00039_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If15e950b569a92b590127d0ca6f20a16     <=
                                             wire_qout_00039_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00039_00002 + 1 :
                                             wire_qout_00039_00002
                                             ;

            Iddc5b5b4501f9f13bcaf22081e5a70f4  <=  wire_qout_00039_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I03e0532841ba39eb1d4ae823c4de2f7d     <=
                                             wire_qout_00039_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00039_00003 + 1 :
                                             wire_qout_00039_00003
                                             ;

            I67f87fbb746dd937fffc534c596f36c4  <=  wire_qout_00039_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1be81a7b73987ee023e396cec87312d1     <=
                                             wire_qout_00039_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00039_00004 + 1 :
                                             wire_qout_00039_00004
                                             ;

            I45bdd0cfe107da0d57cad1333bf95e3b  <=  wire_qout_00039_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4ce1a767a78673590c4074f3f03bad8d     <=
                                             wire_qout_00039_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00039_00005 + 1 :
                                             wire_qout_00039_00005
                                             ;

            I4d54dd2ee2f32909098d3cc2b6689220  <=  wire_qout_00039_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I57806bb7da625881e68ae315543f70d6     <=
                                             wire_qout_00039_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00039_00006 + 1 :
                                             wire_qout_00039_00006
                                             ;

            I7bfb4c5d9e22d1bd8811844d9c74dff8  <=  wire_qout_00039_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8b0ab476b4790150575abb06bcdce2b3     <=
                                             wire_qout_00039_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00039_00007 + 1 :
                                             wire_qout_00039_00007
                                             ;

            Ib9d58222da98f29fa302b4896594fe26  <=  wire_qout_00039_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8846a8961b7d557df4fc62dada679c33     <=
                                             wire_qout_00040_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00040_00000 + 1 :
                                             wire_qout_00040_00000
                                             ;

            Iea3e35ece9fdb3aff3b9ff5369e9a7e0  <=  wire_qout_00040_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7909a0f96a92e93f95023cddc742a5eb     <=
                                             wire_qout_00040_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00040_00001 + 1 :
                                             wire_qout_00040_00001
                                             ;

            Ic44eab478be232721e7a43d14beca32f  <=  wire_qout_00040_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I43ac4857544c0fb79d04e850435ef673     <=
                                             wire_qout_00040_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00040_00002 + 1 :
                                             wire_qout_00040_00002
                                             ;

            Ifab075b1437495268b6a3be4cb022e71  <=  wire_qout_00040_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia6dfa47c465325c1d9fb9b9c5ce08f01     <=
                                             wire_qout_00040_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00040_00003 + 1 :
                                             wire_qout_00040_00003
                                             ;

            I2919272e9ae3996a3e1d602ff72ba86d  <=  wire_qout_00040_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2e9eda5bea0cc3d88359ce8a7a82f21f     <=
                                             wire_qout_00040_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00040_00004 + 1 :
                                             wire_qout_00040_00004
                                             ;

            Ib6fbe376477afa58bfcc17a8564f78b2  <=  wire_qout_00040_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I53ec2486418e41b2ccfa8fd82777eaf0     <=
                                             wire_qout_00040_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00040_00005 + 1 :
                                             wire_qout_00040_00005
                                             ;

            I659322a9fd0d5eac514437b02e0491b3  <=  wire_qout_00040_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I18387c05cef21970ecbc39c20a87aafb     <=
                                             wire_qout_00040_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00040_00006 + 1 :
                                             wire_qout_00040_00006
                                             ;

            Ic68f500938d80460ffdb33a0adc48298  <=  wire_qout_00040_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2b23eae78cb925008ad59f45e80e165b     <=
                                             wire_qout_00040_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00040_00007 + 1 :
                                             wire_qout_00040_00007
                                             ;

            If5ae6fbf843fdeee17945bc5ce81aec8  <=  wire_qout_00040_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic69eb7677638a90b7a54389d47be46de     <=
                                             wire_qout_00040_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00040_00008 + 1 :
                                             wire_qout_00040_00008
                                             ;

            I94460b6ce7b776bcc5eca149eab80c26  <=  wire_qout_00040_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8cb9a216f4da7c27f678386cb214c59d     <=
                                             wire_qout_00041_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00041_00000 + 1 :
                                             wire_qout_00041_00000
                                             ;

            I3347717ba9556e69de30ce7533d4f5a4  <=  wire_qout_00041_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I48cb720a6323697084ac3bbd8fcadfcb     <=
                                             wire_qout_00041_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00041_00001 + 1 :
                                             wire_qout_00041_00001
                                             ;

            I2db290170ddae8dc52ce07edaf48b365  <=  wire_qout_00041_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib8dc3c1885c92cdcce7fcb58d65d03e7     <=
                                             wire_qout_00041_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00041_00002 + 1 :
                                             wire_qout_00041_00002
                                             ;

            Idd775d9fe6fa8dbdbfb07d4071b9caa5  <=  wire_qout_00041_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic3aa51a5c758405fa6e2dbed707555b2     <=
                                             wire_qout_00041_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00041_00003 + 1 :
                                             wire_qout_00041_00003
                                             ;

            I6cbc06919b9c695d99621db6f8d768cb  <=  wire_qout_00041_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4d418179c859feb8bc7d750416bb1004     <=
                                             wire_qout_00041_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00041_00004 + 1 :
                                             wire_qout_00041_00004
                                             ;

            I5b8a1e1a6b904b0f6822c224ee0486e3  <=  wire_qout_00041_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If207b2adc6f668f85cb76bf54673fe18     <=
                                             wire_qout_00041_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00041_00005 + 1 :
                                             wire_qout_00041_00005
                                             ;

            I3f5053e519a928640ae49cf4e5b39d1e  <=  wire_qout_00041_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib08b8067ea75e210e83526ca4a37217e     <=
                                             wire_qout_00041_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00041_00006 + 1 :
                                             wire_qout_00041_00006
                                             ;

            I7c965c047d862c973d09a81abe03a845  <=  wire_qout_00041_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I95b30f641cbf7bec1886643c4468017d     <=
                                             wire_qout_00041_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00041_00007 + 1 :
                                             wire_qout_00041_00007
                                             ;

            I9b8023f4dced915cd52c91bc9d4ed78f  <=  wire_qout_00041_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1978531a6f8d1d25ee6d404025ec4753     <=
                                             wire_qout_00041_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00041_00008 + 1 :
                                             wire_qout_00041_00008
                                             ;

            Idc6b6357741c9887a9db1037ccc2d922  <=  wire_qout_00041_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6c9698ba88db16b8d22ccebd58cc541d     <=
                                             wire_qout_00042_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00042_00000 + 1 :
                                             wire_qout_00042_00000
                                             ;

            Ibe97860165dc5d9a076ebd935385ae51  <=  wire_qout_00042_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0d8ac5e09b200a55bf5ba6f834cc9174     <=
                                             wire_qout_00042_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00042_00001 + 1 :
                                             wire_qout_00042_00001
                                             ;

            I777ee54ff20d0544af18ad8a870d6915  <=  wire_qout_00042_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib58b7d3d77a54ff1a180c6fa5f1400e6     <=
                                             wire_qout_00042_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00042_00002 + 1 :
                                             wire_qout_00042_00002
                                             ;

            Id18c5a1d4eaa73a94e699e5f9e3c3d35  <=  wire_qout_00042_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icf6b990098b7ab91800bfcf1e643153c     <=
                                             wire_qout_00042_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00042_00003 + 1 :
                                             wire_qout_00042_00003
                                             ;

            I72939e49bf2d9c6a84e404419fc644a1  <=  wire_qout_00042_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie4308b9ac6fb6de9329ba02b1eeb0e8a     <=
                                             wire_qout_00042_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00042_00004 + 1 :
                                             wire_qout_00042_00004
                                             ;

            I57b7b48f13436b19a8d6a47e014eb41f  <=  wire_qout_00042_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I01d4f02a356c51d7e4e1993de0d8eebd     <=
                                             wire_qout_00042_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00042_00005 + 1 :
                                             wire_qout_00042_00005
                                             ;

            Ia3ef2f70c5abaa852586a33c505aee0d  <=  wire_qout_00042_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I36c351e3641b01cc43e1dd5de0a649e5     <=
                                             wire_qout_00042_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00042_00006 + 1 :
                                             wire_qout_00042_00006
                                             ;

            I6d423a7d17e05a3c597ec6ef6c5a7cba  <=  wire_qout_00042_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4fc983e94c5b8f7bafca61fb0d351c08     <=
                                             wire_qout_00042_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00042_00007 + 1 :
                                             wire_qout_00042_00007
                                             ;

            I48e3309c61918c3991852b45d9c72ea5  <=  wire_qout_00042_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1fcb82fdf96cda14a55fa6358cb62c1e     <=
                                             wire_qout_00042_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00042_00008 + 1 :
                                             wire_qout_00042_00008
                                             ;

            I472352e7027b9df2fa957d9fd68443ff  <=  wire_qout_00042_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I665e54ea6bdca483149d3b7f3ee42a2b     <=
                                             wire_qout_00043_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00043_00000 + 1 :
                                             wire_qout_00043_00000
                                             ;

            Idbbf2ce4a30787c5f07c3b908a73da75  <=  wire_qout_00043_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I925df2307b5af6d1b166e5435641d3bd     <=
                                             wire_qout_00043_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00043_00001 + 1 :
                                             wire_qout_00043_00001
                                             ;

            Ibc9a860879ccc58c815b9f6caa23320a  <=  wire_qout_00043_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9b14f48aa357d09e460a445da86cdf89     <=
                                             wire_qout_00043_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00043_00002 + 1 :
                                             wire_qout_00043_00002
                                             ;

            Ia71cf07b645c58cffe33be1a9a960eb2  <=  wire_qout_00043_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I78e94ecb6c92fa8ee24edaff33b6f82d     <=
                                             wire_qout_00043_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00043_00003 + 1 :
                                             wire_qout_00043_00003
                                             ;

            I0ceb14ac0187d804f9692e0c55b8e941  <=  wire_qout_00043_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5ebeb9ce5adee72a7c9527ea6d3a3028     <=
                                             wire_qout_00043_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00043_00004 + 1 :
                                             wire_qout_00043_00004
                                             ;

            Ief18a19d451f05f6051e3cc8de16d73c  <=  wire_qout_00043_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I90d7b28ec09142ca8086836fc0c5ea0d     <=
                                             wire_qout_00043_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00043_00005 + 1 :
                                             wire_qout_00043_00005
                                             ;

            I30be0b18e4415ca50f2d8149efaaafe6  <=  wire_qout_00043_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I27d9985415e6d0b117e5a4c2863aa7f8     <=
                                             wire_qout_00043_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00043_00006 + 1 :
                                             wire_qout_00043_00006
                                             ;

            I7ec15b73b2811b44e1e50c74a9f921e9  <=  wire_qout_00043_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idf9b563e5d10c2bdbcc07e81d74467eb     <=
                                             wire_qout_00043_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00043_00007 + 1 :
                                             wire_qout_00043_00007
                                             ;

            I0fd2f706e374a4eb57ee26ab50201e15  <=  wire_qout_00043_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie351922194483938302ff6cafc477e4a     <=
                                             wire_qout_00043_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00043_00008 + 1 :
                                             wire_qout_00043_00008
                                             ;

            I44f170d02bae7fe044456e125a98451d  <=  wire_qout_00043_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifb2da5faf236ca8636677bc1dc35c4db     <=
                                             wire_qout_00044_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00000 + 1 :
                                             wire_qout_00044_00000
                                             ;

            I30c0fcd89e0cc7c5fa348df7b4fa2ccf  <=  wire_qout_00044_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie15825d216685ae241b528fa9c158ff3     <=
                                             wire_qout_00044_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00001 + 1 :
                                             wire_qout_00044_00001
                                             ;

            I13a98f98c54b2e412cd88c96f016c41b  <=  wire_qout_00044_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id92c2d8bc61245c0c8e40bec2424c3c8     <=
                                             wire_qout_00044_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00002 + 1 :
                                             wire_qout_00044_00002
                                             ;

            I9890f7fc708c7b8cf460849b4a30025b  <=  wire_qout_00044_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icd9fd8d7114b6e894dbee493b6797df6     <=
                                             wire_qout_00044_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00003 + 1 :
                                             wire_qout_00044_00003
                                             ;

            I5e69e930a318dcb0594a823b3129d650  <=  wire_qout_00044_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I29ff688c085f2b18e7a3af969f18af76     <=
                                             wire_qout_00044_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00004 + 1 :
                                             wire_qout_00044_00004
                                             ;

            I403303228c0df825f67436f4a7e64061  <=  wire_qout_00044_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6d56db9fcfe69dfcd747521a1ff62297     <=
                                             wire_qout_00044_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00005 + 1 :
                                             wire_qout_00044_00005
                                             ;

            I946246be5b4745508b7d4b578f83aaa2  <=  wire_qout_00044_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2f17f7c79a0118b39a63894917c6affa     <=
                                             wire_qout_00044_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00006 + 1 :
                                             wire_qout_00044_00006
                                             ;

            I95f0acd4f955058041c035789c3a4d99  <=  wire_qout_00044_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7350af5d5ee09ad28c459e3674a829ab     <=
                                             wire_qout_00044_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00007 + 1 :
                                             wire_qout_00044_00007
                                             ;

            I4082b3564c1949a19ed35bd5a88e1ef4  <=  wire_qout_00044_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I67b6415c5135e3d6a41d56d98d3f8315     <=
                                             wire_qout_00044_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00008 + 1 :
                                             wire_qout_00044_00008
                                             ;

            Ia7606050c683ecefc510ba92ac539a9c  <=  wire_qout_00044_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4a6fffd8bb7244599383f2aa3a1c8916     <=
                                             wire_qout_00044_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00009 + 1 :
                                             wire_qout_00044_00009
                                             ;

            I5446c1c323774715371c73bd1be66697  <=  wire_qout_00044_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7dbcd21016231546b76aab175cac9f74     <=
                                             wire_qout_00044_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00010 + 1 :
                                             wire_qout_00044_00010
                                             ;

            I3a8e9e7d2cd6751e8500a5567cef5acc  <=  wire_qout_00044_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9aeff3dc44ed0d0f32518590a900dcc9     <=
                                             wire_qout_00044_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00011 + 1 :
                                             wire_qout_00044_00011
                                             ;

            I621b20d29d3a9a9f41065bc3c3bbd2d8  <=  wire_qout_00044_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I988b7d5d56d22d2c77c5c8c125129a50     <=
                                             wire_qout_00044_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00012 + 1 :
                                             wire_qout_00044_00012
                                             ;

            I263aad78110a1136eb7012c6983b2a8d  <=  wire_qout_00044_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iff35cd97f2a6d37a7861b9cc1a655ef5     <=
                                             wire_qout_00044_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00013 + 1 :
                                             wire_qout_00044_00013
                                             ;

            If4308ed204e33952c9931f8fe257aca4  <=  wire_qout_00044_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifb3f2a1bedfe41c73d198046a2a3f177     <=
                                             wire_qout_00044_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00014 + 1 :
                                             wire_qout_00044_00014
                                             ;

            Iddcfab4a7022e0f12fd20cb34e9b9d02  <=  wire_qout_00044_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I37ddc6ccbc188a3eb8c33a501de820be     <=
                                             wire_qout_00044_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00044_00015 + 1 :
                                             wire_qout_00044_00015
                                             ;

            I759409e242eaeb144a53e630a8cfd514  <=  wire_qout_00044_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ica608f1136da397e2ab61bd4a5d83201     <=
                                             wire_qout_00045_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00000 + 1 :
                                             wire_qout_00045_00000
                                             ;

            I5f96a68d20e3ebc71dad4b43305baa20  <=  wire_qout_00045_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I80636a3df4541bf29780bcb4d0ee48f9     <=
                                             wire_qout_00045_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00001 + 1 :
                                             wire_qout_00045_00001
                                             ;

            I5d92fdff96b9cd64f3af2b28b13e9956  <=  wire_qout_00045_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9ad99d544187db3cc7090b92c9933a31     <=
                                             wire_qout_00045_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00002 + 1 :
                                             wire_qout_00045_00002
                                             ;

            Iab2f643f81921ed8464e1bbd9fa8c68e  <=  wire_qout_00045_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iaa8a2b6fcd469869efcf0b75ca38e68f     <=
                                             wire_qout_00045_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00003 + 1 :
                                             wire_qout_00045_00003
                                             ;

            I17d7f36fdade16dbcf621fe302bd7e57  <=  wire_qout_00045_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9a171d2d8eee362a0073ab7b139d3037     <=
                                             wire_qout_00045_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00004 + 1 :
                                             wire_qout_00045_00004
                                             ;

            I23afd747ecece714e32fbb896b5c022a  <=  wire_qout_00045_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I84cdcba86bc5991feb391003cd7be40b     <=
                                             wire_qout_00045_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00005 + 1 :
                                             wire_qout_00045_00005
                                             ;

            I388528eaf83566cc56b23485a9c05962  <=  wire_qout_00045_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If9e5c3a848acce5daf570458f78f6aad     <=
                                             wire_qout_00045_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00006 + 1 :
                                             wire_qout_00045_00006
                                             ;

            Iea424dd9d8916c4951b8746408b8a521  <=  wire_qout_00045_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I73247d4348333f67a491fc607b15af0e     <=
                                             wire_qout_00045_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00007 + 1 :
                                             wire_qout_00045_00007
                                             ;

            I73bbf90b625d56f663ad10f9d21d8e76  <=  wire_qout_00045_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I021c745eee4b85a2cd91d9d8d2b18b2c     <=
                                             wire_qout_00045_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00008 + 1 :
                                             wire_qout_00045_00008
                                             ;

            I41796b587316c600bf583edc62649bd8  <=  wire_qout_00045_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1381c0a0bd28b1c5542992084635b355     <=
                                             wire_qout_00045_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00009 + 1 :
                                             wire_qout_00045_00009
                                             ;

            I7009c18515dd43d8dd2e5d1ee6779641  <=  wire_qout_00045_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie74eeddc21428254a8fc4c3e293b5eb7     <=
                                             wire_qout_00045_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00010 + 1 :
                                             wire_qout_00045_00010
                                             ;

            I797c9cb725f88c07be28f017871d17f8  <=  wire_qout_00045_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib1d0f94258b45de4bfe610086d8990c5     <=
                                             wire_qout_00045_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00011 + 1 :
                                             wire_qout_00045_00011
                                             ;

            I06b48093d4c9b0327c3efc6fa4ca7daf  <=  wire_qout_00045_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I138d6d5d60df37870cdbb1d9c51a94af     <=
                                             wire_qout_00045_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00012 + 1 :
                                             wire_qout_00045_00012
                                             ;

            I04c734eb876aa722e84d6b9edd297978  <=  wire_qout_00045_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I706378735e63e15c8d5395446ea41db8     <=
                                             wire_qout_00045_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00013 + 1 :
                                             wire_qout_00045_00013
                                             ;

            Ifb89e7ad8ef661959d82b7c22f187243  <=  wire_qout_00045_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If8680a7fc4f5532a660006bf4ca6a66e     <=
                                             wire_qout_00045_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00014 + 1 :
                                             wire_qout_00045_00014
                                             ;

            Id1dce2b9eafc35fa71df33ada4aac539  <=  wire_qout_00045_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic59d1ff3051a95166c3c2d5a2881221b     <=
                                             wire_qout_00045_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00045_00015 + 1 :
                                             wire_qout_00045_00015
                                             ;

            Ied19cb51636bfb029ba8a2c390f97105  <=  wire_qout_00045_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I54a551af28c505601cdfaf8faaa94afb     <=
                                             wire_qout_00046_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00000 + 1 :
                                             wire_qout_00046_00000
                                             ;

            Ie46b71f55aef4d00168202431d47dce0  <=  wire_qout_00046_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6a3124c03eb83d41c16704133bd1cfde     <=
                                             wire_qout_00046_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00001 + 1 :
                                             wire_qout_00046_00001
                                             ;

            I8c0c1a0a35f4f7a688f516c567242d39  <=  wire_qout_00046_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie9ee27b9761af611ab96f0010abd47a3     <=
                                             wire_qout_00046_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00002 + 1 :
                                             wire_qout_00046_00002
                                             ;

            I53222c82827cab7c770e057ae91bc10e  <=  wire_qout_00046_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I305436919f84066a22ab1417ebabd737     <=
                                             wire_qout_00046_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00003 + 1 :
                                             wire_qout_00046_00003
                                             ;

            I8015717cd36aabbf2cf4aa3a5c234690  <=  wire_qout_00046_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I78e63717f436493b756efa32d66cdefd     <=
                                             wire_qout_00046_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00004 + 1 :
                                             wire_qout_00046_00004
                                             ;

            Ic0c13c9a929c8c46e8702cef74de8955  <=  wire_qout_00046_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic965ba971642db19ca773eb68dc0b9bf     <=
                                             wire_qout_00046_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00005 + 1 :
                                             wire_qout_00046_00005
                                             ;

            I71d7f72d83b7410de31e09ea96adb95c  <=  wire_qout_00046_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I579480a66a5f6331fb46de13090ce888     <=
                                             wire_qout_00046_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00006 + 1 :
                                             wire_qout_00046_00006
                                             ;

            I1db4ea6916125702e7fb09d0f742e60a  <=  wire_qout_00046_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I38d78b447217271a63f30f78b424e2ae     <=
                                             wire_qout_00046_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00007 + 1 :
                                             wire_qout_00046_00007
                                             ;

            Idc445d3f5b3b62562b0ac83e5f17e92a  <=  wire_qout_00046_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4c8d7e5474b19a7c63444d0cb6143728     <=
                                             wire_qout_00046_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00008 + 1 :
                                             wire_qout_00046_00008
                                             ;

            Iee6e52d75c093a24eb4e5e0b45feb256  <=  wire_qout_00046_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia4bc4b7414bf31305ec8f63e7eda61e7     <=
                                             wire_qout_00046_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00009 + 1 :
                                             wire_qout_00046_00009
                                             ;

            Id48fe0672aa98f987162931527e9f9bc  <=  wire_qout_00046_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibbebe287d56c7d627f3ffcf706575e77     <=
                                             wire_qout_00046_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00010 + 1 :
                                             wire_qout_00046_00010
                                             ;

            Idce46f6d03376bea1ba361e8c59f8bd1  <=  wire_qout_00046_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I83867e6ee369fff7e39ef5c8d5398fef     <=
                                             wire_qout_00046_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00011 + 1 :
                                             wire_qout_00046_00011
                                             ;

            Ie79ce8adeef2c3c24a3386f054d0cf5b  <=  wire_qout_00046_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1d40df7dbf99674f987bd06db714a702     <=
                                             wire_qout_00046_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00012 + 1 :
                                             wire_qout_00046_00012
                                             ;

            I0d41bef808860bde56d48792764612d5  <=  wire_qout_00046_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I92f42789cb81760ff2973e3a5fe915c3     <=
                                             wire_qout_00046_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00013 + 1 :
                                             wire_qout_00046_00013
                                             ;

            Ib6ae81df8db1dae269437861ee11ec0d  <=  wire_qout_00046_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idbd5f2a25ab05808721cf9c403017565     <=
                                             wire_qout_00046_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00014 + 1 :
                                             wire_qout_00046_00014
                                             ;

            I33ddee677715877c11a1df45cbfb01ac  <=  wire_qout_00046_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7ca5f07d6d3c2a045dfd55ae5214dd65     <=
                                             wire_qout_00046_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00046_00015 + 1 :
                                             wire_qout_00046_00015
                                             ;

            I433dd5092cf1851cd196feade3cfa6d8  <=  wire_qout_00046_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7f4e1445c68abbadce23944b99d206f9     <=
                                             wire_qout_00047_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00000 + 1 :
                                             wire_qout_00047_00000
                                             ;

            I71d3a999d88e591e102398409b3adebf  <=  wire_qout_00047_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id9f28016678e5e2127d9f0aa93e0b534     <=
                                             wire_qout_00047_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00001 + 1 :
                                             wire_qout_00047_00001
                                             ;

            Iebecd2d19f9174d87deedc1a273e7baa  <=  wire_qout_00047_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6b939c57a8b7c7c51ab43e1b1df12f6a     <=
                                             wire_qout_00047_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00002 + 1 :
                                             wire_qout_00047_00002
                                             ;

            I168afc1863f909dbcb6a9230db9f3e00  <=  wire_qout_00047_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic5d0df586d56bf4cb322d4c3ad677385     <=
                                             wire_qout_00047_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00003 + 1 :
                                             wire_qout_00047_00003
                                             ;

            I1c4b29e48d0effac4839037ae5688334  <=  wire_qout_00047_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2e287724873cf6761799eaf464ed6302     <=
                                             wire_qout_00047_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00004 + 1 :
                                             wire_qout_00047_00004
                                             ;

            I431fc2e9533012c8571d8158d4777dea  <=  wire_qout_00047_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia7a10cffe31a53aafa1104b97543280b     <=
                                             wire_qout_00047_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00005 + 1 :
                                             wire_qout_00047_00005
                                             ;

            Ief72606c77113ae37845e4aa4a2ae5e7  <=  wire_qout_00047_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ieeb089c6a18791a2227c8571913d689a     <=
                                             wire_qout_00047_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00006 + 1 :
                                             wire_qout_00047_00006
                                             ;

            I641539560711ff1824bd90baa0f21f96  <=  wire_qout_00047_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib29b00328971c3cd67209a5ea5b63b0a     <=
                                             wire_qout_00047_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00007 + 1 :
                                             wire_qout_00047_00007
                                             ;

            I3ac0799861144b599995318bdade2114  <=  wire_qout_00047_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I517e0868f2bb9a22c287a1f3eeaad2f3     <=
                                             wire_qout_00047_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00008 + 1 :
                                             wire_qout_00047_00008
                                             ;

            Ie83fa8157a7cce44c2e25f46ce897dbb  <=  wire_qout_00047_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2bc9f76469e2a3f9846560ad1975cf54     <=
                                             wire_qout_00047_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00009 + 1 :
                                             wire_qout_00047_00009
                                             ;

            I8be4711146486fea913843e497065b50  <=  wire_qout_00047_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9f089315e435cd69d2929fdd936a8a77     <=
                                             wire_qout_00047_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00010 + 1 :
                                             wire_qout_00047_00010
                                             ;

            I65171c9ee8449407484e5c82d13c6751  <=  wire_qout_00047_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9b54c9fb4179423c731217286e329930     <=
                                             wire_qout_00047_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00011 + 1 :
                                             wire_qout_00047_00011
                                             ;

            I7353ebf3a1cde89d2bb3fa667f7f5485  <=  wire_qout_00047_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I82fb41ab743146badfd2e82258afb310     <=
                                             wire_qout_00047_00012[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00012 + 1 :
                                             wire_qout_00047_00012
                                             ;

            I669d34b955d2991ebbb31c149ad1b6f8  <=  wire_qout_00047_00012[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5619b91de99eead78befdcba1c62411e     <=
                                             wire_qout_00047_00013[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00013 + 1 :
                                             wire_qout_00047_00013
                                             ;

            Iabb01dc9980b4879a7356712b51df0d6  <=  wire_qout_00047_00013[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I83dd2047dece99cd841b2e7955819d57     <=
                                             wire_qout_00047_00014[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00014 + 1 :
                                             wire_qout_00047_00014
                                             ;

            I373841aa2bcbad8232d54ac9035a3ef9  <=  wire_qout_00047_00014[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8c927e66ccbf4d19f07af5ef9fbfe3fb     <=
                                             wire_qout_00047_00015[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00047_00015 + 1 :
                                             wire_qout_00047_00015
                                             ;

            Ib6124faff821158c6a2c9a9c454ab68c  <=  wire_qout_00047_00015[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0793fa8938acdf65486e5582d01b9e5a     <=
                                             wire_qout_00048_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00048_00000 + 1 :
                                             wire_qout_00048_00000
                                             ;

            I6f7a45fe64ffeda9ed120be3a4519aea  <=  wire_qout_00048_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ied68d7ba0ee9974eb33767e737760b4d     <=
                                             wire_qout_00048_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00048_00001 + 1 :
                                             wire_qout_00048_00001
                                             ;

            Id1dafb7e45b860d506e0c2c91b28142e  <=  wire_qout_00048_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I95ba37056659b29fd4318a68d85445e8     <=
                                             wire_qout_00048_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00048_00002 + 1 :
                                             wire_qout_00048_00002
                                             ;

            I5f1609647f1e71cef4ba2d605c6c8445  <=  wire_qout_00048_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I08d7051a18f358d08728f1c401c15c47     <=
                                             wire_qout_00048_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00048_00003 + 1 :
                                             wire_qout_00048_00003
                                             ;

            If17c0096ce34b88007247bf4c429d5c4  <=  wire_qout_00048_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I768b6f55827ac49eb6ac2655e9397be1     <=
                                             wire_qout_00048_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00048_00004 + 1 :
                                             wire_qout_00048_00004
                                             ;

            Ifc2963762403a00c4f3662b2863c991e  <=  wire_qout_00048_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic66f737fe60c55d4c10e5d72b307a061     <=
                                             wire_qout_00048_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00048_00005 + 1 :
                                             wire_qout_00048_00005
                                             ;

            I5fdd8e1550feaecd81b82069fe73ed7e  <=  wire_qout_00048_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5653779f15c6c9b0f3b26927c48d6234     <=
                                             wire_qout_00048_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00048_00006 + 1 :
                                             wire_qout_00048_00006
                                             ;

            I85654bd3a07b4329aba17d8b27777f4e  <=  wire_qout_00048_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iac550729fc437fd67151fab57134ec88     <=
                                             wire_qout_00048_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00048_00007 + 1 :
                                             wire_qout_00048_00007
                                             ;

            Ibf2a253afde05c905d0b2404c5a808a0  <=  wire_qout_00048_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I853b03c5826eedc3c67a2fae7a640212     <=
                                             wire_qout_00048_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00048_00008 + 1 :
                                             wire_qout_00048_00008
                                             ;

            I3ade5535a79ce83857481ac771cd8618  <=  wire_qout_00048_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If46a6b47c1c52243cc0bc92d1edb594f     <=
                                             wire_qout_00049_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00049_00000 + 1 :
                                             wire_qout_00049_00000
                                             ;

            I221524a69e18854f029cad30e8f94e8a  <=  wire_qout_00049_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I75b36a9b429cd657afc8151b9613aca6     <=
                                             wire_qout_00049_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00049_00001 + 1 :
                                             wire_qout_00049_00001
                                             ;

            Ied764ee7730ad129b6f62837ef50774a  <=  wire_qout_00049_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ife682dd9f677da4d27294fb61b141948     <=
                                             wire_qout_00049_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00049_00002 + 1 :
                                             wire_qout_00049_00002
                                             ;

            Ic98f33c6a4613534bcc9b6bc4b4f2d17  <=  wire_qout_00049_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic2b6177a9c586b274b68b25584e6df2c     <=
                                             wire_qout_00049_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00049_00003 + 1 :
                                             wire_qout_00049_00003
                                             ;

            I92eb6f60c14ee9eecb01718b01ea980f  <=  wire_qout_00049_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0d23011c4381496a19cced7bf7960546     <=
                                             wire_qout_00049_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00049_00004 + 1 :
                                             wire_qout_00049_00004
                                             ;

            I97e82e5f6775d1e31537b891597223bd  <=  wire_qout_00049_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic5992d5eaeafd5dded641a7d9801e763     <=
                                             wire_qout_00049_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00049_00005 + 1 :
                                             wire_qout_00049_00005
                                             ;

            Iba1c0ebd9cefeb0dd7f690bdbbbfec58  <=  wire_qout_00049_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic9e7fe68b9045c6c9eb86185b5f5872e     <=
                                             wire_qout_00049_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00049_00006 + 1 :
                                             wire_qout_00049_00006
                                             ;

            I235c3a9fd3e8ea1cee762c10bc8e2c53  <=  wire_qout_00049_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I51ad746720b5e6e09ab50f0283552f1a     <=
                                             wire_qout_00049_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00049_00007 + 1 :
                                             wire_qout_00049_00007
                                             ;

            Idd474d80b50992537d6f527faf279800  <=  wire_qout_00049_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0c8964888a1315507f5d71959dd24cf0     <=
                                             wire_qout_00049_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00049_00008 + 1 :
                                             wire_qout_00049_00008
                                             ;

            I88a89b2d938552458dab9bc34728959b  <=  wire_qout_00049_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id4d4f814a0bb3418cbf70c306acf048f     <=
                                             wire_qout_00050_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00050_00000 + 1 :
                                             wire_qout_00050_00000
                                             ;

            Ib105151d91678f81978495ff94b1e651  <=  wire_qout_00050_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic91bd7b4bd148e526ca21d4a5ba87be9     <=
                                             wire_qout_00050_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00050_00001 + 1 :
                                             wire_qout_00050_00001
                                             ;

            I4edd64d1f1da865b1eb886e22726a033  <=  wire_qout_00050_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7959dddc32f0f181b3ba39149afe1016     <=
                                             wire_qout_00050_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00050_00002 + 1 :
                                             wire_qout_00050_00002
                                             ;

            Ia7c9c24f8e993526e76c6915e56908c4  <=  wire_qout_00050_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I087263600b5f38be072a4f1db787aea7     <=
                                             wire_qout_00050_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00050_00003 + 1 :
                                             wire_qout_00050_00003
                                             ;

            Ib0dadebad37d9ea9d01350054872863c  <=  wire_qout_00050_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I78d17a56de5cbe08191ef23b9731c485     <=
                                             wire_qout_00050_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00050_00004 + 1 :
                                             wire_qout_00050_00004
                                             ;

            I76fd9005abd511c3c5bf6c77de8bf2f3  <=  wire_qout_00050_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I82f713a43596df3b935d6da6f8041dc2     <=
                                             wire_qout_00050_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00050_00005 + 1 :
                                             wire_qout_00050_00005
                                             ;

            Ic124975d36a292816146a2fe61ab3ab9  <=  wire_qout_00050_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I422987396853a6a39dabb6e7ddbf91fb     <=
                                             wire_qout_00050_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00050_00006 + 1 :
                                             wire_qout_00050_00006
                                             ;

            I70a4926e9e6a05fa9ee51a26988862fe  <=  wire_qout_00050_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibb6556671e104141dd33188ea5fc024d     <=
                                             wire_qout_00050_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00050_00007 + 1 :
                                             wire_qout_00050_00007
                                             ;

            Idc5e98f6958786ccf95d39b922b42ea9  <=  wire_qout_00050_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie42ce76076a2a5e887e0112086012da6     <=
                                             wire_qout_00050_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00050_00008 + 1 :
                                             wire_qout_00050_00008
                                             ;

            I8879df010bbdf6e5fc9370e2fb3289b4  <=  wire_qout_00050_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4aea430599b9c0702b3bebd5960b5c91     <=
                                             wire_qout_00051_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00051_00000 + 1 :
                                             wire_qout_00051_00000
                                             ;

            I94a9de743d5bedbea3876de954f479bd  <=  wire_qout_00051_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icbe11a3970136e485eee1bc5053e7273     <=
                                             wire_qout_00051_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00051_00001 + 1 :
                                             wire_qout_00051_00001
                                             ;

            I17c9d8f658dd6b2916b645d103f4702a  <=  wire_qout_00051_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0a7f1ea1719c1f5ff104445a4130a5a8     <=
                                             wire_qout_00051_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00051_00002 + 1 :
                                             wire_qout_00051_00002
                                             ;

            I384e50fa8daa639124f083dda56fac00  <=  wire_qout_00051_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1802d759f26dd919bc315bfd4156238d     <=
                                             wire_qout_00051_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00051_00003 + 1 :
                                             wire_qout_00051_00003
                                             ;

            Ie165d0729542c81ca89f45d15e0afd3d  <=  wire_qout_00051_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2148493e253783fad70f4f2807b83008     <=
                                             wire_qout_00051_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00051_00004 + 1 :
                                             wire_qout_00051_00004
                                             ;

            Ie8e29053f122a9247b0dec291c6ef4f3  <=  wire_qout_00051_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I39e7f78d33aa7f50264908d2efe23634     <=
                                             wire_qout_00051_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00051_00005 + 1 :
                                             wire_qout_00051_00005
                                             ;

            I453dd7d7c0a2f003f0b67e909630d641  <=  wire_qout_00051_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I844be5874def16af98de935019f35fe8     <=
                                             wire_qout_00051_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00051_00006 + 1 :
                                             wire_qout_00051_00006
                                             ;

            I5707d30ca29842b6a96cfaeb44ac6668  <=  wire_qout_00051_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iee5172ba70a6e368b4903f9ff1d93471     <=
                                             wire_qout_00051_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00051_00007 + 1 :
                                             wire_qout_00051_00007
                                             ;

            I3fbd40faa4c3b78b547b8348c466fd1f  <=  wire_qout_00051_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1f34b473283291e0970879465c005e2f     <=
                                             wire_qout_00051_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00051_00008 + 1 :
                                             wire_qout_00051_00008
                                             ;

            I9a403c511fe2d44472ab319a9477199c  <=  wire_qout_00051_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie1e0b5120737a7f4bf845618ccd22239     <=
                                             wire_qout_00052_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00000 + 1 :
                                             wire_qout_00052_00000
                                             ;

            I9db50007841762c9a10f6b7e9d40f858  <=  wire_qout_00052_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8abec3020ee5358f8768e5595e9992b4     <=
                                             wire_qout_00052_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00001 + 1 :
                                             wire_qout_00052_00001
                                             ;

            I89c5af1a6176cefa1f77ee69996473cb  <=  wire_qout_00052_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6fe683073211a484cb6e3c416b365d9f     <=
                                             wire_qout_00052_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00002 + 1 :
                                             wire_qout_00052_00002
                                             ;

            I5ede62333e0f7ddc5446b653ba9a2382  <=  wire_qout_00052_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id7d764da58ade36853e8a45b5ee19dc3     <=
                                             wire_qout_00052_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00003 + 1 :
                                             wire_qout_00052_00003
                                             ;

            I69d82ab774d52c219509e993e7cc4deb  <=  wire_qout_00052_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3cee2fdf353643deac7d6bca20c8fb52     <=
                                             wire_qout_00052_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00004 + 1 :
                                             wire_qout_00052_00004
                                             ;

            I0eaa22f5eca8f33dd254fe241017a098  <=  wire_qout_00052_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie9b8f8f0434fe3783c3d8f68fef30e50     <=
                                             wire_qout_00052_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00005 + 1 :
                                             wire_qout_00052_00005
                                             ;

            I570c036d0237c53bb069c52d621e539e  <=  wire_qout_00052_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I68cba8ad7742cbb34d0b1fb16be4a58a     <=
                                             wire_qout_00052_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00006 + 1 :
                                             wire_qout_00052_00006
                                             ;

            I9d7614d286377329eb3999213889b707  <=  wire_qout_00052_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idcea56657d40e0fdf9a1c2d920938fd6     <=
                                             wire_qout_00052_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00007 + 1 :
                                             wire_qout_00052_00007
                                             ;

            I3eab1582cc42db0ac7739386cce2a712  <=  wire_qout_00052_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic549ffab8f0ce161a177faa2ffd1326d     <=
                                             wire_qout_00052_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00008 + 1 :
                                             wire_qout_00052_00008
                                             ;

            Ie4827dc0983c1a63053c08de6e36d375  <=  wire_qout_00052_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4d463d500f93f74b2724972ec1d62439     <=
                                             wire_qout_00052_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00009 + 1 :
                                             wire_qout_00052_00009
                                             ;

            I2eed3d32a27d51036e17c4a21382b4c1  <=  wire_qout_00052_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iba2f362e263953331649c726afa9c481     <=
                                             wire_qout_00052_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00010 + 1 :
                                             wire_qout_00052_00010
                                             ;

            Ie039ab562e9cf90289047b5425186123  <=  wire_qout_00052_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6a053d931fb030e03d4882856d3bda75     <=
                                             wire_qout_00052_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00052_00011 + 1 :
                                             wire_qout_00052_00011
                                             ;

            Iefbdf686d9452a62cb99cf023a4d9fe7  <=  wire_qout_00052_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I27ede93004e0c240efaa56cc8c570910     <=
                                             wire_qout_00053_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00000 + 1 :
                                             wire_qout_00053_00000
                                             ;

            Idc5dd6caa4ed17a63746d30d381a944e  <=  wire_qout_00053_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I61a11c1711ca10eefea3438722b40bff     <=
                                             wire_qout_00053_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00001 + 1 :
                                             wire_qout_00053_00001
                                             ;

            I17086dc5193aa55e5c6f56ecd365cc00  <=  wire_qout_00053_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia7924c88692cfddf24fb1eff66eacb7e     <=
                                             wire_qout_00053_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00002 + 1 :
                                             wire_qout_00053_00002
                                             ;

            Ib2fe0f68044c11f879e512a200f8099e  <=  wire_qout_00053_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibcfd01e622f7f5a5156dd9b335b4e5e0     <=
                                             wire_qout_00053_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00003 + 1 :
                                             wire_qout_00053_00003
                                             ;

            I768720af835b02a8dab376ef23d17a15  <=  wire_qout_00053_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7f6f418ea51b4298da8758bda3f6a21b     <=
                                             wire_qout_00053_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00004 + 1 :
                                             wire_qout_00053_00004
                                             ;

            I1d98943b01a6a2d8c4db18b98dd62f5c  <=  wire_qout_00053_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7185da8937449e23abdd0f39a4b3ed7d     <=
                                             wire_qout_00053_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00005 + 1 :
                                             wire_qout_00053_00005
                                             ;

            Id3b089fb6edd5bcfdbca142fddd5ff89  <=  wire_qout_00053_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idc3e3ffa31d9b76c7cf9358a5b2e65d7     <=
                                             wire_qout_00053_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00006 + 1 :
                                             wire_qout_00053_00006
                                             ;

            I5196382b75d16892d550f17893de15ec  <=  wire_qout_00053_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I31fe8c887c4aff7c69336676cd31aaa1     <=
                                             wire_qout_00053_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00007 + 1 :
                                             wire_qout_00053_00007
                                             ;

            I6387919f2426c283e2d70e471cda54a6  <=  wire_qout_00053_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I59684d5fe6bbb4b54ac097bd25fceef5     <=
                                             wire_qout_00053_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00008 + 1 :
                                             wire_qout_00053_00008
                                             ;

            I3b84dad6d0dd8730312b3e20c6d5a2a8  <=  wire_qout_00053_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I86a7cd69148f9590ce91d0aa270d6c54     <=
                                             wire_qout_00053_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00009 + 1 :
                                             wire_qout_00053_00009
                                             ;

            I2a4bbedf880a9a7b4e1bf946f9f96c0e  <=  wire_qout_00053_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iabce1ccdd968980f622f0e137b159d11     <=
                                             wire_qout_00053_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00010 + 1 :
                                             wire_qout_00053_00010
                                             ;

            I49d35ec6369de10afb15be8e0cf135c3  <=  wire_qout_00053_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iff02977d7b4c733cca1794246f630931     <=
                                             wire_qout_00053_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00053_00011 + 1 :
                                             wire_qout_00053_00011
                                             ;

            Ic3ba4531855366e9a060cec1c7694844  <=  wire_qout_00053_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9026c904e5ead7ff2994c4f781d61466     <=
                                             wire_qout_00054_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00000 + 1 :
                                             wire_qout_00054_00000
                                             ;

            I4dbabfd592b74aef93b819163130ef5e  <=  wire_qout_00054_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I99d7489ba87c629c6dd9702a9bbfd3c8     <=
                                             wire_qout_00054_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00001 + 1 :
                                             wire_qout_00054_00001
                                             ;

            I9ece87047aec25abc02a5eea72f0e647  <=  wire_qout_00054_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifaf191e0d00ba6da7019c2efcf08e1d9     <=
                                             wire_qout_00054_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00002 + 1 :
                                             wire_qout_00054_00002
                                             ;

            I3ed6426fbdba8aaf1c948cca7442b3a6  <=  wire_qout_00054_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4c295991fb08c90862a2f3ba6489000a     <=
                                             wire_qout_00054_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00003 + 1 :
                                             wire_qout_00054_00003
                                             ;

            I24075f37c6bbd90c83370de1a2e58af2  <=  wire_qout_00054_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iee61d179da125934298400256788cbb8     <=
                                             wire_qout_00054_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00004 + 1 :
                                             wire_qout_00054_00004
                                             ;

            I3175159add7b814df637c2db8feb43f6  <=  wire_qout_00054_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If87c84440426fb24070372dc1d4bf315     <=
                                             wire_qout_00054_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00005 + 1 :
                                             wire_qout_00054_00005
                                             ;

            I0a569f6536789efb7ad2377c11842830  <=  wire_qout_00054_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib9259a807b31c1b7a528d336bfc403ee     <=
                                             wire_qout_00054_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00006 + 1 :
                                             wire_qout_00054_00006
                                             ;

            Iae6ed7748692f2edf1aa9d73380075f0  <=  wire_qout_00054_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I411c4d909b2a571e685cd703245516d7     <=
                                             wire_qout_00054_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00007 + 1 :
                                             wire_qout_00054_00007
                                             ;

            Ib4ae1cedd09d72c235765a6cd7e91366  <=  wire_qout_00054_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If8425453cca8fc8623cb85375c4b8a1d     <=
                                             wire_qout_00054_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00008 + 1 :
                                             wire_qout_00054_00008
                                             ;

            Ie2d946edaddd3c87f328e861f3e72c0a  <=  wire_qout_00054_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I654b497f62df75fa283127b5de29b1ad     <=
                                             wire_qout_00054_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00009 + 1 :
                                             wire_qout_00054_00009
                                             ;

            Id6b508145cd21ba088ab8fda34577c35  <=  wire_qout_00054_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2768519342f7b8a1ee40c1d5ac502b66     <=
                                             wire_qout_00054_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00010 + 1 :
                                             wire_qout_00054_00010
                                             ;

            Ifa6e3541f5e12bf9677ffc51d0392749  <=  wire_qout_00054_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8e354c1c5ba44fe5430887248ce0c43b     <=
                                             wire_qout_00054_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00054_00011 + 1 :
                                             wire_qout_00054_00011
                                             ;

            I21e72a7e5870151c3247d15121e5fb4f  <=  wire_qout_00054_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8970d8a8aea29913e8696c14c153d16e     <=
                                             wire_qout_00055_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00000 + 1 :
                                             wire_qout_00055_00000
                                             ;

            Iba283e99a57d0a3b78ad2e309c316b65  <=  wire_qout_00055_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3555c6e2fd480a6be11549bf95a9b0b1     <=
                                             wire_qout_00055_00001[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00001 + 1 :
                                             wire_qout_00055_00001
                                             ;

            Ifba3e46933049cb093d2c1809f3a8a3e  <=  wire_qout_00055_00001[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8d5600a352e8ba4756f917f912fda6dd     <=
                                             wire_qout_00055_00002[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00002 + 1 :
                                             wire_qout_00055_00002
                                             ;

            I4af3e2bf2ebc913ac902b48da672c5b6  <=  wire_qout_00055_00002[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7e99d73c95e7ae5c3fe07a3c60ef52eb     <=
                                             wire_qout_00055_00003[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00003 + 1 :
                                             wire_qout_00055_00003
                                             ;

            Ifbadefd3a7ab50719a703400ddd742c6  <=  wire_qout_00055_00003[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I831633aebe5c6a52b98d630205376f3a     <=
                                             wire_qout_00055_00004[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00004 + 1 :
                                             wire_qout_00055_00004
                                             ;

            If2042aede3390bd208a281f0380c95a4  <=  wire_qout_00055_00004[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I82e35482de74223be0d2558334ac2dfb     <=
                                             wire_qout_00055_00005[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00005 + 1 :
                                             wire_qout_00055_00005
                                             ;

            I19b73c5c93a71e90f620572f23f0e6d2  <=  wire_qout_00055_00005[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iae2a6f9649ef1bb193e4f0ab5ecbc3e3     <=
                                             wire_qout_00055_00006[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00006 + 1 :
                                             wire_qout_00055_00006
                                             ;

            I4b99891bed4f5c149cd4a5b4f1dde0f0  <=  wire_qout_00055_00006[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie8eca65d791ad2f6e8f4ed244f22ae3d     <=
                                             wire_qout_00055_00007[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00007 + 1 :
                                             wire_qout_00055_00007
                                             ;

            I3472ee8c06644490252e606b62bf9bd5  <=  wire_qout_00055_00007[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic24146b01094df9b9ccd455a791f239d     <=
                                             wire_qout_00055_00008[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00008 + 1 :
                                             wire_qout_00055_00008
                                             ;

            Idb1efe99b5d7fd567a7f82cfd52f7eb8  <=  wire_qout_00055_00008[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1c9031fd54ff9417d44c9fb17dc1fc63     <=
                                             wire_qout_00055_00009[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00009 + 1 :
                                             wire_qout_00055_00009
                                             ;

            I24f82a3f2c0e8df486fe495dd95cf8bc  <=  wire_qout_00055_00009[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idefa20487bc5ba6daff03e6b327d76c6     <=
                                             wire_qout_00055_00010[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00010 + 1 :
                                             wire_qout_00055_00010
                                             ;

            I83ecf12f3b38fc14c3b75e47b71ecc09  <=  wire_qout_00055_00010[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6f984fd9ea27b40ab3afeac8afd29ade     <=
                                             wire_qout_00055_00011[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00055_00011 + 1 :
                                             wire_qout_00055_00011
                                             ;

            I74cbc0ec3bb682e0f927890eef8d7a58  <=  wire_qout_00055_00011[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0be92debced4961df5f461fe81e80bf1     <=
                                             wire_qout_00056_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00056_00000 + 1 :
                                             wire_qout_00056_00000
                                             ;

            I989dda9add29306d7b3c0f376822763a  <=  wire_qout_00056_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia7bdaba4c6601b7146498aea6c9a3e07     <=
                                             wire_qout_00057_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00057_00000 + 1 :
                                             wire_qout_00057_00000
                                             ;

            Ibc929201e2eeb3e61cc8f0acbade497a  <=  wire_qout_00057_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id450c0a1cabe087be051fbf4158e6016     <=
                                             wire_qout_00058_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00058_00000 + 1 :
                                             wire_qout_00058_00000
                                             ;

            Ib0dfbbbca2d3d264065f73b4241caed5  <=  wire_qout_00058_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I656d0d69f6e243746b87ad67764dbc3d     <=
                                             wire_qout_00059_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00059_00000 + 1 :
                                             wire_qout_00059_00000
                                             ;

            I339786aa60d4c71d12c65db27ac420fe  <=  wire_qout_00059_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iab9d870dc1ad159bbaecb20a9b72f005     <=
                                             wire_qout_00060_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00060_00000 + 1 :
                                             wire_qout_00060_00000
                                             ;

            I3ade020bbdf8f954821f737439513043  <=  wire_qout_00060_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id53b60854f19e095c38f2c255dc57f29     <=
                                             wire_qout_00061_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00061_00000 + 1 :
                                             wire_qout_00061_00000
                                             ;

            Ia50526cd3a3174bebc5a7a0889fda661  <=  wire_qout_00061_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If9ba44a2e4a8f0b61692fc69ebeb82bd     <=
                                             wire_qout_00062_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00062_00000 + 1 :
                                             wire_qout_00062_00000
                                             ;

            Ie9f37dba0791359bc426a73639ce33ad  <=  wire_qout_00062_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ief95e8620a1c8ddfd6df673a3a223bd8     <=
                                             wire_qout_00063_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00063_00000 + 1 :
                                             wire_qout_00063_00000
                                             ;

            I9518532a8617fc8290eb6a5e981dea94  <=  wire_qout_00063_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I61519bc0aa02ed461dbb91851d0ae19e     <=
                                             wire_qout_00064_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00064_00000 + 1 :
                                             wire_qout_00064_00000
                                             ;

            If66524125bfde5aa48ac70c4e448b38f  <=  wire_qout_00064_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie0c11d584811174a66ca221baf87c36b     <=
                                             wire_qout_00065_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00065_00000 + 1 :
                                             wire_qout_00065_00000
                                             ;

            Ic3ec6375998b05a3e48f6c5fe7b3910b  <=  wire_qout_00065_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If10f4f45ff0fd17541735934ad20f187     <=
                                             wire_qout_00066_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00066_00000 + 1 :
                                             wire_qout_00066_00000
                                             ;

            I0ac421af6e311b6005c3e02e93ff94ce  <=  wire_qout_00066_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I445919f07a6fa8654211301a9a6126bd     <=
                                             wire_qout_00067_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00067_00000 + 1 :
                                             wire_qout_00067_00000
                                             ;

            Ib9db80f43718305a8a8774d8d80c86c9  <=  wire_qout_00067_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I64102b82893352549abd2e2132b19476     <=
                                             wire_qout_00068_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00068_00000 + 1 :
                                             wire_qout_00068_00000
                                             ;

            I3b775b06b5d78fcd7373c966a62f44ad  <=  wire_qout_00068_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1fc1933fe891ac26f35a42a1b242d919     <=
                                             wire_qout_00069_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00069_00000 + 1 :
                                             wire_qout_00069_00000
                                             ;

            If2372a5956f21f97eeb9c76281b6675e  <=  wire_qout_00069_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I84dfba8bcf8ad3b85f9472fd60d607b5     <=
                                             wire_qout_00070_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00070_00000 + 1 :
                                             wire_qout_00070_00000
                                             ;

            I7b32c2b108e24750e2a24785668af3ea  <=  wire_qout_00070_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4302fccefe5ee13161f9ad49f9ddf43c     <=
                                             wire_qout_00071_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00071_00000 + 1 :
                                             wire_qout_00071_00000
                                             ;

            I8ec99197a7d823f5745d382c10161430  <=  wire_qout_00071_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I59d7153724d3b3805af799692fbe245a     <=
                                             wire_qout_00072_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00072_00000 + 1 :
                                             wire_qout_00072_00000
                                             ;

            Ib895fec0b3756932b85962c1d129a03e  <=  wire_qout_00072_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id1650d0e39be078027493f58e9bbcbdd     <=
                                             wire_qout_00073_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00073_00000 + 1 :
                                             wire_qout_00073_00000
                                             ;

            I76aab345d13c6678fe37a4a7133cfd7d  <=  wire_qout_00073_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If40ad4aca8dbb3bf7dde8c2ff2e5b8f2     <=
                                             wire_qout_00074_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00074_00000 + 1 :
                                             wire_qout_00074_00000
                                             ;

            Ib4f368fa3d3ec11d9ffb2ae9a2ae6310  <=  wire_qout_00074_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie49f173549396caeab1d13da36e37c65     <=
                                             wire_qout_00075_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00075_00000 + 1 :
                                             wire_qout_00075_00000
                                             ;

            Idd0f3cfc5599481c954a2bfe69f044e5  <=  wire_qout_00075_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3002a0e0cdf8e79bc7186a876410d106     <=
                                             wire_qout_00076_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00076_00000 + 1 :
                                             wire_qout_00076_00000
                                             ;

            Ie624c4dad5036a25ca314b94cf3c4b95  <=  wire_qout_00076_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2b50fa03f584d10e9af3be085a02a12c     <=
                                             wire_qout_00077_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00077_00000 + 1 :
                                             wire_qout_00077_00000
                                             ;

            Ibf4b3caa5655cfb6663f9b7e2383bbbf  <=  wire_qout_00077_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If473d172a7bff5aeae99245bbb72978d     <=
                                             wire_qout_00078_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00078_00000 + 1 :
                                             wire_qout_00078_00000
                                             ;

            I049d1c09c15def12ba7bae95fc1c3d55  <=  wire_qout_00078_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib89f7b5625995290a64bcfb143d978ca     <=
                                             wire_qout_00079_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00079_00000 + 1 :
                                             wire_qout_00079_00000
                                             ;

            Ide06ba186ddb179b489ba6e3e209e3e8  <=  wire_qout_00079_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iebe0c9b4a87d58a1c55e2ee6b01603c4     <=
                                             wire_qout_00080_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00080_00000 + 1 :
                                             wire_qout_00080_00000
                                             ;

            I1b78785ebe2e7f77a3125a6334c4dc54  <=  wire_qout_00080_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I104411bb641d2445c7e1385a809bb682     <=
                                             wire_qout_00081_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00081_00000 + 1 :
                                             wire_qout_00081_00000
                                             ;

            Ie79c93f1703121713fb9401617f349a8  <=  wire_qout_00081_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I47dd28b4ae4f7151aff5bb271e35b716     <=
                                             wire_qout_00082_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00082_00000 + 1 :
                                             wire_qout_00082_00000
                                             ;

            Icf25f076eec2bf81c899c66f6cfbebc0  <=  wire_qout_00082_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3a27d5573b748df459b90a5a347f9d09     <=
                                             wire_qout_00083_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00083_00000 + 1 :
                                             wire_qout_00083_00000
                                             ;

            Ic5c837a0556d1cb66edbf0294d08283a  <=  wire_qout_00083_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2dbef85d2b2b95af39c3a98c4e143253     <=
                                             wire_qout_00084_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00084_00000 + 1 :
                                             wire_qout_00084_00000
                                             ;

            I51ff4bda38746682e3cd4c68118c3216  <=  wire_qout_00084_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I510d39830ae7b0a857ac11baa7c144d3     <=
                                             wire_qout_00085_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00085_00000 + 1 :
                                             wire_qout_00085_00000
                                             ;

            I1c074a53e6c0f2467bcdd7c952f51670  <=  wire_qout_00085_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2751a94a66ea4cb44c512df4c509937f     <=
                                             wire_qout_00086_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00086_00000 + 1 :
                                             wire_qout_00086_00000
                                             ;

            I37c49c5a2af240496f5a5706b0d42ea6  <=  wire_qout_00086_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic9a003bfb70ac2da6c229fcad09246d4     <=
                                             wire_qout_00087_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00087_00000 + 1 :
                                             wire_qout_00087_00000
                                             ;

            Ia94c439131e1df5c95fc8ad3cfdba473  <=  wire_qout_00087_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I34ed986182a3311a8cb005b3dccc224b     <=
                                             wire_qout_00088_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00088_00000 + 1 :
                                             wire_qout_00088_00000
                                             ;

            I723a6fee3b2496f23c48b3584f8bf9ce  <=  wire_qout_00088_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic79281755397f6099ff30c5d07d7e6de     <=
                                             wire_qout_00089_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00089_00000 + 1 :
                                             wire_qout_00089_00000
                                             ;

            I648b62fa0bc2185c1756ee531e8e34de  <=  wire_qout_00089_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8d6559ccc33cbc663584923a55b928b5     <=
                                             wire_qout_00090_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00090_00000 + 1 :
                                             wire_qout_00090_00000
                                             ;

            Ife631f9a3c4c64a3d92aa9586ae75f3c  <=  wire_qout_00090_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4f0a4c241844e390318f11899a0f2c5a     <=
                                             wire_qout_00091_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00091_00000 + 1 :
                                             wire_qout_00091_00000
                                             ;

            Iaac1d82f0846fce1bd88ebf8e60300ac  <=  wire_qout_00091_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I45fffa266ce3838f82d755b59216a4d6     <=
                                             wire_qout_00092_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00092_00000 + 1 :
                                             wire_qout_00092_00000
                                             ;

            I48cd09f035f668536cd288a23010b07b  <=  wire_qout_00092_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8f0e65f5db47d5460d4ec2172807a3e1     <=
                                             wire_qout_00093_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00093_00000 + 1 :
                                             wire_qout_00093_00000
                                             ;

            I119b2e5c2fea5338244c4019884af26f  <=  wire_qout_00093_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I34127c0d1af2438e13b6f4709ece80ba     <=
                                             wire_qout_00094_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00094_00000 + 1 :
                                             wire_qout_00094_00000
                                             ;

            I2bd34b2fd12f12bc301fd0d5d69c0fb6  <=  wire_qout_00094_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3a67de0e76bbf29d8c77c21865abda2f     <=
                                             wire_qout_00095_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00095_00000 + 1 :
                                             wire_qout_00095_00000
                                             ;

            Ib715b1e0061b84ce614a30d961a83e7e  <=  wire_qout_00095_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic64e64aeb754249b868e14311ea19759     <=
                                             wire_qout_00096_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00096_00000 + 1 :
                                             wire_qout_00096_00000
                                             ;

            Ief8c2838abac83370fd7ec25c06d509b  <=  wire_qout_00096_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic4aa0dc9014c8445f8d9a7723d7263f5     <=
                                             wire_qout_00097_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00097_00000 + 1 :
                                             wire_qout_00097_00000
                                             ;

            I561d79eb079915c0b1732cbddb119c2d  <=  wire_qout_00097_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I47b988d017580bdfe8f443904b1f3aac     <=
                                             wire_qout_00098_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00098_00000 + 1 :
                                             wire_qout_00098_00000
                                             ;

            I8bb75bf828d5ef337fa6a965808e4638  <=  wire_qout_00098_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ica9ff13e8c3850be6c70b0b06c1d9fbf     <=
                                             wire_qout_00099_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00099_00000 + 1 :
                                             wire_qout_00099_00000
                                             ;

            I11ba339c8250d07b497c88a39a6df1ac  <=  wire_qout_00099_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If2efeb489911f295dd7722cb22ea521d     <=
                                             wire_qout_00100_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00100_00000 + 1 :
                                             wire_qout_00100_00000
                                             ;

            I173aa69cf52114e223ac1410d90b4bfe  <=  wire_qout_00100_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iaa16dffcc01e41e6ff17e92bdefe3df5     <=
                                             wire_qout_00101_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00101_00000 + 1 :
                                             wire_qout_00101_00000
                                             ;

            Ia4e89e99acb95f4183474b94798ca35d  <=  wire_qout_00101_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie8857b9841fbd795a4192976ef7ecc25     <=
                                             wire_qout_00102_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00102_00000 + 1 :
                                             wire_qout_00102_00000
                                             ;

            If4c36727ab1c29bf78f72e8acfc00d7c  <=  wire_qout_00102_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If12aef69eea28052aa3bdb6ac31af205     <=
                                             wire_qout_00103_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00103_00000 + 1 :
                                             wire_qout_00103_00000
                                             ;

            I6426943b4ab66f17c2b7b399ccc7a6a9  <=  wire_qout_00103_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0b3c6162ae2b9221738a18a29489887f     <=
                                             wire_qout_00104_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00104_00000 + 1 :
                                             wire_qout_00104_00000
                                             ;

            Iddcffa815489773b3688fd68dba18bd8  <=  wire_qout_00104_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I08211bba29e87faf4079152bcc973e7d     <=
                                             wire_qout_00105_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00105_00000 + 1 :
                                             wire_qout_00105_00000
                                             ;

            Id00642563679fa9a6696f8e7bbdf6576  <=  wire_qout_00105_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibff3da265f1c3f21548f5b019e1a9dc1     <=
                                             wire_qout_00106_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00106_00000 + 1 :
                                             wire_qout_00106_00000
                                             ;

            Ifda1c55899cd3506853cc82b450b3936  <=  wire_qout_00106_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie9fa1762d7844b0d781afdfb0771cea9     <=
                                             wire_qout_00107_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00107_00000 + 1 :
                                             wire_qout_00107_00000
                                             ;

            Ib5d1a7cdbcba0b654c12063d4f1768e1  <=  wire_qout_00107_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia677d504b9f7fc2698c0345f236428ba     <=
                                             wire_qout_00108_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00108_00000 + 1 :
                                             wire_qout_00108_00000
                                             ;

            I5e8ed024e2f2548bb375a2ecf1918a5f  <=  wire_qout_00108_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idebce29121c0481df83d755b60ff632c     <=
                                             wire_qout_00109_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00109_00000 + 1 :
                                             wire_qout_00109_00000
                                             ;

            Id25deba967318f049de8163e67262f4b  <=  wire_qout_00109_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iad2c780a6386674d50cca54d8c4ebd86     <=
                                             wire_qout_00110_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00110_00000 + 1 :
                                             wire_qout_00110_00000
                                             ;

            I925f6b549a25cdc8f85152eb21ea3b58  <=  wire_qout_00110_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If1d7944e7c4828ddb91ffea28609cbc7     <=
                                             wire_qout_00111_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00111_00000 + 1 :
                                             wire_qout_00111_00000
                                             ;

            I9b49e1acb81ef5b088b808d2e4ce9954  <=  wire_qout_00111_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I843a68ceb0adab829091f31d0de56eb6     <=
                                             wire_qout_00112_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00112_00000 + 1 :
                                             wire_qout_00112_00000
                                             ;

            I6386a4dd26e7c36165dc265b3a2c93cf  <=  wire_qout_00112_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I59701b9eb54dda2744a79cebe7d73f3b     <=
                                             wire_qout_00113_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00113_00000 + 1 :
                                             wire_qout_00113_00000
                                             ;

            Ia20709f08cfff3a51d4af1e81d640400  <=  wire_qout_00113_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If63cf5e8f47e4e51176401f0d954ea23     <=
                                             wire_qout_00114_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00114_00000 + 1 :
                                             wire_qout_00114_00000
                                             ;

            I1ff042bdb52aac5d69791e96e2f9706c  <=  wire_qout_00114_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id09454844b525697de3e3727d89551e4     <=
                                             wire_qout_00115_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00115_00000 + 1 :
                                             wire_qout_00115_00000
                                             ;

            Iaa2cbf59f6f61198b4fcf5a741cd5bc8  <=  wire_qout_00115_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6d1b2ce4368945b56eee7814638471cc     <=
                                             wire_qout_00116_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00116_00000 + 1 :
                                             wire_qout_00116_00000
                                             ;

            I01c94743a11042e75638ba6618356203  <=  wire_qout_00116_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6079945faa57335b1c902ccf7f960a70     <=
                                             wire_qout_00117_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00117_00000 + 1 :
                                             wire_qout_00117_00000
                                             ;

            I0a0340a0e52145f3597accfe4a4e8624  <=  wire_qout_00117_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie7752906ac55cf51f3e96e8c0046f1aa     <=
                                             wire_qout_00118_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00118_00000 + 1 :
                                             wire_qout_00118_00000
                                             ;

            I3bb4d24caaa0882a75125e466070f0b1  <=  wire_qout_00118_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2d7d4135a94f5df949283c043228791f     <=
                                             wire_qout_00119_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00119_00000 + 1 :
                                             wire_qout_00119_00000
                                             ;

            I44ead0ab5ccc53226fccc03024643771  <=  wire_qout_00119_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I99c75e3d26c5d01f6ae9abcd05407d8c     <=
                                             wire_qout_00120_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00120_00000 + 1 :
                                             wire_qout_00120_00000
                                             ;

            Iaded125f7fd5c833e7206dd7071069be  <=  wire_qout_00120_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I81e6f97621dbfb2fed6fc236005a2b19     <=
                                             wire_qout_00121_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00121_00000 + 1 :
                                             wire_qout_00121_00000
                                             ;

            I373be7c3f9511a2906584e33e5048abf  <=  wire_qout_00121_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ieac60532dcfc916a65054e35cf31d6d2     <=
                                             wire_qout_00122_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00122_00000 + 1 :
                                             wire_qout_00122_00000
                                             ;

            Ie0b5f51835ebdb508a596eeebf0e4847  <=  wire_qout_00122_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ib7eb83ba73e0dc17f69c357b6ca555bf     <=
                                             wire_qout_00123_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00123_00000 + 1 :
                                             wire_qout_00123_00000
                                             ;

            Iddb75e0197b9a76b36a59ac2a7ccdf3a  <=  wire_qout_00123_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5139d8a7a099e3c619c60647c15b7420     <=
                                             wire_qout_00124_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00124_00000 + 1 :
                                             wire_qout_00124_00000
                                             ;

            I08c03198b9599b2f4590e3022e398f7c  <=  wire_qout_00124_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6ccd2e11ebd5b2de80b120e20650a602     <=
                                             wire_qout_00125_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00125_00000 + 1 :
                                             wire_qout_00125_00000
                                             ;

            Ia4f3cff223e24815ee1d86bf41756f06  <=  wire_qout_00125_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie669cebe5fe39e1a841f8dd3c1f6bc57     <=
                                             wire_qout_00126_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00126_00000 + 1 :
                                             wire_qout_00126_00000
                                             ;

            I56592e1452c4b559af19465b30230ec0  <=  wire_qout_00126_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If32acb9fc212c4af34099acf6df2bc5a     <=
                                             wire_qout_00127_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00127_00000 + 1 :
                                             wire_qout_00127_00000
                                             ;

            I213ce488e5345fa405a9c5df297d6f74  <=  wire_qout_00127_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I075ce236a181bf925c8ccce91d9bc8cd     <=
                                             wire_qout_00128_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00128_00000 + 1 :
                                             wire_qout_00128_00000
                                             ;

            Iefac1e428116a797c2c0803410ac5601  <=  wire_qout_00128_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I541d4e422b999a0dfca44d275178e1d9     <=
                                             wire_qout_00129_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00129_00000 + 1 :
                                             wire_qout_00129_00000
                                             ;

            I8b419d5827e5b1af9649d602401c189a  <=  wire_qout_00129_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I3e02657f3d9f79338cd083ed024bf96c     <=
                                             wire_qout_00130_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00130_00000 + 1 :
                                             wire_qout_00130_00000
                                             ;

            Ie989550c9101de382056dd60d5da0e01  <=  wire_qout_00130_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia5e5537405ab8edcc7cd43c86837d43d     <=
                                             wire_qout_00131_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00131_00000 + 1 :
                                             wire_qout_00131_00000
                                             ;

            I259010e323e1e8dcd9dd719091131f6c  <=  wire_qout_00131_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I07ff388e3b6c7288f0f6c35a345023fe     <=
                                             wire_qout_00132_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00132_00000 + 1 :
                                             wire_qout_00132_00000
                                             ;

            I389ac86954fd70464c9550e3fed4ed33  <=  wire_qout_00132_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I56cb3b3e193ca5068734417fd0ec4e02     <=
                                             wire_qout_00133_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00133_00000 + 1 :
                                             wire_qout_00133_00000
                                             ;

            I77371f0e55b4684d1af196ed52d3d997  <=  wire_qout_00133_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I5bbf1765d8f81581d0cf31c0bc755fb3     <=
                                             wire_qout_00134_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00134_00000 + 1 :
                                             wire_qout_00134_00000
                                             ;

            I5a21996f5724a2a49fcf8e928c01b062  <=  wire_qout_00134_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iaa1643095e518846cdede4d5a90dff84     <=
                                             wire_qout_00135_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00135_00000 + 1 :
                                             wire_qout_00135_00000
                                             ;

            Id46108963921efa50aff64d4dd7d1701  <=  wire_qout_00135_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iee6e12f4717a3279dd31b874eabae69e     <=
                                             wire_qout_00136_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00136_00000 + 1 :
                                             wire_qout_00136_00000
                                             ;

            I8da50e5093acefb6f809aed64564a53e  <=  wire_qout_00136_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic52a9edbbc5283844d2514ea142ca6e2     <=
                                             wire_qout_00137_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00137_00000 + 1 :
                                             wire_qout_00137_00000
                                             ;

            I03b0694777d0160a83cbc82ac1397736  <=  wire_qout_00137_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ice3e978c8da2a7de5b28542a5589f0a2     <=
                                             wire_qout_00138_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00138_00000 + 1 :
                                             wire_qout_00138_00000
                                             ;

            I85c2bffb93569d9fe1b1bcb10b98bcac  <=  wire_qout_00138_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I336a425aed221c85ca80b9a97d21d6b1     <=
                                             wire_qout_00139_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00139_00000 + 1 :
                                             wire_qout_00139_00000
                                             ;

            Id00274c88b93867a80606343add1cdab  <=  wire_qout_00139_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie477c0f3b77bb299ba8b1a410d211ef7     <=
                                             wire_qout_00140_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00140_00000 + 1 :
                                             wire_qout_00140_00000
                                             ;

            I61e829cbf7d6c0ef8ddc11677981e2cf  <=  wire_qout_00140_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie62920d089ae762603cd33fbf97d92bb     <=
                                             wire_qout_00141_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00141_00000 + 1 :
                                             wire_qout_00141_00000
                                             ;

            I9e8ae2aed048068b01b3bd46f30baae8  <=  wire_qout_00141_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2ca952e4e676537fd5a8fc71ecfa10e9     <=
                                             wire_qout_00142_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00142_00000 + 1 :
                                             wire_qout_00142_00000
                                             ;

            I7dab71adbe62687846fc027d2789451d  <=  wire_qout_00142_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iefd31e7ff3c829c88f60bc89d70afcf7     <=
                                             wire_qout_00143_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00143_00000 + 1 :
                                             wire_qout_00143_00000
                                             ;

            If1295608bd218ed60922a0b95bf1d098  <=  wire_qout_00143_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iafa987a413fd8fcacfe872bc0f5bc2d6     <=
                                             wire_qout_00144_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00144_00000 + 1 :
                                             wire_qout_00144_00000
                                             ;

            Idf04e08c120ed116af14a62659675b44  <=  wire_qout_00144_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I305c1ea420d666f258e38c5a65847367     <=
                                             wire_qout_00145_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00145_00000 + 1 :
                                             wire_qout_00145_00000
                                             ;

            Ieb7614ad1b1bfed3e2b0089a72fe214a  <=  wire_qout_00145_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9f040c4088bfab72d74e5332e9710d1a     <=
                                             wire_qout_00146_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00146_00000 + 1 :
                                             wire_qout_00146_00000
                                             ;

            I589062eca318b25dfe5735da455b6fe1  <=  wire_qout_00146_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia2f41f9778324a06daeb185c736516a4     <=
                                             wire_qout_00147_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00147_00000 + 1 :
                                             wire_qout_00147_00000
                                             ;

            If3db87afb3ea184c9e4020c5e45cb161  <=  wire_qout_00147_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id9778ba5fbdbed4d33a092da6b68c414     <=
                                             wire_qout_00148_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00148_00000 + 1 :
                                             wire_qout_00148_00000
                                             ;

            Ia14bc1fcd5bbdcb60b8e68298f7d716a  <=  wire_qout_00148_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I27c2c79d0d719c71c8e28218d1174a13     <=
                                             wire_qout_00149_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00149_00000 + 1 :
                                             wire_qout_00149_00000
                                             ;

            I268b60cb371b3d46dc3f8b0009f541b1  <=  wire_qout_00149_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2a9d6a774769b12ae20bc0cee0c36f5c     <=
                                             wire_qout_00150_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00150_00000 + 1 :
                                             wire_qout_00150_00000
                                             ;

            If2cd93b57cd1c2b91ee7a73a97dd19f2  <=  wire_qout_00150_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I2c567b75f1399c069b95284f4c36b6d1     <=
                                             wire_qout_00151_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00151_00000 + 1 :
                                             wire_qout_00151_00000
                                             ;

            Id81305359a07db527e49fda05cd2784f  <=  wire_qout_00151_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If3d3eb609abfd6e315eec803d2e94490     <=
                                             wire_qout_00152_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00152_00000 + 1 :
                                             wire_qout_00152_00000
                                             ;

            Id8292eca087c1a17dc8b5a572a76f21f  <=  wire_qout_00152_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9c58aea7ce986b1d28f5808b347c015d     <=
                                             wire_qout_00153_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00153_00000 + 1 :
                                             wire_qout_00153_00000
                                             ;

            Iddb19725b093506e5e521d8d68dcb8e1  <=  wire_qout_00153_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Id139c7a783196941100003b6cb0cd1e7     <=
                                             wire_qout_00154_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00154_00000 + 1 :
                                             wire_qout_00154_00000
                                             ;

            I0b573d3a86a3111451da661e46384876  <=  wire_qout_00154_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I524d7614b01460778da3ce98f6aaa3d9     <=
                                             wire_qout_00155_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00155_00000 + 1 :
                                             wire_qout_00155_00000
                                             ;

            I0ff479e61d1a0cede88ebffb073c60be  <=  wire_qout_00155_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8acda65f116d5c91cbe2662ac282aa31     <=
                                             wire_qout_00156_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00156_00000 + 1 :
                                             wire_qout_00156_00000
                                             ;

            Icd6f8f5df6b4ca4c81855e974db76526  <=  wire_qout_00156_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If67dbe22f8d22b3430215fb0deae8204     <=
                                             wire_qout_00157_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00157_00000 + 1 :
                                             wire_qout_00157_00000
                                             ;

            I7ce064a756dad56d37684d5d7d168047  <=  wire_qout_00157_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9a35cd7512787263abedd6d9913cf507     <=
                                             wire_qout_00158_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00158_00000 + 1 :
                                             wire_qout_00158_00000
                                             ;

            Ied2ea62cfb21602645babc36e27b8218  <=  wire_qout_00158_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If9cca23469c5e6001650f1f8b1360ae8     <=
                                             wire_qout_00159_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00159_00000 + 1 :
                                             wire_qout_00159_00000
                                             ;

            I79b85da6e5ce0b02ebd1619115c98e24  <=  wire_qout_00159_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icc2606ae8f9a3b425225ae7339112b9d     <=
                                             wire_qout_00160_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00160_00000 + 1 :
                                             wire_qout_00160_00000
                                             ;

            I8e1ddd7e4185c28caa71d30bc28138f3  <=  wire_qout_00160_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I34aa1802d24e074ae54563898929abfa     <=
                                             wire_qout_00161_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00161_00000 + 1 :
                                             wire_qout_00161_00000
                                             ;

            Iab0bff1633e2f3ea0bfbc291f3ab5d29  <=  wire_qout_00161_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Icb85b3464dc40e8504c53c377e889c45     <=
                                             wire_qout_00162_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00162_00000 + 1 :
                                             wire_qout_00162_00000
                                             ;

            I5f0751fceaa008feba5c6867ced453dc  <=  wire_qout_00162_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie595a7d10b5ac84c0301fb55bebd3680     <=
                                             wire_qout_00163_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00163_00000 + 1 :
                                             wire_qout_00163_00000
                                             ;

            I9f6751c15237c20b0cf2175575195ea7  <=  wire_qout_00163_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9c217a672cabc05efbdff218637123ba     <=
                                             wire_qout_00164_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00164_00000 + 1 :
                                             wire_qout_00164_00000
                                             ;

            I6ea50be10bc990a1206cdc9e28e0c4c2  <=  wire_qout_00164_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If20f3780b4af857ffe8083056085517a     <=
                                             wire_qout_00165_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00165_00000 + 1 :
                                             wire_qout_00165_00000
                                             ;

            I43c2fab87f70ea883321ab82de85f133  <=  wire_qout_00165_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic2e275bfa8ab3d2002d2aa374ac9bfe2     <=
                                             wire_qout_00166_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00166_00000 + 1 :
                                             wire_qout_00166_00000
                                             ;

            I1af02ed6cf00d4cb0704b5e44c83bfa3  <=  wire_qout_00166_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Iac5798fd9915b6778700da6a14f6a381     <=
                                             wire_qout_00167_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00167_00000 + 1 :
                                             wire_qout_00167_00000
                                             ;

            Ib71611afdd0381cc1884f5ddbbae1acc  <=  wire_qout_00167_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ide3204bf317fdfb993410d338085b174     <=
                                             wire_qout_00168_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00168_00000 + 1 :
                                             wire_qout_00168_00000
                                             ;

            I38fc49afce0298846ae8ed63ae715e81  <=  wire_qout_00168_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ic3a95140fc1029efa17a6557bc977719     <=
                                             wire_qout_00169_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00169_00000 + 1 :
                                             wire_qout_00169_00000
                                             ;

            Iddc3e44d83e8253e5129b6cbf5082df7  <=  wire_qout_00169_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I647d3a46bb2c7ed0f1ec08760b3858be     <=
                                             wire_qout_00170_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00170_00000 + 1 :
                                             wire_qout_00170_00000
                                             ;

            I975a87bdda30c5b6be8d2f0e4b107450  <=  wire_qout_00170_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4816747af9d9fc8dc85fd831336ec710     <=
                                             wire_qout_00171_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00171_00000 + 1 :
                                             wire_qout_00171_00000
                                             ;

            I582bd96afa764ded148202f738b7a1df  <=  wire_qout_00171_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1f66c026a5437320bd1f4df2ff71663d     <=
                                             wire_qout_00172_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00172_00000 + 1 :
                                             wire_qout_00172_00000
                                             ;

            I6fb88d97bc9ed37a06b729020a1df140  <=  wire_qout_00172_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If347c58c328193f420286ea27a4afa20     <=
                                             wire_qout_00173_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00173_00000 + 1 :
                                             wire_qout_00173_00000
                                             ;

            I1500943c4a550e78fc169437b0a663b7  <=  wire_qout_00173_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I7a126c8304be920f2a920315dc61ba7f     <=
                                             wire_qout_00174_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00174_00000 + 1 :
                                             wire_qout_00174_00000
                                             ;

            I0b83f4ef8ba9badb27e81b32765ec5b6  <=  wire_qout_00174_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I237327d6a74df1fb05537dc3691ebf11     <=
                                             wire_qout_00175_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00175_00000 + 1 :
                                             wire_qout_00175_00000
                                             ;

            I2c420acf428e44cdd9ca9998e276f258  <=  wire_qout_00175_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I64a3e8bb4c87b066806d33a5306a2c53     <=
                                             wire_qout_00176_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00176_00000 + 1 :
                                             wire_qout_00176_00000
                                             ;

            Ic7b6dae3017b55dd3cd27423d5f1b0ec  <=  wire_qout_00176_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ibbca6ec39234473fb517447a8beacafc     <=
                                             wire_qout_00177_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00177_00000 + 1 :
                                             wire_qout_00177_00000
                                             ;

            I4a91a7c9b2a0f3552b8f2ef4e2398be2  <=  wire_qout_00177_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I78327356176a16fc996188b83b058cbc     <=
                                             wire_qout_00178_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00178_00000 + 1 :
                                             wire_qout_00178_00000
                                             ;

            I99ff29c7ba68b5d0819f1e1bead51287  <=  wire_qout_00178_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifec496c87a7a2474855067305ac8cba3     <=
                                             wire_qout_00179_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00179_00000 + 1 :
                                             wire_qout_00179_00000
                                             ;

            If06b00be0356a2be5074d958ddcdb2f9  <=  wire_qout_00179_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I41584165a62caaa37ddebbf79bb8b617     <=
                                             wire_qout_00180_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00180_00000 + 1 :
                                             wire_qout_00180_00000
                                             ;

            I604283449f13c7b225ea03f99f2e296a  <=  wire_qout_00180_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Idf0916d6b025aad6eccb98ada5ba3aca     <=
                                             wire_qout_00181_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00181_00000 + 1 :
                                             wire_qout_00181_00000
                                             ;

            I2b600e5f5c146ee97c4044c08e1f5ad5  <=  wire_qout_00181_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I00ef133d5a53f8f99f35b50327e5272b     <=
                                             wire_qout_00182_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00182_00000 + 1 :
                                             wire_qout_00182_00000
                                             ;

            I9fe16403fc21bb1159a5e0305fd1ef69  <=  wire_qout_00182_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I6f0e302d38d75982d0761e306ce9f146     <=
                                             wire_qout_00183_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00183_00000 + 1 :
                                             wire_qout_00183_00000
                                             ;

            Iabdb9374e5caee281c25b003624b2c4e  <=  wire_qout_00183_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I127eed5de00e10a020717e796de76c7d     <=
                                             wire_qout_00184_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00184_00000 + 1 :
                                             wire_qout_00184_00000
                                             ;

            Ibd12036702fe60b57354b3aac921559d  <=  wire_qout_00184_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If9aad73aefb1b225f35e8c813b85fe87     <=
                                             wire_qout_00185_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00185_00000 + 1 :
                                             wire_qout_00185_00000
                                             ;

            Ib1639811de6eb1c38257800c201fb704  <=  wire_qout_00185_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I00a89ac37676521a081a21b1ec1a0798     <=
                                             wire_qout_00186_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00186_00000 + 1 :
                                             wire_qout_00186_00000
                                             ;

            If926d98f659e8fe4bbf36ad2c5c852c5  <=  wire_qout_00186_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I06f3a34f2b1770ef82ddc2a732b3d4fb     <=
                                             wire_qout_00187_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00187_00000 + 1 :
                                             wire_qout_00187_00000
                                             ;

            I211f8d7f97ebb8eb3e50313513abfb1b  <=  wire_qout_00187_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I4744d64a746f16004e3bedaaa41465f1     <=
                                             wire_qout_00188_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00188_00000 + 1 :
                                             wire_qout_00188_00000
                                             ;

            I304ac9f96945546cdf1b6f1fa7136731  <=  wire_qout_00188_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ifae0cc6cc1c65d24bbe84c4ba938e2ea     <=
                                             wire_qout_00189_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00189_00000 + 1 :
                                             wire_qout_00189_00000
                                             ;

            I7a9800418bd5c195fc47a72370680b56  <=  wire_qout_00189_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1223c21129382d41e4f38ef4bbe60c2f     <=
                                             wire_qout_00190_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00190_00000 + 1 :
                                             wire_qout_00190_00000
                                             ;

            I5f6a61c9f0c67510e148e596f553a4d6  <=  wire_qout_00190_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I14e36e16df00adcd7dc1973d3852d2d9     <=
                                             wire_qout_00191_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00191_00000 + 1 :
                                             wire_qout_00191_00000
                                             ;

            I8e313ceb21359bcc44114ab217b1c394  <=  wire_qout_00191_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0d05ae27b53fb6939e4c2f862a8d20b2     <=
                                             wire_qout_00192_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00192_00000 + 1 :
                                             wire_qout_00192_00000
                                             ;

            I4c9518755c33d725221ad79ee6badba9  <=  wire_qout_00192_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I97a6fcc08929c3b7d15e36d7706ed13d     <=
                                             wire_qout_00193_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00193_00000 + 1 :
                                             wire_qout_00193_00000
                                             ;

            I3c3cffec9f47c9979cb9503f222f370c  <=  wire_qout_00193_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I1f04e86bf27596718836d0a09adbe120     <=
                                             wire_qout_00194_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00194_00000 + 1 :
                                             wire_qout_00194_00000
                                             ;

            I68d6769541fdc3df321e192f645c667f  <=  wire_qout_00194_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie40873cfd6d10a61a94a761becf588a8     <=
                                             wire_qout_00195_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00195_00000 + 1 :
                                             wire_qout_00195_00000
                                             ;

            Ided55428cbb77f454c2607ac783d7548  <=  wire_qout_00195_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I61960ed74fee948cc12bd1fd8384559a     <=
                                             wire_qout_00196_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00196_00000 + 1 :
                                             wire_qout_00196_00000
                                             ;

            Ifd3d4f3e2a388b3c70e7704d6351e0ba  <=  wire_qout_00196_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I8533a3ec4be4c49166184c94761eaebc     <=
                                             wire_qout_00197_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00197_00000 + 1 :
                                             wire_qout_00197_00000
                                             ;

            I17d32f292758416fe02527dfd938fa0d  <=  wire_qout_00197_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I00be319b5bdb85ffaf3bb0eca0b348b6     <=
                                             wire_qout_00198_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00198_00000 + 1 :
                                             wire_qout_00198_00000
                                             ;

            I9ce3942aba354c1fd7d6b9a39c994d7b  <=  wire_qout_00198_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ie889c916b5af185b52ff5e2e3cc23045     <=
                                             wire_qout_00199_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00199_00000 + 1 :
                                             wire_qout_00199_00000
                                             ;

            I2c6c6041c9c69c84f4d64af6458955f5  <=  wire_qout_00199_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I89697be6dcb2e7f972db498c1b1dea71     <=
                                             wire_qout_00200_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00200_00000 + 1 :
                                             wire_qout_00200_00000
                                             ;

            I830a4fffe1244e071eb82c28ddc4a308  <=  wire_qout_00200_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If13dfbfff7cd8e197bb44006a3db73bf     <=
                                             wire_qout_00201_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00201_00000 + 1 :
                                             wire_qout_00201_00000
                                             ;

            Ifad8e46fc3844bbfaf434a14f6b5869d  <=  wire_qout_00201_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I87ed6c3e172c7a06bf6aefe7bf718d70     <=
                                             wire_qout_00202_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00202_00000 + 1 :
                                             wire_qout_00202_00000
                                             ;

            I10a6c6a8fdb0003de1f360c148777d0f  <=  wire_qout_00202_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I0db87adc849839fab3a4c9884d5a4882     <=
                                             wire_qout_00203_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00203_00000 + 1 :
                                             wire_qout_00203_00000
                                             ;

            I4cde586fc28f8d03fc9934d56f7ff7b8  <=  wire_qout_00203_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I535e01a6c35fd7b455e4b79b1d4bb414     <=
                                             wire_qout_00204_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00204_00000 + 1 :
                                             wire_qout_00204_00000
                                             ;

            Ib83a067fb08e118dcf794902beef9405  <=  wire_qout_00204_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            Ia2d1c752cc4b405adb97a815e90a7b96     <=
                                             wire_qout_00205_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00205_00000 + 1 :
                                             wire_qout_00205_00000
                                             ;

            I358cf9609272a4562423a85f9b2f56bf  <=  wire_qout_00205_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            I9ac12eb3878f6fc7dc428fe5e7f35d97     <=
                                             wire_qout_00206_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00206_00000 + 1 :
                                             wire_qout_00206_00000
                                             ;

            Ic1e9d9113150ad57954c0e369259dc62  <=  wire_qout_00206_00000[SGN_MAX_SUM_WDTH] ;

           end
           if (start_d2) begin
            If46fa11dfadb0691eaaa0a40836e08d8     <=
                                             wire_qout_00207_00000[SGN_MAX_SUM_WDTH] ?
                                             ~wire_qout_00207_00000 + 1 :
                                             wire_qout_00207_00000
                                             ;

            If7fe3f5ccbb5b279e41fd183c8ff3974  <=  wire_qout_00207_00000[SGN_MAX_SUM_WDTH] ;

           end
       end

   end

assign wire_qout_00000_00000      = sum0_00000 +  ~Iea07d1adf9016a29cffd61d183e268d0 +1;
assign wire_qout_00000_00001      = sum0_00000 +  ~If92db65b39a83e1c699e4cc6d7f9e57b +1;
assign wire_qout_00000_00002      = sum0_00000 +  ~I8f2986bc015fcc64ac5e5395ac6dd851 +1;
assign wire_qout_00000_00003      = sum0_00000 +  ~I355725a804e0df68b4acf96ca98f2448 +1;
assign wire_qout_00000_00004      = sum0_00000 +  ~I78212ae965ab2dcb2eed0b060d6b253f +1;
assign wire_qout_00000_00005      = sum0_00000 +  ~I0b56aa7a1b7549c91dddd3a06ecbaacf +1;
assign wire_qout_00000_00006      = sum0_00000 +  ~I71412803cc5229025487255aec62ec4f +1;
assign wire_qout_00000_00007      = sum0_00000 +  ~I32fcb28a27356bc6f403528836ea4c1f +1;
assign wire_qout_00000_00008      = sum0_00000 +  ~Iad354d876cb9fc72fc0143e6f7da9357 +1;
assign wire_qout_00000_00009      = sum0_00000 +  ~If6e745bb85abba7282dae1f6f701225e +1;
assign wire_qout_00000_00010      = sum0_00000 +  ~I93bb43c1b89d4c70a57bdc019d64fd22 +1;
assign wire_qout_00000_00011      = sum0_00000 +  ~I7a2e554d07bbea291f2cfc18694fca3a +1;
assign wire_qout_00000_00012      = sum0_00000 +  ~I3e59b2419c7dd1553b792d536208514e +1;
assign wire_qout_00000_00013      = sum0_00000 +  ~I46894c6526983bf1ce4b503159131b41 +1;
assign wire_qout_00000_00014      = sum0_00000 +  ~I6404d0df952b5bf8292c753e4c6f35d8 +1;
assign wire_qout_00000_00015      = sum0_00000 +  ~I8522c402e654d007abffcb0e904af5e6 +1;
assign wire_qout_00000_00016      = sum0_00000 +  ~I5ed85845c39337c37791f16e718069b4 +1;
assign wire_qout_00000_00017      = sum0_00000 +  ~I89013d61c1ea8da8b1c6071cc21c316f +1;
assign wire_qout_00000_00018      = sum0_00000 +  ~I4102100fa5f1dd299af0190862efcc42 +1;
assign wire_qout_00000_00019      = sum0_00000 +  ~I4939f69abb1eac56d5021e06406a93b5 +1;
assign wire_qout_00000_00020      = sum0_00000 +  ~Iadbd245bf842aebb456417579a3e6296 +1;
assign wire_qout_00000_00021      = sum0_00000 +  ~Ifc8ece44a4e68c3117eda9e65f3084d2 +1;
assign wire_qout_00001_00000      = sum0_00001 +  ~I91679dfab57a372eddc7f9b94a231edb +1;
assign wire_qout_00001_00001      = sum0_00001 +  ~I2213c1a2b831f421707a261f5a58b1b1 +1;
assign wire_qout_00001_00002      = sum0_00001 +  ~Ic53b875b2ddcba11406eb2ca39354757 +1;
assign wire_qout_00001_00003      = sum0_00001 +  ~I634484f00590216c0f74f975c9c83400 +1;
assign wire_qout_00001_00004      = sum0_00001 +  ~Ib3b1db2d8b669988c887ed780e439b26 +1;
assign wire_qout_00001_00005      = sum0_00001 +  ~I735db8b0ee0ec98e4cce0030b11508da +1;
assign wire_qout_00001_00006      = sum0_00001 +  ~If1607e907e626902ee26d15020a64c21 +1;
assign wire_qout_00001_00007      = sum0_00001 +  ~I081b38dbb37d4c14a6a9fd3fefa13daa +1;
assign wire_qout_00001_00008      = sum0_00001 +  ~Ibac5e7b6d4bf5cd6926358318f0c418f +1;
assign wire_qout_00001_00009      = sum0_00001 +  ~Iadfc60386481092ae85cc148a2c40abb +1;
assign wire_qout_00001_00010      = sum0_00001 +  ~Ie0ee5445c56a5f9b41640b57422206de +1;
assign wire_qout_00001_00011      = sum0_00001 +  ~Ie5f8620371236cb11c9e88c16b509ee8 +1;
assign wire_qout_00001_00012      = sum0_00001 +  ~I8d7c1fe2e33bbd45379b0325a3c5e989 +1;
assign wire_qout_00001_00013      = sum0_00001 +  ~I4fbdc4ee57a3be42b62d9bd43078d6ef +1;
assign wire_qout_00001_00014      = sum0_00001 +  ~I5510b88bfd65811b3200adf4ef975b48 +1;
assign wire_qout_00001_00015      = sum0_00001 +  ~Ib57ef2f577cca54713c16717cbbd1ce9 +1;
assign wire_qout_00001_00016      = sum0_00001 +  ~I15943aa74e9fbbaebdc0d54eb6a3bffa +1;
assign wire_qout_00001_00017      = sum0_00001 +  ~I6ac24c46319a787daa5c545de8c6eeea +1;
assign wire_qout_00001_00018      = sum0_00001 +  ~I52403a0454e5fa002e79eaab7ea497bd +1;
assign wire_qout_00001_00019      = sum0_00001 +  ~I634f0ce28934600a1a31ab0d8e59b4a9 +1;
assign wire_qout_00001_00020      = sum0_00001 +  ~I7103aa739616a39c03e675ea0efb0335 +1;
assign wire_qout_00001_00021      = sum0_00001 +  ~I0296d01fd3f9a269a617efd4beea9b8b +1;
assign wire_qout_00002_00000      = sum0_00002 +  ~I065a81ba25962785215583e7ece27661 +1;
assign wire_qout_00002_00001      = sum0_00002 +  ~I631a3300cb6685f47da7781940ec5d27 +1;
assign wire_qout_00002_00002      = sum0_00002 +  ~I8bbe1a2ace8f51aa22cca5d9fc66f136 +1;
assign wire_qout_00002_00003      = sum0_00002 +  ~I38c3e3e136acb79c8a0ff850bcc55f16 +1;
assign wire_qout_00002_00004      = sum0_00002 +  ~I35b2c7e9cdc53a98913e1c16a3a47b37 +1;
assign wire_qout_00002_00005      = sum0_00002 +  ~Ib1a2b31d49ae476e2f1fb9acba2d5af0 +1;
assign wire_qout_00002_00006      = sum0_00002 +  ~Ic72f41f9bbf470aee3c9b9b8787b31c3 +1;
assign wire_qout_00002_00007      = sum0_00002 +  ~I3ea4c33a9419820ed54460eb64134dff +1;
assign wire_qout_00002_00008      = sum0_00002 +  ~Ia0d940e16c8cbd4f7544f5a5cd7d83b2 +1;
assign wire_qout_00002_00009      = sum0_00002 +  ~I4a8abfa0896ce414d9b98093ef84455f +1;
assign wire_qout_00002_00010      = sum0_00002 +  ~I680be647bf2a62e0ee9b5d379dc87b4f +1;
assign wire_qout_00002_00011      = sum0_00002 +  ~If4d75f83299a21802b6fbe136913489f +1;
assign wire_qout_00002_00012      = sum0_00002 +  ~Ibddfda6413e3dd2f483c3174ea836b6a +1;
assign wire_qout_00002_00013      = sum0_00002 +  ~I33bddb0adcc2af7b12a83bf843036385 +1;
assign wire_qout_00002_00014      = sum0_00002 +  ~I529f92b82248efe2cf64f7da0ec8283c +1;
assign wire_qout_00002_00015      = sum0_00002 +  ~I2f34af0036985cd94ade9cc905bec065 +1;
assign wire_qout_00002_00016      = sum0_00002 +  ~Ia1a0d8d7dfd6e877f15cce773f85f5b7 +1;
assign wire_qout_00002_00017      = sum0_00002 +  ~I5dd29fd1a73df5662d2b636e7285bad9 +1;
assign wire_qout_00002_00018      = sum0_00002 +  ~Ide530e6f4622c8a7b101b6dce9650e42 +1;
assign wire_qout_00002_00019      = sum0_00002 +  ~Ibaf00a6780325882067a79f0c4d693d2 +1;
assign wire_qout_00002_00020      = sum0_00002 +  ~I16e3559c63ebfed83d6698fc9a9cd93a +1;
assign wire_qout_00002_00021      = sum0_00002 +  ~I9747a02384abb1c2dd1f52b3a5a999cc +1;
assign wire_qout_00003_00000      = sum0_00003 +  ~Iceb7a1d4c23806b8f5824016779ad129 +1;
assign wire_qout_00003_00001      = sum0_00003 +  ~I40ef50004a60ae58aedc49eb5e6797c9 +1;
assign wire_qout_00003_00002      = sum0_00003 +  ~I753f92da60980736440aba814a156f1e +1;
assign wire_qout_00003_00003      = sum0_00003 +  ~I4ac79b67a8904b95f7912d24af420585 +1;
assign wire_qout_00003_00004      = sum0_00003 +  ~Iad44c932cfa5c249c5e59f8c706173a8 +1;
assign wire_qout_00003_00005      = sum0_00003 +  ~I10f14b6433498e3b9e9bf021b60115e8 +1;
assign wire_qout_00003_00006      = sum0_00003 +  ~I96008f47b9f134c9c4274cfcfb28e550 +1;
assign wire_qout_00003_00007      = sum0_00003 +  ~Id0344146d1a53d418add6d2b185377dd +1;
assign wire_qout_00003_00008      = sum0_00003 +  ~I1eede74f12d37331b399eb7136bc621f +1;
assign wire_qout_00003_00009      = sum0_00003 +  ~I3e4754acc31d99bc71525789bdee0c1a +1;
assign wire_qout_00003_00010      = sum0_00003 +  ~I11c1fc94a3bd6dffa17e1571cc6ae97c +1;
assign wire_qout_00003_00011      = sum0_00003 +  ~I5395ee57418c31e11cf847f0f514ec19 +1;
assign wire_qout_00003_00012      = sum0_00003 +  ~Iff125392fa39afebae1637a19c4e23ec +1;
assign wire_qout_00003_00013      = sum0_00003 +  ~Ia6308e16fae5428f4ab6560f5b21479a +1;
assign wire_qout_00003_00014      = sum0_00003 +  ~I5ea02b5349cd4d99ccbcb6b26f0cfdd7 +1;
assign wire_qout_00003_00015      = sum0_00003 +  ~I21de4f6194dec9e3c401934db92c25e7 +1;
assign wire_qout_00003_00016      = sum0_00003 +  ~I57d0920119f8901bd4dea2d5f8fb5d90 +1;
assign wire_qout_00003_00017      = sum0_00003 +  ~I89537301987d6da0dbe6cff3caab3ff4 +1;
assign wire_qout_00003_00018      = sum0_00003 +  ~Iaf0bbbe791bb71d0f557dc71caa5fb87 +1;
assign wire_qout_00003_00019      = sum0_00003 +  ~Ic7ff9cde71054c1ee9eef81eabdd7061 +1;
assign wire_qout_00003_00020      = sum0_00003 +  ~I88c10c47ae424fbdcb852fbf1e94127c +1;
assign wire_qout_00003_00021      = sum0_00003 +  ~Icd2e75e47cab1d539ba9ff1b6e1d7155 +1;
assign wire_qout_00004_00000      = sum0_00004 +  ~I37e6bc7aff363ed0ed1f84b23c5f3e34 +1;
assign wire_qout_00004_00001      = sum0_00004 +  ~I733605337bf6972630c089d32fd7f98f +1;
assign wire_qout_00004_00002      = sum0_00004 +  ~Idcb1d8bbdeaed6768c2a418c3048e6ee +1;
assign wire_qout_00004_00003      = sum0_00004 +  ~Ia89da2f1890524ad3519ab403dd0686c +1;
assign wire_qout_00004_00004      = sum0_00004 +  ~Ie33a780b0221084898c9fc5b237b244a +1;
assign wire_qout_00004_00005      = sum0_00004 +  ~Iabbd1668e0014df518ede5216232834c +1;
assign wire_qout_00004_00006      = sum0_00004 +  ~Ibd89458312687610aa166a9538968851 +1;
assign wire_qout_00004_00007      = sum0_00004 +  ~Icbaf92a8e9875bcb19a1d074779a9ea5 +1;
assign wire_qout_00004_00008      = sum0_00004 +  ~I80f3c8559da8e97bc5397bb8b621a0bd +1;
assign wire_qout_00004_00009      = sum0_00004 +  ~I7a0eada108891aba06cecab5071232c9 +1;
assign wire_qout_00004_00010      = sum0_00004 +  ~Ie21a2c9b22e7bf8425fb5c0f33e5f4f7 +1;
assign wire_qout_00004_00011      = sum0_00004 +  ~Iaa5b2807e5cc2403c5787eeb3d10ca6b +1;
assign wire_qout_00004_00012      = sum0_00004 +  ~I6da2b3a481ee71b85f3087b36b399288 +1;
assign wire_qout_00004_00013      = sum0_00004 +  ~I11094e852295755925c3c61f1df81643 +1;
assign wire_qout_00004_00014      = sum0_00004 +  ~I9c633aa620cca127b0ff8cf882178e76 +1;
assign wire_qout_00004_00015      = sum0_00004 +  ~I694d471fd353eb54aae08a2afa7b645a +1;
assign wire_qout_00004_00016      = sum0_00004 +  ~I816704585ad393f685731104ad3ec64f +1;
assign wire_qout_00004_00017      = sum0_00004 +  ~I85d95015a9ce27a18ccbf73bbbcdbd70 +1;
assign wire_qout_00004_00018      = sum0_00004 +  ~I992e7c551b4aa818606c3465d33eb798 +1;
assign wire_qout_00004_00019      = sum0_00004 +  ~I2ead0e9941e2280309ab53535b1e1ac1 +1;
assign wire_qout_00004_00020      = sum0_00004 +  ~I56873feb8418005b5661c7382f2dbeec +1;
assign wire_qout_00004_00021      = sum0_00004 +  ~Ib6ea4a822da2ea32e0abf6cf8a33d295 +1;
assign wire_qout_00004_00022      = sum0_00004 +  ~Id1659ccdeaea3e59eb2d3f65a65ebd05 +1;
assign wire_qout_00005_00000      = sum0_00005 +  ~Ic2171967791a0329f3e39fc19d0a6bc8 +1;
assign wire_qout_00005_00001      = sum0_00005 +  ~I7d5041a6796c00188f74936d283defe6 +1;
assign wire_qout_00005_00002      = sum0_00005 +  ~Iba7608ee0a01af103e022bcaf564bf6b +1;
assign wire_qout_00005_00003      = sum0_00005 +  ~Iedbe9d0e48bd36064f59faea51afddb9 +1;
assign wire_qout_00005_00004      = sum0_00005 +  ~Ic3871325d57b310c95ca02fcaca529eb +1;
assign wire_qout_00005_00005      = sum0_00005 +  ~I42f9b1f8ef24ad56c10086852678b456 +1;
assign wire_qout_00005_00006      = sum0_00005 +  ~I3ed5d0fca86f35b3d4b4a89c6147d0cd +1;
assign wire_qout_00005_00007      = sum0_00005 +  ~Ib0126fb335e32793c400a97c5a4a337c +1;
assign wire_qout_00005_00008      = sum0_00005 +  ~I20590d8fb97ec0b2164ffe17826136a7 +1;
assign wire_qout_00005_00009      = sum0_00005 +  ~I3c128efc9f80c9b8334bf7b61de71b43 +1;
assign wire_qout_00005_00010      = sum0_00005 +  ~Ic7147944f8835e26b9838fdbdc18ca41 +1;
assign wire_qout_00005_00011      = sum0_00005 +  ~I698b1dbc9d8664d1c86c7a763d97b3b7 +1;
assign wire_qout_00005_00012      = sum0_00005 +  ~I508bbade361787127e1a2e8687ec884c +1;
assign wire_qout_00005_00013      = sum0_00005 +  ~I2afeb2a7b199c0c6738938f156ae4274 +1;
assign wire_qout_00005_00014      = sum0_00005 +  ~I86255756ddd1f88b74e070b19f8c3bfa +1;
assign wire_qout_00005_00015      = sum0_00005 +  ~I7d4924388dc5373ad7936dca76797473 +1;
assign wire_qout_00005_00016      = sum0_00005 +  ~Ie317e5ea2ca4ba2060d0f491290af96f +1;
assign wire_qout_00005_00017      = sum0_00005 +  ~I56ea52c50a188ec47e48740839a031c9 +1;
assign wire_qout_00005_00018      = sum0_00005 +  ~Id9b9a8fe43992ec0793845715dd2226c +1;
assign wire_qout_00005_00019      = sum0_00005 +  ~I93b69bfb228db4b569a6772179d603be +1;
assign wire_qout_00005_00020      = sum0_00005 +  ~I71afab29cdb962e1f1ca21b61dfb50c6 +1;
assign wire_qout_00005_00021      = sum0_00005 +  ~I9905e2686b350e8a6e7f790563a91294 +1;
assign wire_qout_00005_00022      = sum0_00005 +  ~I524e78ae6a4204e17ba4532dba047d4b +1;
assign wire_qout_00006_00000      = sum0_00006 +  ~I71228fe4188ab1d9796081184a422094 +1;
assign wire_qout_00006_00001      = sum0_00006 +  ~Ie19b39200436b0bfca13502ad36c21b9 +1;
assign wire_qout_00006_00002      = sum0_00006 +  ~If6657f90c84ca5e2ba08ec705f34be03 +1;
assign wire_qout_00006_00003      = sum0_00006 +  ~I60ec7459bbe99fce295406bee1f2af46 +1;
assign wire_qout_00006_00004      = sum0_00006 +  ~I29ab844f80c105d247c5c15faa35863c +1;
assign wire_qout_00006_00005      = sum0_00006 +  ~I856fa68463aa5ef1ae53442699d38b33 +1;
assign wire_qout_00006_00006      = sum0_00006 +  ~Ic3d00a27f15f8983a120395082854d6b +1;
assign wire_qout_00006_00007      = sum0_00006 +  ~I6b1d01c3cb8fb51e43cdb788b89816be +1;
assign wire_qout_00006_00008      = sum0_00006 +  ~Ib74a56900c1f8b159ad381f61acee801 +1;
assign wire_qout_00006_00009      = sum0_00006 +  ~Ia5eba52d169755c507b9e0094e467fab +1;
assign wire_qout_00006_00010      = sum0_00006 +  ~I0899e8fec1a7209cd94757c0b2f87c9a +1;
assign wire_qout_00006_00011      = sum0_00006 +  ~I08ece7cd684e593e02321612b7a88cee +1;
assign wire_qout_00006_00012      = sum0_00006 +  ~I691c84d81c60a462e28e2b2bae3ea845 +1;
assign wire_qout_00006_00013      = sum0_00006 +  ~I58dc9cce6384160c0a85c6efb3319cdb +1;
assign wire_qout_00006_00014      = sum0_00006 +  ~I56bf74b5890ec67090f499afdc0a9c88 +1;
assign wire_qout_00006_00015      = sum0_00006 +  ~Ibaf2f1f8bda2f6b932dc30f8369c0e1f +1;
assign wire_qout_00006_00016      = sum0_00006 +  ~Id9364a29fd79b52d0442e18dc0227854 +1;
assign wire_qout_00006_00017      = sum0_00006 +  ~Ica3a41ace27f7d94377981079952f4f7 +1;
assign wire_qout_00006_00018      = sum0_00006 +  ~Ib57795a63d642a73456324bab41384b6 +1;
assign wire_qout_00006_00019      = sum0_00006 +  ~Iabf572c97b48c6a7dcc19e56676e3a82 +1;
assign wire_qout_00006_00020      = sum0_00006 +  ~Iefd370d0df1a93639af482f78a1e8706 +1;
assign wire_qout_00006_00021      = sum0_00006 +  ~I995d2809ffaf0ecda6a004d01cb9c8c4 +1;
assign wire_qout_00006_00022      = sum0_00006 +  ~I4e8ebc46bc068c3f9889d970db131112 +1;
assign wire_qout_00007_00000      = sum0_00007 +  ~I7b561638da1b4a45ff59be81243e4471 +1;
assign wire_qout_00007_00001      = sum0_00007 +  ~If0a3b88a66a816b25f17ced5d0e8f775 +1;
assign wire_qout_00007_00002      = sum0_00007 +  ~I0374ada4fe50717f2158468b7ad205d4 +1;
assign wire_qout_00007_00003      = sum0_00007 +  ~I357137b41bb91e0659b1ac6ead9b5c12 +1;
assign wire_qout_00007_00004      = sum0_00007 +  ~I5d70bc64cf7b3d3ef4180e082e533237 +1;
assign wire_qout_00007_00005      = sum0_00007 +  ~I7d9ad929660cd212387d893266b681da +1;
assign wire_qout_00007_00006      = sum0_00007 +  ~I34be4b353cf75603301372840c2f91c2 +1;
assign wire_qout_00007_00007      = sum0_00007 +  ~I14834fc8e6489775359bcecf5a37ff4d +1;
assign wire_qout_00007_00008      = sum0_00007 +  ~I633a74e4dfa841c9fd13dbb6564c8493 +1;
assign wire_qout_00007_00009      = sum0_00007 +  ~I157bd468200e63385583b9045758d81e +1;
assign wire_qout_00007_00010      = sum0_00007 +  ~I918c46173eebc5b2a95e041cfd91d958 +1;
assign wire_qout_00007_00011      = sum0_00007 +  ~I4f8792c18bd07b23e82bbc44b4ca947f +1;
assign wire_qout_00007_00012      = sum0_00007 +  ~I8d0a1ae4c47edf1f2b99d1175aaa7197 +1;
assign wire_qout_00007_00013      = sum0_00007 +  ~I734e601f5f9d568a44a48834559e04db +1;
assign wire_qout_00007_00014      = sum0_00007 +  ~Ie421da1dc5aaea57c50d0c7d9c5a2717 +1;
assign wire_qout_00007_00015      = sum0_00007 +  ~Ief5cbddfbfb98fce4812a676849b9a98 +1;
assign wire_qout_00007_00016      = sum0_00007 +  ~Id113cab2dd1949d32e3c1c15273185c8 +1;
assign wire_qout_00007_00017      = sum0_00007 +  ~Icfe1a689e33b2b9aa9dba692d6d610b9 +1;
assign wire_qout_00007_00018      = sum0_00007 +  ~Ia4b671f3360f3ce55db0dc0e4d78ddbe +1;
assign wire_qout_00007_00019      = sum0_00007 +  ~I60cbd4369e7ba9b6532f279e5c59084c +1;
assign wire_qout_00007_00020      = sum0_00007 +  ~Ifb6c65a00d9a2c31d8b1119b949828d8 +1;
assign wire_qout_00007_00021      = sum0_00007 +  ~I4a777f0dd62b19dd340ad31517c4e789 +1;
assign wire_qout_00007_00022      = sum0_00007 +  ~Ib75747cb32130d44b338ed8c8af8ca11 +1;
assign wire_qout_00008_00000      = sum0_00008 +  ~Ic7e35cf8d5cd230b94c40714f16e2418 +1;
assign wire_qout_00008_00001      = sum0_00008 +  ~Ic51bb9184dfd103703cd0c6ad6edff4b +1;
assign wire_qout_00008_00002      = sum0_00008 +  ~I103f1449c78c47396d6a54dc1c810934 +1;
assign wire_qout_00008_00003      = sum0_00008 +  ~I56b3a97dc3037f0bb2eed93a9482c813 +1;
assign wire_qout_00008_00004      = sum0_00008 +  ~I51e98035b35a35fdc52f5bab8f19c152 +1;
assign wire_qout_00008_00005      = sum0_00008 +  ~Ia6a7f9beaceb08d81012f0e72171252f +1;
assign wire_qout_00008_00006      = sum0_00008 +  ~I21b062856ced09cb9131c01b5e166f32 +1;
assign wire_qout_00008_00007      = sum0_00008 +  ~I4f1221ce7880729fe584b42ef3afe6b2 +1;
assign wire_qout_00008_00008      = sum0_00008 +  ~Ie7f3f1d6cee7f02ae1b17740ed54c049 +1;
assign wire_qout_00008_00009      = sum0_00008 +  ~Ib196f5bcf9152703dc32c5101076600a +1;
assign wire_qout_00009_00000      = sum0_00009 +  ~Ide9ef5a16d8fe32353c2c2a30e8ee3b0 +1;
assign wire_qout_00009_00001      = sum0_00009 +  ~Iee6f2484a381bd42e441ff072ec582e4 +1;
assign wire_qout_00009_00002      = sum0_00009 +  ~I53121a39de0bcba91a4d0438be2ae958 +1;
assign wire_qout_00009_00003      = sum0_00009 +  ~Iff7950f24f0a6b0073942c37fff49d37 +1;
assign wire_qout_00009_00004      = sum0_00009 +  ~Ide86f019e9573706c25bd8b4552396a8 +1;
assign wire_qout_00009_00005      = sum0_00009 +  ~I2370042234b0e93bb66e44b97fca3e43 +1;
assign wire_qout_00009_00006      = sum0_00009 +  ~If9efe7a1c359ec03014a52870ac13aec +1;
assign wire_qout_00009_00007      = sum0_00009 +  ~I6a6eb62960b616043415406ebfc21346 +1;
assign wire_qout_00009_00008      = sum0_00009 +  ~I06c7728ef64be8311f48d10d766d0c44 +1;
assign wire_qout_00009_00009      = sum0_00009 +  ~I9fe11f6c8147391aa4a5afd1a4e4f731 +1;
assign wire_qout_00010_00000      = sum0_00010 +  ~Id50edc56fce48130247fdbc42eeff9ea +1;
assign wire_qout_00010_00001      = sum0_00010 +  ~If3e5161254eb9056914c46263b865c10 +1;
assign wire_qout_00010_00002      = sum0_00010 +  ~I58703e8b6d04f8c69ac38f5fcfdc4efc +1;
assign wire_qout_00010_00003      = sum0_00010 +  ~Ie1f41720e296ced1b74cb325b666d88f +1;
assign wire_qout_00010_00004      = sum0_00010 +  ~I5d5701435c96f1078e741921b56e3c65 +1;
assign wire_qout_00010_00005      = sum0_00010 +  ~Id96e744d9b10dcddd1ae0115ea57a76a +1;
assign wire_qout_00010_00006      = sum0_00010 +  ~I0c0060fe260afa3cdc72f35ffb6938ff +1;
assign wire_qout_00010_00007      = sum0_00010 +  ~Iaec1f186cb4a65da21d41e637fc628f7 +1;
assign wire_qout_00010_00008      = sum0_00010 +  ~I9c15a6a5c0db11ede80ff6d04c9a56d8 +1;
assign wire_qout_00010_00009      = sum0_00010 +  ~I8922487573e02d684a3d71448c3828f5 +1;
assign wire_qout_00011_00000      = sum0_00011 +  ~I47f17afcd5871fc3ac378316fd3d7ae9 +1;
assign wire_qout_00011_00001      = sum0_00011 +  ~Ia9642d79bb50567348083b4435c7d66d +1;
assign wire_qout_00011_00002      = sum0_00011 +  ~I2b2bd845428c49346ef8e94e95b618f8 +1;
assign wire_qout_00011_00003      = sum0_00011 +  ~Ib730fdb59198f23d1e590f6d6039e96a +1;
assign wire_qout_00011_00004      = sum0_00011 +  ~I644e83f0a7d432fba38ffb2d99088eca +1;
assign wire_qout_00011_00005      = sum0_00011 +  ~I97f2b15ce0a74e68d5a4438111adcb0a +1;
assign wire_qout_00011_00006      = sum0_00011 +  ~I84c88b631bed5311cb6e99e58941149e +1;
assign wire_qout_00011_00007      = sum0_00011 +  ~I45c5e6710240685bf54b73b0d7a64271 +1;
assign wire_qout_00011_00008      = sum0_00011 +  ~I5827bc87b5db1801b7db16e1e61515db +1;
assign wire_qout_00011_00009      = sum0_00011 +  ~I1c85c8f73ef80a6808c6aec0c8eca8ab +1;
assign wire_qout_00012_00000      = sum0_00012 +  ~Id13c99b7f7500c8195b54627efbc4232 +1;
assign wire_qout_00012_00001      = sum0_00012 +  ~I4636821315d702a677dc93113872e647 +1;
assign wire_qout_00012_00002      = sum0_00012 +  ~I9c981b0614a29386ca5e8ebc06a17f15 +1;
assign wire_qout_00012_00003      = sum0_00012 +  ~I4df3d4dac24877b14e6d361bafc1a800 +1;
assign wire_qout_00012_00004      = sum0_00012 +  ~I913d818403024510c55b65b56a38dd89 +1;
assign wire_qout_00013_00000      = sum0_00013 +  ~I57015930f5b09a6c6b030ed01dad2177 +1;
assign wire_qout_00013_00001      = sum0_00013 +  ~Ib54d55a70605119e37e9898b940ff636 +1;
assign wire_qout_00013_00002      = sum0_00013 +  ~If7e146da4f3bd255b8457fd6902005f6 +1;
assign wire_qout_00013_00003      = sum0_00013 +  ~Ied00d87af99ae55144fdde41ebfc1357 +1;
assign wire_qout_00013_00004      = sum0_00013 +  ~I7774313f1ae5a2de98855aad572b3676 +1;
assign wire_qout_00014_00000      = sum0_00014 +  ~I679baea452c3c6d04c53baa88edd8eb3 +1;
assign wire_qout_00014_00001      = sum0_00014 +  ~If4132b39ddb92aa02d8d0346fb0e6691 +1;
assign wire_qout_00014_00002      = sum0_00014 +  ~Iba70e737d52e6812a67c159520e5192f +1;
assign wire_qout_00014_00003      = sum0_00014 +  ~Ib9ceb8315f0cd848f861bab677c2c694 +1;
assign wire_qout_00014_00004      = sum0_00014 +  ~I7846bc2cc11e08d05f7c853c4920d555 +1;
assign wire_qout_00015_00000      = sum0_00015 +  ~I0865623d3350645e63fa6e6c9b78ac57 +1;
assign wire_qout_00015_00001      = sum0_00015 +  ~I0262b30a4efa9f1cfb11d1c3940de9e7 +1;
assign wire_qout_00015_00002      = sum0_00015 +  ~I7a2e79d42779ad235bca6ce3757cf588 +1;
assign wire_qout_00015_00003      = sum0_00015 +  ~I09e9a3cd4c12d204f760758e873a177b +1;
assign wire_qout_00015_00004      = sum0_00015 +  ~I30b0b1d54912c1a41a02a25ab238bb54 +1;
assign wire_qout_00016_00000      = sum0_00016 +  ~I49fb0909ddf66fc0073e6400f1a07844 +1;
assign wire_qout_00016_00001      = sum0_00016 +  ~I9938397dc94002481984f5b560fadc58 +1;
assign wire_qout_00016_00002      = sum0_00016 +  ~I4378d139db4b710e3587aa72df22b70d +1;
assign wire_qout_00016_00003      = sum0_00016 +  ~Ifa43d74fa91b7b9884969f575ef9ca8e +1;
assign wire_qout_00016_00004      = sum0_00016 +  ~I7c19a79f441ecbb73685db5a505e7479 +1;
assign wire_qout_00017_00000      = sum0_00017 +  ~If2af8106efc1f7dd02c074af68278b3d +1;
assign wire_qout_00017_00001      = sum0_00017 +  ~I89a3f8d5f760d1a650f85814cbfdc017 +1;
assign wire_qout_00017_00002      = sum0_00017 +  ~Ifae345c79662c3df3dff0fe68ad68746 +1;
assign wire_qout_00017_00003      = sum0_00017 +  ~I88a61cf72347d695489909d0819332ab +1;
assign wire_qout_00017_00004      = sum0_00017 +  ~I9aaa036a6158d11c235bdc8406d79f4c +1;
assign wire_qout_00018_00000      = sum0_00018 +  ~Ie8df350430970b5f1229cda772440f85 +1;
assign wire_qout_00018_00001      = sum0_00018 +  ~I7d77ac9b64b2e8cae21c6e36947e3ca2 +1;
assign wire_qout_00018_00002      = sum0_00018 +  ~Ic1faed76fca5a9ceb7db26c2f43623d9 +1;
assign wire_qout_00018_00003      = sum0_00018 +  ~I3ca2b9b77ed8d78a10aff42a07a53b07 +1;
assign wire_qout_00018_00004      = sum0_00018 +  ~I1f00849ea055a7893df386aed162a7b6 +1;
assign wire_qout_00019_00000      = sum0_00019 +  ~Iaf8a19fde3de660c3fa925593bebbe0c +1;
assign wire_qout_00019_00001      = sum0_00019 +  ~Icd1da43a4d95230e79dbd35a7ae41066 +1;
assign wire_qout_00019_00002      = sum0_00019 +  ~Ice9079fb6e08d629f8c0c9ce332c8f11 +1;
assign wire_qout_00019_00003      = sum0_00019 +  ~I15fafe2baba4d2f28037023a81ce0a81 +1;
assign wire_qout_00019_00004      = sum0_00019 +  ~If4d5b48882e9e628cf51ad2ac2f38c22 +1;
assign wire_qout_00020_00000      = sum0_00020 +  ~Id0eef1adba01447c14a6f005782dd9a2 +1;
assign wire_qout_00020_00001      = sum0_00020 +  ~I1d1a7c5928982c278d068ebd262254da +1;
assign wire_qout_00020_00002      = sum0_00020 +  ~I6354a0e638340378124e4df7f3d145b8 +1;
assign wire_qout_00020_00003      = sum0_00020 +  ~I0236c912c6d684bf4862b725be9d5951 +1;
assign wire_qout_00020_00004      = sum0_00020 +  ~I6f3be51d69b2b64a04e55b8946d5dd56 +1;
assign wire_qout_00020_00005      = sum0_00020 +  ~Icde3e6dbcf985682041f30903ad95572 +1;
assign wire_qout_00020_00006      = sum0_00020 +  ~I46ee30b46020d91707689f3468f00e26 +1;
assign wire_qout_00020_00007      = sum0_00020 +  ~I2605f078c1a9006c93855a9a2b0cf6b9 +1;
assign wire_qout_00020_00008      = sum0_00020 +  ~I4d226dd2f0bfcdbea6a2e6a6613c1b64 +1;
assign wire_qout_00020_00009      = sum0_00020 +  ~I5c942076b173cf527e1be2ddb8560e84 +1;
assign wire_qout_00020_00010      = sum0_00020 +  ~Ic95191bccb18e26c10e56be395ca6b1a +1;
assign wire_qout_00020_00011      = sum0_00020 +  ~Ia284f974dd8a526f31eb81ed71a06e94 +1;
assign wire_qout_00020_00012      = sum0_00020 +  ~Icc93450a007cee4c0a42717ed7600528 +1;
assign wire_qout_00020_00013      = sum0_00020 +  ~I9ec9f389d0489908d497487e44c6edcd +1;
assign wire_qout_00021_00000      = sum0_00021 +  ~If8a527cc7f06a9963a80a880d225d34c +1;
assign wire_qout_00021_00001      = sum0_00021 +  ~I39ff4663007dbc89b403f3b08a69bb6c +1;
assign wire_qout_00021_00002      = sum0_00021 +  ~I9590eb28a81c730b83b92ef7653e71a1 +1;
assign wire_qout_00021_00003      = sum0_00021 +  ~I2ba1acca919bddcc22a41a28d43a4e3e +1;
assign wire_qout_00021_00004      = sum0_00021 +  ~I62d8efd4227cb3dc88aa08b6585fafc8 +1;
assign wire_qout_00021_00005      = sum0_00021 +  ~I749e987266a20840bb8a4b1a2a2fc5b0 +1;
assign wire_qout_00021_00006      = sum0_00021 +  ~I7607af5d98e8070e3d15cee23cdf877e +1;
assign wire_qout_00021_00007      = sum0_00021 +  ~I2e11a697d7f17ac30302eadb500de72d +1;
assign wire_qout_00021_00008      = sum0_00021 +  ~Ia0886ce792e062e22d0c224158cdfb7d +1;
assign wire_qout_00021_00009      = sum0_00021 +  ~I6b3cd79aa87235ff174c0299b855dd3d +1;
assign wire_qout_00021_00010      = sum0_00021 +  ~Ie4ae993ddb776bdffec843db0def2f5c +1;
assign wire_qout_00021_00011      = sum0_00021 +  ~I3ed2da9b53daac0852a06ad1acfad21b +1;
assign wire_qout_00021_00012      = sum0_00021 +  ~Idefa29d4d4e2a6e9147f84893520096f +1;
assign wire_qout_00021_00013      = sum0_00021 +  ~Id1fbbe0594dae272856566522633bb3d +1;
assign wire_qout_00022_00000      = sum0_00022 +  ~I8070a3b7d8b1a7ae90c1a2d27aed09aa +1;
assign wire_qout_00022_00001      = sum0_00022 +  ~Ie88285ce2b9c71de02ebd62e8f44ca72 +1;
assign wire_qout_00022_00002      = sum0_00022 +  ~Ica1997c6c569c1d1f45224fbaa4e6b59 +1;
assign wire_qout_00022_00003      = sum0_00022 +  ~Iaf08bcaaeb15bb0c971432f7f8b16d0a +1;
assign wire_qout_00022_00004      = sum0_00022 +  ~Idcb37cfc357cc088c775409fb9225b51 +1;
assign wire_qout_00022_00005      = sum0_00022 +  ~Ic419255414995e7168afb97b051fa64f +1;
assign wire_qout_00022_00006      = sum0_00022 +  ~Iee6da3120d73373627b25ab7c0dedd28 +1;
assign wire_qout_00022_00007      = sum0_00022 +  ~I56fc99a22960232b305d6e683c66fcc7 +1;
assign wire_qout_00022_00008      = sum0_00022 +  ~I0a9a09b0ab43d2a0f1d1d01e13f0333c +1;
assign wire_qout_00022_00009      = sum0_00022 +  ~Ibc73d07e0c97a6fcae791e04106cb082 +1;
assign wire_qout_00022_00010      = sum0_00022 +  ~I224bbdf94ac86c5c376d1db4f4d4e060 +1;
assign wire_qout_00022_00011      = sum0_00022 +  ~I43f2b69c6b427de3095c44d4166b77cd +1;
assign wire_qout_00022_00012      = sum0_00022 +  ~I1e50c90010a3df1a8ce1cff811cc7a0c +1;
assign wire_qout_00022_00013      = sum0_00022 +  ~Ie1817cbf3a80dae435a5571dfbd2f5ad +1;
assign wire_qout_00023_00000      = sum0_00023 +  ~I0052d562fb3182890c8828e52d437b11 +1;
assign wire_qout_00023_00001      = sum0_00023 +  ~I1eedecb1d8ff505c75be7787199afada +1;
assign wire_qout_00023_00002      = sum0_00023 +  ~I7ef544597a185b1de63b4ffc4a1d44c2 +1;
assign wire_qout_00023_00003      = sum0_00023 +  ~Iadeedf3870f0b1eae98d0f7dbbeff04a +1;
assign wire_qout_00023_00004      = sum0_00023 +  ~I70ae07db9b44d530be220f06401d3d3d +1;
assign wire_qout_00023_00005      = sum0_00023 +  ~I7992ea31927b4f0e268462a3b0f18c5d +1;
assign wire_qout_00023_00006      = sum0_00023 +  ~Iadf927d18644a232ad1f1eba7db82934 +1;
assign wire_qout_00023_00007      = sum0_00023 +  ~I2a9c673cdd7ded79e09ada38c0f47e6f +1;
assign wire_qout_00023_00008      = sum0_00023 +  ~Ia86740e870d8063f0266b68ad6d7481d +1;
assign wire_qout_00023_00009      = sum0_00023 +  ~I6627bcdbaa8afb115123777abd45435b +1;
assign wire_qout_00023_00010      = sum0_00023 +  ~I96fe3eb633eff6958ac575b997460bb9 +1;
assign wire_qout_00023_00011      = sum0_00023 +  ~Iefdcb71f2903b11f5cb0b8857f7a1727 +1;
assign wire_qout_00023_00012      = sum0_00023 +  ~I2eb90278aaa54b9c8212b3b4af7c3617 +1;
assign wire_qout_00023_00013      = sum0_00023 +  ~I43493f70f0336453d77caf7f27503daa +1;
assign wire_qout_00024_00000      = sum0_00024 +  ~I26a7fe395eb583258c1ac58aaaa3234a +1;
assign wire_qout_00024_00001      = sum0_00024 +  ~I21668ff77cf75570cae97f575cbcf644 +1;
assign wire_qout_00024_00002      = sum0_00024 +  ~Ie48be9e6b6fd63baa104d0a6a4561a1a +1;
assign wire_qout_00024_00003      = sum0_00024 +  ~I05370777439b01811fe7f750d2f724f4 +1;
assign wire_qout_00024_00004      = sum0_00024 +  ~Icdcd83341f6b5c404f91ec7e97d0550c +1;
assign wire_qout_00024_00005      = sum0_00024 +  ~Ibba4e82d1510ddc16eb4ef64893cec02 +1;
assign wire_qout_00024_00006      = sum0_00024 +  ~Ifb00ae47340bc99669c71da34cccc59e +1;
assign wire_qout_00025_00000      = sum0_00025 +  ~I75a4cf2948bebc58e12bb039ed273ff2 +1;
assign wire_qout_00025_00001      = sum0_00025 +  ~I5a9fdec7d7ff99fe33ad6cd8afd9e059 +1;
assign wire_qout_00025_00002      = sum0_00025 +  ~I47b1695a74e4d27389b97543415dcc67 +1;
assign wire_qout_00025_00003      = sum0_00025 +  ~Ieb38fa62119a5a77c060d6634e051298 +1;
assign wire_qout_00025_00004      = sum0_00025 +  ~I3459d98131faef5a5040a03847890b55 +1;
assign wire_qout_00025_00005      = sum0_00025 +  ~Ie9b9221b2122087cd5f309570b6d31ca +1;
assign wire_qout_00025_00006      = sum0_00025 +  ~Id4451722e8e2393d627dcd0175dc9903 +1;
assign wire_qout_00026_00000      = sum0_00026 +  ~Ic10356f9069e3651b9c045c906e63512 +1;
assign wire_qout_00026_00001      = sum0_00026 +  ~Ic3a431f39c678b7175ed30fde1fa6424 +1;
assign wire_qout_00026_00002      = sum0_00026 +  ~Ib01cfd833a63500e03333f263805db3d +1;
assign wire_qout_00026_00003      = sum0_00026 +  ~I0b7b4c0a8503c751229edfe0237cc903 +1;
assign wire_qout_00026_00004      = sum0_00026 +  ~Iace01234164c8a9f7c98eeb83268745b +1;
assign wire_qout_00026_00005      = sum0_00026 +  ~Iace8b3b3a4c16763132b5aaa6b24212d +1;
assign wire_qout_00026_00006      = sum0_00026 +  ~I80a89644e278e96b1cd1c4b7f764dc34 +1;
assign wire_qout_00027_00000      = sum0_00027 +  ~Ia92d2276a8a23521ad1b88df7c27bc2e +1;
assign wire_qout_00027_00001      = sum0_00027 +  ~I39bbec42c442d1e8c818f46ad9c096a8 +1;
assign wire_qout_00027_00002      = sum0_00027 +  ~I88f1b5c12759a5efb2d2ded8483c9ed2 +1;
assign wire_qout_00027_00003      = sum0_00027 +  ~Iaf4ae293c576af16f5f43a8b86c1aa3d +1;
assign wire_qout_00027_00004      = sum0_00027 +  ~I68b575fcbc5321d4d26a22bcdbb506f6 +1;
assign wire_qout_00027_00005      = sum0_00027 +  ~Idf600b93ee1018ecf969ed7944b6bc7b +1;
assign wire_qout_00027_00006      = sum0_00027 +  ~I1cd93172cf5996bc870063aa642188a2 +1;
assign wire_qout_00028_00000      = sum0_00028 +  ~I4af080cb4e5cc525db95e5f401019e8c +1;
assign wire_qout_00028_00001      = sum0_00028 +  ~I6fc8044eb226a14ff1a786ddc96d2414 +1;
assign wire_qout_00028_00002      = sum0_00028 +  ~I27fd0073dbcdee599fbe85cf48806efc +1;
assign wire_qout_00028_00003      = sum0_00028 +  ~Iaee6d725a8b2653eeac6d5acb91f8f36 +1;
assign wire_qout_00028_00004      = sum0_00028 +  ~I4afdeba4fc2a12a6cbe3567a519367fc +1;
assign wire_qout_00028_00005      = sum0_00028 +  ~Ib42816335dd8475dcc78662c4c0786c1 +1;
assign wire_qout_00028_00006      = sum0_00028 +  ~I343c9efe71164c01e9c7d599e032864a +1;
assign wire_qout_00028_00007      = sum0_00028 +  ~I108c269ceec4adcff9afeda01101b838 +1;
assign wire_qout_00028_00008      = sum0_00028 +  ~I761983331fb6e3c6c437b3f1660f0b6b +1;
assign wire_qout_00028_00009      = sum0_00028 +  ~I70d32affde22f9dcb2d77430fca39069 +1;
assign wire_qout_00028_00010      = sum0_00028 +  ~Ic08e85346f61da036a15345a13ac12f0 +1;
assign wire_qout_00028_00011      = sum0_00028 +  ~If5dfdadb3868ed5a495007362f7db648 +1;
assign wire_qout_00028_00012      = sum0_00028 +  ~Ia1ee5579358b564de06c08ca418a9bf4 +1;
assign wire_qout_00029_00000      = sum0_00029 +  ~I9bb81dda8102b829441be46460eb8900 +1;
assign wire_qout_00029_00001      = sum0_00029 +  ~I8eef6ca0a61a21882ea28b3d63735228 +1;
assign wire_qout_00029_00002      = sum0_00029 +  ~I438522d92cce6f7010246424746ca255 +1;
assign wire_qout_00029_00003      = sum0_00029 +  ~I92496f68b44a94565af28a2c28d6fbae +1;
assign wire_qout_00029_00004      = sum0_00029 +  ~I66528f43f614f0edb715564eba3c77c1 +1;
assign wire_qout_00029_00005      = sum0_00029 +  ~I8cab9fba615b94fd4bb6934325be8ab8 +1;
assign wire_qout_00029_00006      = sum0_00029 +  ~I92d9fec22d36b1baac8bd78abfc1bbd5 +1;
assign wire_qout_00029_00007      = sum0_00029 +  ~I4eadce87f47df6d8f0e4acd057de5a09 +1;
assign wire_qout_00029_00008      = sum0_00029 +  ~I73203143fe37933c16fff873c1abf512 +1;
assign wire_qout_00029_00009      = sum0_00029 +  ~Ibed2a63af723a7abf96dacf1951e5266 +1;
assign wire_qout_00029_00010      = sum0_00029 +  ~Id667c80003b5541de9f84d3b8709c828 +1;
assign wire_qout_00029_00011      = sum0_00029 +  ~I02cbb4255db2b21ea32140f9e9ddb36b +1;
assign wire_qout_00029_00012      = sum0_00029 +  ~I65354f2069de0c25bbe7cd50fbe892aa +1;
assign wire_qout_00030_00000      = sum0_00030 +  ~Ic279867ebf3055980f3d813d5dc8dec6 +1;
assign wire_qout_00030_00001      = sum0_00030 +  ~I5c05da8a222ad5effb9815cbf3ec25f3 +1;
assign wire_qout_00030_00002      = sum0_00030 +  ~Ib8bf21f32c0e8b9cfa42a53807bfe3a3 +1;
assign wire_qout_00030_00003      = sum0_00030 +  ~I7208256bb198bfce1be71390b01bc028 +1;
assign wire_qout_00030_00004      = sum0_00030 +  ~I49f2a06ceb3a59773c65b19f54ff362b +1;
assign wire_qout_00030_00005      = sum0_00030 +  ~I86e495dc894d2aace15c1aff89798bf7 +1;
assign wire_qout_00030_00006      = sum0_00030 +  ~I0d53bb5344cabe5fa5ce3ecf7122a260 +1;
assign wire_qout_00030_00007      = sum0_00030 +  ~Ib2f5f5fc77ea8b529f2471c54388f2d1 +1;
assign wire_qout_00030_00008      = sum0_00030 +  ~Idcada1bfb3c0d1f2a09aab58a2071a57 +1;
assign wire_qout_00030_00009      = sum0_00030 +  ~I814b62120953991f9da055f118967e05 +1;
assign wire_qout_00030_00010      = sum0_00030 +  ~I123a212546a8ac394051425db4924812 +1;
assign wire_qout_00030_00011      = sum0_00030 +  ~Ie95f1a7e0effcec0aa423dc803056a13 +1;
assign wire_qout_00030_00012      = sum0_00030 +  ~I106deaff50b8480eac31ddbae2ec7c61 +1;
assign wire_qout_00031_00000      = sum0_00031 +  ~I68528be9951f5b8805411711cd11ea59 +1;
assign wire_qout_00031_00001      = sum0_00031 +  ~I0f034a8f077b0ab231727b6298e366d8 +1;
assign wire_qout_00031_00002      = sum0_00031 +  ~If9c12f8662333fb54a45cfa1bc5da487 +1;
assign wire_qout_00031_00003      = sum0_00031 +  ~Ie1681d905517daafcc7584725cd6014c +1;
assign wire_qout_00031_00004      = sum0_00031 +  ~I2ff3edcdb6158f1e3c9a555aeefc0850 +1;
assign wire_qout_00031_00005      = sum0_00031 +  ~I43b380be6df7df0d354223d0a0d6d6b6 +1;
assign wire_qout_00031_00006      = sum0_00031 +  ~I23eb1dc4d1c992f804dd04a2d823c778 +1;
assign wire_qout_00031_00007      = sum0_00031 +  ~I7f90f96c0260560ad5e6dc7448b2670a +1;
assign wire_qout_00031_00008      = sum0_00031 +  ~I07b417cdcc99eaea3413f563e26ddc73 +1;
assign wire_qout_00031_00009      = sum0_00031 +  ~I2f3ab9654e515a54e22e73d6c130ccc3 +1;
assign wire_qout_00031_00010      = sum0_00031 +  ~Iebdc41368d57498a04fa73e30b10a966 +1;
assign wire_qout_00031_00011      = sum0_00031 +  ~I5b4305bef5b4350c1d7ae143667afddd +1;
assign wire_qout_00031_00012      = sum0_00031 +  ~I2795d21d343b83a69146314a2407cfa2 +1;
assign wire_qout_00032_00000      = sum0_00032 +  ~Ic6386d7d8813731d612e24b715740275 +1;
assign wire_qout_00032_00001      = sum0_00032 +  ~I4c366a57920ff090a98a2cb8b9caa00b +1;
assign wire_qout_00032_00002      = sum0_00032 +  ~I14cf5d43fc9864820a8a25efcc5c6d86 +1;
assign wire_qout_00032_00003      = sum0_00032 +  ~I33b99994abbb5ecf8eed4de39033e4f8 +1;
assign wire_qout_00032_00004      = sum0_00032 +  ~I7c3291f0250d13ca94802b0b071a95c6 +1;
assign wire_qout_00032_00005      = sum0_00032 +  ~I2c926fd9d306e9ae13364e07c4b0395b +1;
assign wire_qout_00033_00000      = sum0_00033 +  ~Ib23edc35fa5bbfe0415fcf0861a22d9b +1;
assign wire_qout_00033_00001      = sum0_00033 +  ~I3e0e682047f7cc36142e668828cbff1e +1;
assign wire_qout_00033_00002      = sum0_00033 +  ~I99fb9030e8361e57818c07511479a9b8 +1;
assign wire_qout_00033_00003      = sum0_00033 +  ~Ic87c3d7762a18772972552162e1d1a8c +1;
assign wire_qout_00033_00004      = sum0_00033 +  ~I7e393e6c1d1bc44daaab120d55f5dd59 +1;
assign wire_qout_00033_00005      = sum0_00033 +  ~I448f126fd3932d5065abbe7bb2d92c56 +1;
assign wire_qout_00034_00000      = sum0_00034 +  ~Ifc8c6df8904b97674f2970ebc95b523c +1;
assign wire_qout_00034_00001      = sum0_00034 +  ~Icd0622a90782b9c451950e7ab0399567 +1;
assign wire_qout_00034_00002      = sum0_00034 +  ~I6493b3c087d4685a6b3f98c73dc2ff49 +1;
assign wire_qout_00034_00003      = sum0_00034 +  ~I20c2057240417146df144b518b43d052 +1;
assign wire_qout_00034_00004      = sum0_00034 +  ~Ied029d0bdea3bf134744c99426fa72dc +1;
assign wire_qout_00034_00005      = sum0_00034 +  ~Icb82c9ff4cb58159a1c3115c6fdd5f8c +1;
assign wire_qout_00035_00000      = sum0_00035 +  ~Ia3450e134e4086c35acbdee1e6042396 +1;
assign wire_qout_00035_00001      = sum0_00035 +  ~I5a0f27df5158309f32f0df31e8ae3ae3 +1;
assign wire_qout_00035_00002      = sum0_00035 +  ~I17d9e19854cef197fd3267618617efc3 +1;
assign wire_qout_00035_00003      = sum0_00035 +  ~I2993acb61f1abe529f8a60c94a438550 +1;
assign wire_qout_00035_00004      = sum0_00035 +  ~Ic8be2c94235fb40f78da33179ce4873a +1;
assign wire_qout_00035_00005      = sum0_00035 +  ~Ib3367565e4456da15e7c2315dccdb5e4 +1;
assign wire_qout_00036_00000      = sum0_00036 +  ~I15a1671def323cd294591564ae6ef8b1 +1;
assign wire_qout_00036_00001      = sum0_00036 +  ~Ic512effb493a06ece58a2af155135004 +1;
assign wire_qout_00036_00002      = sum0_00036 +  ~I2c72248cbe49ec0a0febac2437b8a6dc +1;
assign wire_qout_00036_00003      = sum0_00036 +  ~I964e17c41a134c080e9c43412a514f3f +1;
assign wire_qout_00036_00004      = sum0_00036 +  ~I94f1724740defe5bb7e40041d0e266a0 +1;
assign wire_qout_00036_00005      = sum0_00036 +  ~Ic19486b6ab0373b9c0ad8f7597782d8f +1;
assign wire_qout_00036_00006      = sum0_00036 +  ~I31243de90dc2a1656ca9d5e03bdd78da +1;
assign wire_qout_00036_00007      = sum0_00036 +  ~I242a30bdc8699d8ff550b25dd53d6c59 +1;
assign wire_qout_00037_00000      = sum0_00037 +  ~I9d15f76bb68b214057566cba4b511214 +1;
assign wire_qout_00037_00001      = sum0_00037 +  ~I9cc16a00912e7dfc05fb505a9db23cd8 +1;
assign wire_qout_00037_00002      = sum0_00037 +  ~Iacf9640cbf486411d6ceb8fe1a2fd5c9 +1;
assign wire_qout_00037_00003      = sum0_00037 +  ~I9015033ab0caf3fa41dae4de43f24a82 +1;
assign wire_qout_00037_00004      = sum0_00037 +  ~Ia630e59cbce82a570ae3890a6c0221e5 +1;
assign wire_qout_00037_00005      = sum0_00037 +  ~I4904ab14b19fa1b6befc218bc7be3842 +1;
assign wire_qout_00037_00006      = sum0_00037 +  ~I282d2eb4e74e034694e33273b9cb19d5 +1;
assign wire_qout_00037_00007      = sum0_00037 +  ~I3f33901c407a87e10d86c13c83dd52eb +1;
assign wire_qout_00038_00000      = sum0_00038 +  ~I43f41bf07836cee48069e9890c1de2a0 +1;
assign wire_qout_00038_00001      = sum0_00038 +  ~Id88480a0a350bb5fcf01ed5fff0bbd4c +1;
assign wire_qout_00038_00002      = sum0_00038 +  ~I1d9b9ff357667a362f0442f19986f451 +1;
assign wire_qout_00038_00003      = sum0_00038 +  ~Ice73589836da9028def6efb24a04dbbd +1;
assign wire_qout_00038_00004      = sum0_00038 +  ~Idb72c046c5996fbbd80b706666ffbd92 +1;
assign wire_qout_00038_00005      = sum0_00038 +  ~Ie5757e7b1647ab7d43cdbcf98cbb77fc +1;
assign wire_qout_00038_00006      = sum0_00038 +  ~I6072331f838d82329a07a4ffa340c7b6 +1;
assign wire_qout_00038_00007      = sum0_00038 +  ~Idf6875955525d80dc660ce956f4a84e7 +1;
assign wire_qout_00039_00000      = sum0_00039 +  ~Ia96955d9c0a8a587e0afab37c8415d8c +1;
assign wire_qout_00039_00001      = sum0_00039 +  ~Ifec374bce7f5507438f550df22d61a01 +1;
assign wire_qout_00039_00002      = sum0_00039 +  ~Ief67e897e57b96e2ec200e82bbc7caeb +1;
assign wire_qout_00039_00003      = sum0_00039 +  ~Ide604e9bbe35cb55892a4602e18b2527 +1;
assign wire_qout_00039_00004      = sum0_00039 +  ~I262f2390e77ec486ccd3a6ed05816e2d +1;
assign wire_qout_00039_00005      = sum0_00039 +  ~I280e20c20c0b4f26278b3de9b2ff84e4 +1;
assign wire_qout_00039_00006      = sum0_00039 +  ~Ib3a0307176d424a4733720416d71069d +1;
assign wire_qout_00039_00007      = sum0_00039 +  ~I76060709de3ea188748849f043c59ac0 +1;
assign wire_qout_00040_00000      = sum0_00040 +  ~I8be20605d26d218911e80a883a90d085 +1;
assign wire_qout_00040_00001      = sum0_00040 +  ~Ieafa9d74d4a61d28ac4a913db460bf33 +1;
assign wire_qout_00040_00002      = sum0_00040 +  ~I6fd1b4395af175eff85b3bfeef4c329b +1;
assign wire_qout_00040_00003      = sum0_00040 +  ~I39e6d3fb468aa40ea73535e81556ea65 +1;
assign wire_qout_00040_00004      = sum0_00040 +  ~Iae449b74e50e0907feae9e60f2329426 +1;
assign wire_qout_00040_00005      = sum0_00040 +  ~Iebf769a6bdaf214c1006c55c608d4eda +1;
assign wire_qout_00040_00006      = sum0_00040 +  ~Ia030c08757123aae947f86ab8bfb6d94 +1;
assign wire_qout_00040_00007      = sum0_00040 +  ~I8c35c5b343b552c22000e194c517ca12 +1;
assign wire_qout_00040_00008      = sum0_00040 +  ~Ibf80bb564263ea85bd886a8617f09bb2 +1;
assign wire_qout_00041_00000      = sum0_00041 +  ~Ib8dfd9b8badef282ca00a4f793c3c868 +1;
assign wire_qout_00041_00001      = sum0_00041 +  ~I596ad7e132f272cb196b74faa8c75aa4 +1;
assign wire_qout_00041_00002      = sum0_00041 +  ~Idc629414f6d0236ce0714cfaae23f065 +1;
assign wire_qout_00041_00003      = sum0_00041 +  ~I157fdf8775206858c08682db3039b084 +1;
assign wire_qout_00041_00004      = sum0_00041 +  ~Iacbb4daf5ce5c7eb1a2afe30d0cb5382 +1;
assign wire_qout_00041_00005      = sum0_00041 +  ~I4e08021c0235fafb60200aab97827a8f +1;
assign wire_qout_00041_00006      = sum0_00041 +  ~I730634ea15ac94d241f3ad2d6393a227 +1;
assign wire_qout_00041_00007      = sum0_00041 +  ~Iee367c535d9c39f872d2ec043e7e7b33 +1;
assign wire_qout_00041_00008      = sum0_00041 +  ~I68bb1f26f878862f288c1f57049cf58b +1;
assign wire_qout_00042_00000      = sum0_00042 +  ~Ia9b5d9ede006c56a6d83905529c77b7b +1;
assign wire_qout_00042_00001      = sum0_00042 +  ~I1487170cb1f3370ad45efc801cefc8ab +1;
assign wire_qout_00042_00002      = sum0_00042 +  ~Id88568dd34fbee42c9cb8cc15ac5c31d +1;
assign wire_qout_00042_00003      = sum0_00042 +  ~Ia30539545e66c4cfc16828140149180a +1;
assign wire_qout_00042_00004      = sum0_00042 +  ~Icbfbb37bad6344005dd233b3605a784f +1;
assign wire_qout_00042_00005      = sum0_00042 +  ~I91a6408a11fab36a8ba3dbd3f895a803 +1;
assign wire_qout_00042_00006      = sum0_00042 +  ~I47b878f27c30f79a37e97e022307e9e9 +1;
assign wire_qout_00042_00007      = sum0_00042 +  ~Ie76b0739aec66f8860870e66e87a6445 +1;
assign wire_qout_00042_00008      = sum0_00042 +  ~I50383e3d7c172eedfa00aa50a9faac4c +1;
assign wire_qout_00043_00000      = sum0_00043 +  ~Ifeaa99e03bda8ded058f98387de3d49d +1;
assign wire_qout_00043_00001      = sum0_00043 +  ~I4255ac1af4367c321567c4e46b06ab25 +1;
assign wire_qout_00043_00002      = sum0_00043 +  ~Ia445bdc7def7d8c1eec31ab892c25c41 +1;
assign wire_qout_00043_00003      = sum0_00043 +  ~Ic3b4752136ac08e343933ccc3a4ec47c +1;
assign wire_qout_00043_00004      = sum0_00043 +  ~Ica6707efd6d44ba6bbb87c0593a3d828 +1;
assign wire_qout_00043_00005      = sum0_00043 +  ~I739267bcc50c54b8a685cb3c6afc5cc1 +1;
assign wire_qout_00043_00006      = sum0_00043 +  ~I9160d11439c5140c0109b5190eb82e6b +1;
assign wire_qout_00043_00007      = sum0_00043 +  ~I6ff7b86cd7f63f9243646f1be10b2577 +1;
assign wire_qout_00043_00008      = sum0_00043 +  ~I165653ab165cfafe2b74cd441331f9e1 +1;
assign wire_qout_00044_00000      = sum0_00044 +  ~I08a8cd6965c23af6650568b654831b20 +1;
assign wire_qout_00044_00001      = sum0_00044 +  ~I9b6a674dbcbfcf65f1ae0deb8fc3566d +1;
assign wire_qout_00044_00002      = sum0_00044 +  ~Ie3a336de822ac7baf8486b1618ef1126 +1;
assign wire_qout_00044_00003      = sum0_00044 +  ~I5fc3c26d6c5aa893dfd5caa0f677233a +1;
assign wire_qout_00044_00004      = sum0_00044 +  ~Ie22b94121b58f17af14c75bfb27f96dd +1;
assign wire_qout_00044_00005      = sum0_00044 +  ~I0d9f8c99194d9d6e187b4ad02fcce8b4 +1;
assign wire_qout_00044_00006      = sum0_00044 +  ~I71e101962e766a4d1484b3235359a4b5 +1;
assign wire_qout_00044_00007      = sum0_00044 +  ~If2539da6722562bbf31786fd0036666a +1;
assign wire_qout_00044_00008      = sum0_00044 +  ~I22c8ccd4a9018ad1c129aa058bf579d8 +1;
assign wire_qout_00044_00009      = sum0_00044 +  ~I83330fef69470d2f5def8e6d7d9c50d2 +1;
assign wire_qout_00044_00010      = sum0_00044 +  ~I0539d598bbe3d50940329a282c801328 +1;
assign wire_qout_00044_00011      = sum0_00044 +  ~I202f88fdc946494d55fc8831c2e8a34c +1;
assign wire_qout_00044_00012      = sum0_00044 +  ~I3ee10f6a7785a236db317515fdd23a2d +1;
assign wire_qout_00044_00013      = sum0_00044 +  ~I453fdf4fbb5af5bd28a20d7643da9eb2 +1;
assign wire_qout_00044_00014      = sum0_00044 +  ~Ic4a6c02880a9aead7353332708e3f388 +1;
assign wire_qout_00044_00015      = sum0_00044 +  ~I7fb3b66cb48521f8715f66bf5642cdb2 +1;
assign wire_qout_00045_00000      = sum0_00045 +  ~I2fd872df07f50688486c0d602cfc5549 +1;
assign wire_qout_00045_00001      = sum0_00045 +  ~Iccefa45795486757515d95e5908b306a +1;
assign wire_qout_00045_00002      = sum0_00045 +  ~Ib1357cb20f471f1670ac2448f964f8eb +1;
assign wire_qout_00045_00003      = sum0_00045 +  ~Iab953a8974a1eb619dc0f074c003b5f9 +1;
assign wire_qout_00045_00004      = sum0_00045 +  ~I6e37582849c2c98fd15ad92d22c222da +1;
assign wire_qout_00045_00005      = sum0_00045 +  ~If004de0cac6e5f7701a1fce48c6936d5 +1;
assign wire_qout_00045_00006      = sum0_00045 +  ~Ic1efa395cc1fd2c5a1d1559fb169a5a0 +1;
assign wire_qout_00045_00007      = sum0_00045 +  ~I8e96c69e7d872be23229353808c34953 +1;
assign wire_qout_00045_00008      = sum0_00045 +  ~Ib6aded6c73a8cc3cb964b0ae895b859e +1;
assign wire_qout_00045_00009      = sum0_00045 +  ~I939368b76d98b43826c68c7f468a5632 +1;
assign wire_qout_00045_00010      = sum0_00045 +  ~I544f6263f16cd5e0b7cf28c511a8f6e3 +1;
assign wire_qout_00045_00011      = sum0_00045 +  ~I484545c4d2c869d79eb17f51e11070a3 +1;
assign wire_qout_00045_00012      = sum0_00045 +  ~I39289e6385a9bc378a9b8dd440249a7f +1;
assign wire_qout_00045_00013      = sum0_00045 +  ~Ie9cce5746a83479a567bbaeac6dbf497 +1;
assign wire_qout_00045_00014      = sum0_00045 +  ~Ic044d7419cc43736d278c2df33b4a3cc +1;
assign wire_qout_00045_00015      = sum0_00045 +  ~I6714551e8885ef5e4490673fe1b2dad1 +1;
assign wire_qout_00046_00000      = sum0_00046 +  ~Ie9ab3c88ac62369e3d92d110165a94a8 +1;
assign wire_qout_00046_00001      = sum0_00046 +  ~If38feb4f76f761dce6145731ad235d7f +1;
assign wire_qout_00046_00002      = sum0_00046 +  ~I6359856a1843d8c8b65dc478bccb3acd +1;
assign wire_qout_00046_00003      = sum0_00046 +  ~If6f3d91c3c7a43622b9a522492cd83d3 +1;
assign wire_qout_00046_00004      = sum0_00046 +  ~Id023a6298e65da1f4da3831f5136afc2 +1;
assign wire_qout_00046_00005      = sum0_00046 +  ~I6b24690f394792edb0d82b3b9e110851 +1;
assign wire_qout_00046_00006      = sum0_00046 +  ~I5b55c285f7e3e78447fee68532ab9f7f +1;
assign wire_qout_00046_00007      = sum0_00046 +  ~I32701d9e4b96853c53f0ab651a6a4ba2 +1;
assign wire_qout_00046_00008      = sum0_00046 +  ~I82f266e5792cdb6e7ebd264e246161f5 +1;
assign wire_qout_00046_00009      = sum0_00046 +  ~Ibfacfe5b83819afe7fbd4bffa2d6d4e2 +1;
assign wire_qout_00046_00010      = sum0_00046 +  ~Ib8e68a77ad8b9e7cf415bee17645c3f9 +1;
assign wire_qout_00046_00011      = sum0_00046 +  ~I644ee0055a55f54ab3544bb532e39c61 +1;
assign wire_qout_00046_00012      = sum0_00046 +  ~Ic5467e42aa377c6ffd8f70673808774f +1;
assign wire_qout_00046_00013      = sum0_00046 +  ~Ic57eb4a034247a4c952d8224ea9f2bac +1;
assign wire_qout_00046_00014      = sum0_00046 +  ~Ia642db613c0ec1ca4e69afde7a14a839 +1;
assign wire_qout_00046_00015      = sum0_00046 +  ~I432aa7cb844286c442356954f8814260 +1;
assign wire_qout_00047_00000      = sum0_00047 +  ~If520c1cd27f9d4bc52d0d029f693b660 +1;
assign wire_qout_00047_00001      = sum0_00047 +  ~Ie87075ac979410cc11099a356966b8a2 +1;
assign wire_qout_00047_00002      = sum0_00047 +  ~I6fab46b1766878b26b53f352fee98223 +1;
assign wire_qout_00047_00003      = sum0_00047 +  ~Ieaf14683f40374c4531326d228cb43c3 +1;
assign wire_qout_00047_00004      = sum0_00047 +  ~I5149125aaaad943d891df6a3c2be93a0 +1;
assign wire_qout_00047_00005      = sum0_00047 +  ~I770dff588ee1f52f58bea1921cb23383 +1;
assign wire_qout_00047_00006      = sum0_00047 +  ~I8f0a90e761111a613d2488285534a500 +1;
assign wire_qout_00047_00007      = sum0_00047 +  ~I765a8825e42180a6c63f7b33703bb483 +1;
assign wire_qout_00047_00008      = sum0_00047 +  ~I512cc8f6519aa08aee18225b56d47c9f +1;
assign wire_qout_00047_00009      = sum0_00047 +  ~If08370fd0e8af818c6db20f43e74034d +1;
assign wire_qout_00047_00010      = sum0_00047 +  ~I0ff382edfc8051459657ffa3899f5f73 +1;
assign wire_qout_00047_00011      = sum0_00047 +  ~I9d2864024148337277523ef7fa2e1600 +1;
assign wire_qout_00047_00012      = sum0_00047 +  ~I1c85a2d1df6749a194072eb731506bfe +1;
assign wire_qout_00047_00013      = sum0_00047 +  ~I3e3ce8b4ead150a6eae2e5c701c7b598 +1;
assign wire_qout_00047_00014      = sum0_00047 +  ~I45bc13ae0e0554a79c62cd9c6aa8f2a5 +1;
assign wire_qout_00047_00015      = sum0_00047 +  ~I92678f5b52c9c55556ff7f17f0f607b7 +1;
assign wire_qout_00048_00000      = sum0_00048 +  ~Ib4bdc9069d0c08655f5e87f705943eda +1;
assign wire_qout_00048_00001      = sum0_00048 +  ~Idbf9094c94c931f16fba468b9dd59a25 +1;
assign wire_qout_00048_00002      = sum0_00048 +  ~I1c3c4ce44610e04c5eef2fcbc2ea5114 +1;
assign wire_qout_00048_00003      = sum0_00048 +  ~Ie84be0ae8311d906eff08f7f5b214943 +1;
assign wire_qout_00048_00004      = sum0_00048 +  ~Ic90b98708faa8c8b75d4bd9a52c292f7 +1;
assign wire_qout_00048_00005      = sum0_00048 +  ~I8eba6f14f42701d22859fbea94bd1871 +1;
assign wire_qout_00048_00006      = sum0_00048 +  ~I6d83efa9f988328f487e9232bf2633a2 +1;
assign wire_qout_00048_00007      = sum0_00048 +  ~Ic23e01562c8a753fd70c343297be288a +1;
assign wire_qout_00048_00008      = sum0_00048 +  ~I5669856f88f5e2c98f64df696db76414 +1;
assign wire_qout_00049_00000      = sum0_00049 +  ~Ic3a608b850709286ea0ad2f67425d9ac +1;
assign wire_qout_00049_00001      = sum0_00049 +  ~I5267fa34449e6eebe891017fc32d0749 +1;
assign wire_qout_00049_00002      = sum0_00049 +  ~I599d01cfe6e54d8e45d64446c446818d +1;
assign wire_qout_00049_00003      = sum0_00049 +  ~I8f94dbafaac589ac9f14b56d4556ff96 +1;
assign wire_qout_00049_00004      = sum0_00049 +  ~I754563caea429d3d0e22df5d193b84eb +1;
assign wire_qout_00049_00005      = sum0_00049 +  ~If7f373506cac70f8ba1222db135c27e8 +1;
assign wire_qout_00049_00006      = sum0_00049 +  ~I69f563e7b7ad483893ac9c4684349769 +1;
assign wire_qout_00049_00007      = sum0_00049 +  ~Ia0a02781c674fe5d769206448d475245 +1;
assign wire_qout_00049_00008      = sum0_00049 +  ~I1b7a401bc11741e6f011fb9895b5c797 +1;
assign wire_qout_00050_00000      = sum0_00050 +  ~Ieb528d666fdb708279184bb59eac25d9 +1;
assign wire_qout_00050_00001      = sum0_00050 +  ~Ic3ff7ce12c836bf0693252b9a7a7cfe8 +1;
assign wire_qout_00050_00002      = sum0_00050 +  ~I19bba6a58ad3ef959b33701f82761984 +1;
assign wire_qout_00050_00003      = sum0_00050 +  ~I8acc93b34974c1e708b0e1591f7b2d3d +1;
assign wire_qout_00050_00004      = sum0_00050 +  ~Ib60d4ac0fcadcdfce5a14fb92f58423f +1;
assign wire_qout_00050_00005      = sum0_00050 +  ~I039f05d5be891a37e04556f1eae674d2 +1;
assign wire_qout_00050_00006      = sum0_00050 +  ~Id0f75e19b94541ed5c5c352d13390d2d +1;
assign wire_qout_00050_00007      = sum0_00050 +  ~Ife1190f76c2e251704c2960c23330a48 +1;
assign wire_qout_00050_00008      = sum0_00050 +  ~Id3e0c98bff2636e216b4d3a0ffd51054 +1;
assign wire_qout_00051_00000      = sum0_00051 +  ~If4d3b31b87c0f723241d35ce7e854eba +1;
assign wire_qout_00051_00001      = sum0_00051 +  ~I72369dedfe36cb22269033cc305b730c +1;
assign wire_qout_00051_00002      = sum0_00051 +  ~Iec71fe7fcebccf1ae0d10a5d187fcc44 +1;
assign wire_qout_00051_00003      = sum0_00051 +  ~Ie11da10808c4ca84f399535df6261307 +1;
assign wire_qout_00051_00004      = sum0_00051 +  ~I280fa9d114e227cd649bf0e55e845651 +1;
assign wire_qout_00051_00005      = sum0_00051 +  ~I94c4e11670b4233fa072517a8f19c901 +1;
assign wire_qout_00051_00006      = sum0_00051 +  ~I4dca2dd40a7127ce44f83b430a34c738 +1;
assign wire_qout_00051_00007      = sum0_00051 +  ~I1a24e98165afa62bd14986911a36fb6e +1;
assign wire_qout_00051_00008      = sum0_00051 +  ~Ife1164cad7cda4aa9a08d94dfe86add6 +1;
assign wire_qout_00052_00000      = sum0_00052 +  ~I8d8d95ff26f33f69a182b32ccde23905 +1;
assign wire_qout_00052_00001      = sum0_00052 +  ~I2508854bcbab37bd09c9465c377c06aa +1;
assign wire_qout_00052_00002      = sum0_00052 +  ~I140078292f7209eccacd53a8bab18016 +1;
assign wire_qout_00052_00003      = sum0_00052 +  ~I141fb1cbe09f9abe282cffd4de815d25 +1;
assign wire_qout_00052_00004      = sum0_00052 +  ~If79d1d378f7c6fd29fc3335ec5f5c51d +1;
assign wire_qout_00052_00005      = sum0_00052 +  ~I4a41999cea9357a85c73a0af509eeac9 +1;
assign wire_qout_00052_00006      = sum0_00052 +  ~I8e517c401d62dbb10dcc96ab536f6afb +1;
assign wire_qout_00052_00007      = sum0_00052 +  ~I8ad3627f171eadcc960a688ac0afcbc0 +1;
assign wire_qout_00052_00008      = sum0_00052 +  ~I85c4d3d6c8408c6f38741257ed177ca6 +1;
assign wire_qout_00052_00009      = sum0_00052 +  ~Id66c47fd69c175a4393e975a269cf053 +1;
assign wire_qout_00052_00010      = sum0_00052 +  ~I37dca40506d61bdeab1255ed4892ca20 +1;
assign wire_qout_00052_00011      = sum0_00052 +  ~I340c98b886123c541a1b8d9fc8a6d48c +1;
assign wire_qout_00053_00000      = sum0_00053 +  ~I2dc64c3b06588542b027f997437bee63 +1;
assign wire_qout_00053_00001      = sum0_00053 +  ~Id92a37c091100e9df08e24498ecb4022 +1;
assign wire_qout_00053_00002      = sum0_00053 +  ~I74a4b9365391fd20c34588002ad40547 +1;
assign wire_qout_00053_00003      = sum0_00053 +  ~I461195b7ae78743e09ee50486ad6ebe5 +1;
assign wire_qout_00053_00004      = sum0_00053 +  ~I356d747600182675699a2d2634d4c5ce +1;
assign wire_qout_00053_00005      = sum0_00053 +  ~I87d6a5d30c3e4202cf51f33c7a770c51 +1;
assign wire_qout_00053_00006      = sum0_00053 +  ~I960768a84aec9d5b8bc7c1c523024a25 +1;
assign wire_qout_00053_00007      = sum0_00053 +  ~I09b5273bb15d48a7fd78559930fa6d1c +1;
assign wire_qout_00053_00008      = sum0_00053 +  ~I5814a85c45fd0f7be21ed325235fe4b7 +1;
assign wire_qout_00053_00009      = sum0_00053 +  ~Ib06b60cf9933dd8952206c5f3ccced8e +1;
assign wire_qout_00053_00010      = sum0_00053 +  ~I67347c413b5efd8ff9e0d5bc7ab2a047 +1;
assign wire_qout_00053_00011      = sum0_00053 +  ~I72b1bb104bf2843f161448baf7aab44b +1;
assign wire_qout_00054_00000      = sum0_00054 +  ~Ib23d889edb5a6d9f27de977d3b1a2616 +1;
assign wire_qout_00054_00001      = sum0_00054 +  ~Ifaff9dd032cf96487be819c59b03000a +1;
assign wire_qout_00054_00002      = sum0_00054 +  ~I028ce03be0618b816e0ecdf43d4cd6e6 +1;
assign wire_qout_00054_00003      = sum0_00054 +  ~I6ae2523095237282533e0b5f1c26b488 +1;
assign wire_qout_00054_00004      = sum0_00054 +  ~I5aba6218461e8d571be03a3ef041ebaa +1;
assign wire_qout_00054_00005      = sum0_00054 +  ~I6ca8a1fa2c72b1c61d11dc7d1ba5f37b +1;
assign wire_qout_00054_00006      = sum0_00054 +  ~I3ec5819176ad4b0895a9118d90ab22b5 +1;
assign wire_qout_00054_00007      = sum0_00054 +  ~I49b64469d298012dbb131d879bff38d6 +1;
assign wire_qout_00054_00008      = sum0_00054 +  ~I95361d5f524ccb9feb42811af5c482e2 +1;
assign wire_qout_00054_00009      = sum0_00054 +  ~I9c4b34b5fb1d59c132bcaeb6258675df +1;
assign wire_qout_00054_00010      = sum0_00054 +  ~I613d4b1e3b9e812b785c9cf14fefdfe6 +1;
assign wire_qout_00054_00011      = sum0_00054 +  ~I848ed394bd4f0b199d11c0ff458394a7 +1;
assign wire_qout_00055_00000      = sum0_00055 +  ~Ie65a0634454381e24bb3223a333e3ad0 +1;
assign wire_qout_00055_00001      = sum0_00055 +  ~Iad166146f7df5e8068fc6efe4d3e4141 +1;
assign wire_qout_00055_00002      = sum0_00055 +  ~I63e45abd4d27219bddcef06108b72021 +1;
assign wire_qout_00055_00003      = sum0_00055 +  ~Id1bacd13718f7c29c26b63c239d04dd8 +1;
assign wire_qout_00055_00004      = sum0_00055 +  ~Ia3104c69fb4f7abfb5efa3874169a7ad +1;
assign wire_qout_00055_00005      = sum0_00055 +  ~Ie1b7257c99831ec5864f65958ecf14fb +1;
assign wire_qout_00055_00006      = sum0_00055 +  ~I4accbad1b451ed2b622e15ef9ae16d13 +1;
assign wire_qout_00055_00007      = sum0_00055 +  ~I5ce8b2f633011e89356243a1a71edeb6 +1;
assign wire_qout_00055_00008      = sum0_00055 +  ~I3e5139f24e3d082eb31b0e61ea9fa1aa +1;
assign wire_qout_00055_00009      = sum0_00055 +  ~I61cc8a0f49e393721a62a776e4793deb +1;
assign wire_qout_00055_00010      = sum0_00055 +  ~Ie631e40caade823a196370fc3358f042 +1;
assign wire_qout_00055_00011      = sum0_00055 +  ~I4c971e714427664c59c6371e14781bae +1;
assign wire_qout_00056_00000      = sum0_00056 +  ~I36ca732e811d67cd742d24fd4cae887b +1;
assign wire_qout_00057_00000      = sum0_00057 +  ~I354fdd241d5d07f0d8380fe8924e0a8c +1;
assign wire_qout_00058_00000      = sum0_00058 +  ~Id38b705f5d2863a020a475ffffc8afd6 +1;
assign wire_qout_00059_00000      = sum0_00059 +  ~Id6e5d67e7bb7c4b999459374ea80459a +1;
assign wire_qout_00060_00000      = sum0_00060 +  ~I05341013abd4206eb66fcddfd63bfe26 +1;
assign wire_qout_00061_00000      = sum0_00061 +  ~I15da71a21f5842cb65b543d9bc3e267b +1;
assign wire_qout_00062_00000      = sum0_00062 +  ~Iccf255fb3422c558465e45226068a16d +1;
assign wire_qout_00063_00000      = sum0_00063 +  ~I1c2674b2e6b269ed539827412c5199a5 +1;
assign wire_qout_00064_00000      = sum0_00064 +  ~I6a3f405bb4a0c4448d9b9d3dd95d036c +1;
assign wire_qout_00065_00000      = sum0_00065 +  ~Ib528bb7a64cce4f694081d151fa6fa86 +1;
assign wire_qout_00066_00000      = sum0_00066 +  ~Iaa40bd3abf668a21e0f87c7bda7b3f69 +1;
assign wire_qout_00067_00000      = sum0_00067 +  ~I919d36a7f6ad42c4bbc23222beb73106 +1;
assign wire_qout_00068_00000      = sum0_00068 +  ~I648d2a279dd1f587b1e45eeb35f2fa90 +1;
assign wire_qout_00069_00000      = sum0_00069 +  ~I194a64bef92ecf6714141eaa5d41c9d4 +1;
assign wire_qout_00070_00000      = sum0_00070 +  ~Id332e7f482524adeac7f7cdafcf5ca46 +1;
assign wire_qout_00071_00000      = sum0_00071 +  ~I226383d68f89db716cfd8d08b837865a +1;
assign wire_qout_00072_00000      = sum0_00072 +  ~I2bdf5d319ba9089a4da34b108f5c5ae5 +1;
assign wire_qout_00073_00000      = sum0_00073 +  ~Ia91800792941ec7cc60415c3f844e4ed +1;
assign wire_qout_00074_00000      = sum0_00074 +  ~Id7c507d96098ee7a955af8a48ee5d72a +1;
assign wire_qout_00075_00000      = sum0_00075 +  ~Ie15e4c1bcdb0e18085d4b320ac6a925c +1;
assign wire_qout_00076_00000      = sum0_00076 +  ~I5485d9edcafc6202f6e5f0969979802f +1;
assign wire_qout_00077_00000      = sum0_00077 +  ~I7fe364f9f537cbef782e7007848a1c10 +1;
assign wire_qout_00078_00000      = sum0_00078 +  ~I52dcf5bace9cadcf8a895aaa6a8c1da8 +1;
assign wire_qout_00079_00000      = sum0_00079 +  ~I13a9eec6175e695ab8bc4516cf57d6ec +1;
assign wire_qout_00080_00000      = sum0_00080 +  ~Iee73a7c685a4cee03f33d3ef379b1c8a +1;
assign wire_qout_00081_00000      = sum0_00081 +  ~I740dc91716e3906ad078e2c7cc3c925a +1;
assign wire_qout_00082_00000      = sum0_00082 +  ~I514d2dc697e9b39ba027c418a6df6cb9 +1;
assign wire_qout_00083_00000      = sum0_00083 +  ~I782726e317a2aada9e755bcbc4b0d3fa +1;
assign wire_qout_00084_00000      = sum0_00084 +  ~I11eb26cf0f0b3a334e8f7317bf8d9eb0 +1;
assign wire_qout_00085_00000      = sum0_00085 +  ~I26cb63ba20245b2c332b09e25c4409aa +1;
assign wire_qout_00086_00000      = sum0_00086 +  ~Idd7691d31f8d0c09ee988116d574ec59 +1;
assign wire_qout_00087_00000      = sum0_00087 +  ~Iecc02842a2d2b9b9e8187f2d39e62e05 +1;
assign wire_qout_00088_00000      = sum0_00088 +  ~I5551342f1751fc64f32744a46b9649be +1;
assign wire_qout_00089_00000      = sum0_00089 +  ~Iff7c29299f005c1cd5a16b64601e727e +1;
assign wire_qout_00090_00000      = sum0_00090 +  ~I17a5446e942bcc1dc2c96930e0a87a70 +1;
assign wire_qout_00091_00000      = sum0_00091 +  ~I719b67f84e07e90dfd29a8cd5d94cf39 +1;
assign wire_qout_00092_00000      = sum0_00092 +  ~I2c835dfb3596b8bf057a7cc21122c81f +1;
assign wire_qout_00093_00000      = sum0_00093 +  ~Ib71b3d357c98dcdfae5c777ca3082275 +1;
assign wire_qout_00094_00000      = sum0_00094 +  ~I086bf19f620c8a8f6888e775cb1ed7f4 +1;
assign wire_qout_00095_00000      = sum0_00095 +  ~I802c554d5b04af6b949677819a4966ed +1;
assign wire_qout_00096_00000      = sum0_00096 +  ~Iceefb06cb3715e1b41e6f7d89420e5ba +1;
assign wire_qout_00097_00000      = sum0_00097 +  ~I56948bc48c0220893d68004615a6ebaa +1;
assign wire_qout_00098_00000      = sum0_00098 +  ~Iec1368f034655d61354ab5b5e94d7d89 +1;
assign wire_qout_00099_00000      = sum0_00099 +  ~I1e43c0aeeb8a2461d208eba24967af30 +1;
assign wire_qout_00100_00000      = sum0_00100 +  ~Ia6eb85b127cf9c1a437611556296b967 +1;
assign wire_qout_00101_00000      = sum0_00101 +  ~Ieba89aa901e61218074af53a2484a74b +1;
assign wire_qout_00102_00000      = sum0_00102 +  ~I8b3b875c6c07bd97ba598a5139156fa4 +1;
assign wire_qout_00103_00000      = sum0_00103 +  ~I7b33ddad346077928620344542b9481e +1;
assign wire_qout_00104_00000      = sum0_00104 +  ~I11d967a5c5d14c88b5587d4cfed1d05f +1;
assign wire_qout_00105_00000      = sum0_00105 +  ~I27458d76b3ac6520fb379405c6b2956f +1;
assign wire_qout_00106_00000      = sum0_00106 +  ~I2525111a2fb5f10d64bbd16e148653b8 +1;
assign wire_qout_00107_00000      = sum0_00107 +  ~I7b7cbcd1c6d2a2eeaaff474536a69eed +1;
assign wire_qout_00108_00000      = sum0_00108 +  ~Id2a7f0781d18dccc7c4e0b383b7cddfa +1;
assign wire_qout_00109_00000      = sum0_00109 +  ~If8bc141d98ebe1be7fa81cde5c65868e +1;
assign wire_qout_00110_00000      = sum0_00110 +  ~I8645e1326c66f5efef4b9c923599d1a3 +1;
assign wire_qout_00111_00000      = sum0_00111 +  ~I0426ef66185128dd1ef4dbb68dcda585 +1;
assign wire_qout_00112_00000      = sum0_00112 +  ~Iddd954df5bae9b4240e0512f746669a9 +1;
assign wire_qout_00113_00000      = sum0_00113 +  ~I29e940970d87e8e09b26ab1b0b8f2286 +1;
assign wire_qout_00114_00000      = sum0_00114 +  ~I488f6d9676aa85a55d030bf12e8997a7 +1;
assign wire_qout_00115_00000      = sum0_00115 +  ~I99d761b75ade1fb2e8afbb1a77752609 +1;
assign wire_qout_00116_00000      = sum0_00116 +  ~Iac4e3d20178049f9c59abf374752dccc +1;
assign wire_qout_00117_00000      = sum0_00117 +  ~I618d33f26badabfa578908903a613bce +1;
assign wire_qout_00118_00000      = sum0_00118 +  ~I822d7973afe090b2764335f1b72dfd0e +1;
assign wire_qout_00119_00000      = sum0_00119 +  ~I12c1035353e553b3b6a13bb174ce6020 +1;
assign wire_qout_00120_00000      = sum0_00120 +  ~Ia6d61947d36fc128c689808c82db80f6 +1;
assign wire_qout_00121_00000      = sum0_00121 +  ~Ie9b042f686381739b9ff219041f1e0ce +1;
assign wire_qout_00122_00000      = sum0_00122 +  ~I0c4268c01aed70ce4fc71531bf4bb862 +1;
assign wire_qout_00123_00000      = sum0_00123 +  ~Ia34e42f8de91fa4861b0c6cac5dcfc29 +1;
assign wire_qout_00124_00000      = sum0_00124 +  ~Ib7c5850b4f7cc77be2048d114a2128d9 +1;
assign wire_qout_00125_00000      = sum0_00125 +  ~I32bb50faa2b246b2d3b462a79be597c5 +1;
assign wire_qout_00126_00000      = sum0_00126 +  ~Idc6d40a49f05c5422758cee50f787eb1 +1;
assign wire_qout_00127_00000      = sum0_00127 +  ~Ide1d7dc22a4b271ef764df14ac22366a +1;
assign wire_qout_00128_00000      = sum0_00128 +  ~I7ace6778ac86b3e05939a3fcc716136f +1;
assign wire_qout_00129_00000      = sum0_00129 +  ~I044e01e8d2df46e03f00a0af2beb0bf5 +1;
assign wire_qout_00130_00000      = sum0_00130 +  ~I45a7ddcda2662e36b7617dfe64514346 +1;
assign wire_qout_00131_00000      = sum0_00131 +  ~Idada779a1ac7b844867571d77054b657 +1;
assign wire_qout_00132_00000      = sum0_00132 +  ~Ieeba01b18a244ab8c0ac263c138fabcc +1;
assign wire_qout_00133_00000      = sum0_00133 +  ~Ie4c9797a955778694dd8615219cb51e7 +1;
assign wire_qout_00134_00000      = sum0_00134 +  ~I28a5ed4c239e64c76bb6e566b50cfd23 +1;
assign wire_qout_00135_00000      = sum0_00135 +  ~I79a705ee1e414fe4a5fb14e9b3ce9597 +1;
assign wire_qout_00136_00000      = sum0_00136 +  ~I04f90a907f10a7fa1ae3591b48094d5c +1;
assign wire_qout_00137_00000      = sum0_00137 +  ~I31d25b1b49e65216e90b39aa27acd6be +1;
assign wire_qout_00138_00000      = sum0_00138 +  ~I1f6540c5f037d861dee2c0091cba01ec +1;
assign wire_qout_00139_00000      = sum0_00139 +  ~I9632bb500b7faaaaeb649d74c21cbe8c +1;
assign wire_qout_00140_00000      = sum0_00140 +  ~Idd0217a35c3adc8abc7bb581a5df7a2d +1;
assign wire_qout_00141_00000      = sum0_00141 +  ~Ic05b46168884322644db4e331d37d759 +1;
assign wire_qout_00142_00000      = sum0_00142 +  ~I53c88dc237bb2cd02d50fd7f0a168a48 +1;
assign wire_qout_00143_00000      = sum0_00143 +  ~I7450d4ab3ef0227e93a02bfd620d047b +1;
assign wire_qout_00144_00000      = sum0_00144 +  ~I2b16e5b4e279bb29c3c675b72083e5fe +1;
assign wire_qout_00145_00000      = sum0_00145 +  ~I70c92e8ada46476d15ef4b3c620d2601 +1;
assign wire_qout_00146_00000      = sum0_00146 +  ~Ib193b07804d6d5f111b06bda487bfa5f +1;
assign wire_qout_00147_00000      = sum0_00147 +  ~I885433b0ab16c6d87abe45af13c9e529 +1;
assign wire_qout_00148_00000      = sum0_00148 +  ~I198c055930cb89d0390c336eda8fed4f +1;
assign wire_qout_00149_00000      = sum0_00149 +  ~I688a2c72e69b217d2673e8da75146a83 +1;
assign wire_qout_00150_00000      = sum0_00150 +  ~I3b6fde4ed14cd68af1468ae1d4cc1a22 +1;
assign wire_qout_00151_00000      = sum0_00151 +  ~I5d3df1e7563630311f56143ee6d97a8e +1;
assign wire_qout_00152_00000      = sum0_00152 +  ~I90a7ea789d3bf7f9126c786474a56da0 +1;
assign wire_qout_00153_00000      = sum0_00153 +  ~I5029424c9d9fe923eeb858b1e62cd758 +1;
assign wire_qout_00154_00000      = sum0_00154 +  ~I1e805c70d50c2765b4a03ad2982dc421 +1;
assign wire_qout_00155_00000      = sum0_00155 +  ~Iba58175a7fd5c5da650222193caff0b3 +1;
assign wire_qout_00156_00000      = sum0_00156 +  ~I7401a0501ba69c5559fbf00c77e58dc5 +1;
assign wire_qout_00157_00000      = sum0_00157 +  ~Idd9f7ea657ea9cdcb45a7e4b573b9d50 +1;
assign wire_qout_00158_00000      = sum0_00158 +  ~I53f275395dd6be17961a5edc3e8da7f2 +1;
assign wire_qout_00159_00000      = sum0_00159 +  ~Icab010d78cd66b02e089c74f04bf4e75 +1;
assign wire_qout_00160_00000      = sum0_00160 +  ~I376a48b7e0195a5aacc76a0ad8bd14b2 +1;
assign wire_qout_00161_00000      = sum0_00161 +  ~I241622b0367dde514f96ece55c8c3964 +1;
assign wire_qout_00162_00000      = sum0_00162 +  ~If94a1abfb972f63629d07e64dc23863c +1;
assign wire_qout_00163_00000      = sum0_00163 +  ~I07b9b1f4fa01b16cc69356057d3b6154 +1;
assign wire_qout_00164_00000      = sum0_00164 +  ~I2288a6ad3b748b716249f4adc42d52c4 +1;
assign wire_qout_00165_00000      = sum0_00165 +  ~I022df337bcc05ac5648b8ae2e42f3a76 +1;
assign wire_qout_00166_00000      = sum0_00166 +  ~I60d9a7f95fb8623753002ecaf9a4efcc +1;
assign wire_qout_00167_00000      = sum0_00167 +  ~I23a74ea5e7174d95e6d16a5e85ac236b +1;
assign wire_qout_00168_00000      = sum0_00168 +  ~Ie697d28d757df82b3901564bda43251c +1;
assign wire_qout_00169_00000      = sum0_00169 +  ~I8572aedc94f7243ce5eacb332c81eae2 +1;
assign wire_qout_00170_00000      = sum0_00170 +  ~I6734123aaf6320da75638b212812732f +1;
assign wire_qout_00171_00000      = sum0_00171 +  ~I7f6dc6f0f403c58f9aaaa70c2383a666 +1;
assign wire_qout_00172_00000      = sum0_00172 +  ~I66391978843c39b6acbdb4847a01050a +1;
assign wire_qout_00173_00000      = sum0_00173 +  ~I4f756e4125c8af5c412944b273e01cb0 +1;
assign wire_qout_00174_00000      = sum0_00174 +  ~Id2c9f7ac95de07148c54803f69347f56 +1;
assign wire_qout_00175_00000      = sum0_00175 +  ~I5061e13a179d27e1ba5f89ce8ee0fd4a +1;
assign wire_qout_00176_00000      = sum0_00176 +  ~I0f7c32fc1548fb49b8041f55c157498a +1;
assign wire_qout_00177_00000      = sum0_00177 +  ~I89ffab735ee30423c82e079ed98216c5 +1;
assign wire_qout_00178_00000      = sum0_00178 +  ~I9494921d8487ee0b314f75cf0380fd2f +1;
assign wire_qout_00179_00000      = sum0_00179 +  ~If2b3e7d1541cbd8ffc2b4cfc3ad13a57 +1;
assign wire_qout_00180_00000      = sum0_00180 +  ~Idf3d79da44f2d686f5bd43c3c1427430 +1;
assign wire_qout_00181_00000      = sum0_00181 +  ~If8125ad3c9e7f0a2b84106064d320996 +1;
assign wire_qout_00182_00000      = sum0_00182 +  ~Ic9018b88fa91fb638bbab0613795ae13 +1;
assign wire_qout_00183_00000      = sum0_00183 +  ~Iad4ea0196eb32f9a152c9e6fe5059e46 +1;
assign wire_qout_00184_00000      = sum0_00184 +  ~Ia8ff29ed728e7f2ae4213f00328b495d +1;
assign wire_qout_00185_00000      = sum0_00185 +  ~I70717726200ec02929f679ef05496455 +1;
assign wire_qout_00186_00000      = sum0_00186 +  ~Iaf1e4c7dae6ad89567836877c08f57d2 +1;
assign wire_qout_00187_00000      = sum0_00187 +  ~Icd09aa81e9b43528af73e23b2f0f80cb +1;
assign wire_qout_00188_00000      = sum0_00188 +  ~I6ebb2b94f0f80425f8401ae823d92a1d +1;
assign wire_qout_00189_00000      = sum0_00189 +  ~I4a2c3204a6a9936d4a215b46c0ffd045 +1;
assign wire_qout_00190_00000      = sum0_00190 +  ~Ib02c0694762c4815448b2c8d3df767c2 +1;
assign wire_qout_00191_00000      = sum0_00191 +  ~I98cee6efbbe565d3a4de16703189782f +1;
assign wire_qout_00192_00000      = sum0_00192 +  ~Ibf981c01a9d44cbea3c6d8ead92bc2ab +1;
assign wire_qout_00193_00000      = sum0_00193 +  ~I864c33e8ea204d20a9baef4584f22d4e +1;
assign wire_qout_00194_00000      = sum0_00194 +  ~I6ad3228e0e2e1f19648d73e83ba5a229 +1;
assign wire_qout_00195_00000      = sum0_00195 +  ~Ie099210a99a4899c53baf39559592690 +1;
assign wire_qout_00196_00000      = sum0_00196 +  ~Ieeec71d9df4613555fade2ced7b3baf1 +1;
assign wire_qout_00197_00000      = sum0_00197 +  ~I4931884e3544af182bcda9061091a42d +1;
assign wire_qout_00198_00000      = sum0_00198 +  ~Ib3fb10da528d450251764a9b9ede0dba +1;
assign wire_qout_00199_00000      = sum0_00199 +  ~Icdc9e676957b2223d60c413331fa982f +1;
assign wire_qout_00200_00000      = sum0_00200 +  ~I381f6051282c062ccf53866830344cd4 +1;
assign wire_qout_00201_00000      = sum0_00201 +  ~Icfc21935c007fbbceb2a67ebe1a68a0b +1;
assign wire_qout_00202_00000      = sum0_00202 +  ~I120d597a80158374726e064fb0f099fb +1;
assign wire_qout_00203_00000      = sum0_00203 +  ~I2520aa556aadf851f58f0b1820498730 +1;
assign wire_qout_00204_00000      = sum0_00204 +  ~I6203f49a08107f7185ebadeecf2c16b0 +1;
assign wire_qout_00205_00000      = sum0_00205 +  ~Ia706fb593b63cebbee0321c154cb859b +1;
assign wire_qout_00206_00000      = sum0_00206 +  ~Ia4b5f2b07556629673fc6576bc49a5dc +1;
assign wire_qout_00207_00000      = sum0_00207 +  ~Ic532c6b85b156f821e0742f47239a65c +1;









   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
            sgnprod_00000 <=  1'b0;
            I5033323484d90d6bfbe03749019fc6dd <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00001 <=  1'b0;
            If5dad13ac41b3034bdb034bc86c9b348 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00002 <=  1'b0;
            Iac428f9f798618e1ef495c626c41892b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00003 <=  1'b0;
            I5a6427c8f18b36d2ea18fe60a0831ef1 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00004 <=  1'b0;
            Icc29441eac6ca7a138d45743d37505e3 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00005 <=  1'b0;
            I0e7754dcbc04a4850e052ae4a2fbe328 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00006 <=  1'b0;
            Ia30c019ed8ce395556494a92e7b42a92 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00007 <=  1'b0;
            I9799695ea8244992a6694eaf5c8ae64d <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00008 <=  1'b0;
            I4524cd664b4cb41f642c675fa484c84b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00009 <=  1'b0;
            I64e959d80af111ed2fcd54a5407d21bf <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00010 <=  1'b0;
            I3e0da4bcbab4804b5397fb3aa2c94f51 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00011 <=  1'b0;
            I3740b30d31f3c61d93a14a46e3199c4d <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00012 <=  1'b0;
            Ibf0a30abfec9031737eada436ac1a0d4 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00013 <=  1'b0;
            Id36e8953a02400a5ab1f4dfdb0422e6d <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00014 <=  1'b0;
            Ica71108a53bfcfd1892b4d03ef68110c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00015 <=  1'b0;
            I7c97629ec6e594f9b2160815ddd133cc <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00016 <=  1'b0;
            I4823c8239ace86dc399e906c1b5a0d74 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00017 <=  1'b0;
            I10ad572ca72c2ea991487c39f7eabd7b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00018 <=  1'b0;
            Ie9f3fd3a6d16316e55addbe0e336519f <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00019 <=  1'b0;
            I07965bca84276dd56da1af98e64b0adc <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00020 <=  1'b0;
            Ic2ade31b8bcf68c4dcc1a371ff14074b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00021 <=  1'b0;
            Ic0edcf240048fbfde4e938c3e4c5e281 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00022 <=  1'b0;
            I8b42e89ff5f780d4ef8cd1cd5c99ef61 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00023 <=  1'b0;
            I70b1b8521b36920707e95fc9418eb8a9 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00024 <=  1'b0;
            I4fb1c32a62cbbaeb585c6564a3c938f9 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00025 <=  1'b0;
            Iefc37daeec14e14ef2fe0716f73109dc <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00026 <=  1'b0;
            Ibd15f164f6d2ac9e5721a21464bc2c5c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00027 <=  1'b0;
            I951dfff9507bb70214d48e03a0ebb3a7 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00028 <=  1'b0;
            Ie78e30b2a2eda75d0df7d10fd67b5e36 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00029 <=  1'b0;
            Ia0b83a372dd4115dc4d61eb8ff0811b9 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00030 <=  1'b0;
            If5c5bcbbea01aa22f242b913f0d01929 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00031 <=  1'b0;
            Iccba58cd3519fb4cc75a61b50da1d562 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00032 <=  1'b0;
            Ibc0999e4d0b3cc2650f9348b8c204b14 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00033 <=  1'b0;
            I2aeff1fb4b839a581acaf26f90f9113c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00034 <=  1'b0;
            I7d60d53f883f8187700c4e78b4c22f1c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00035 <=  1'b0;
            Id6fcf4b7af4a37c854a12e2ae80851fa <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00036 <=  1'b0;
            Ifa5e5f7d753964f14f0f16dbe552fd85 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00037 <=  1'b0;
            I900d471b087cf5a436c2ad66a84d8280 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00038 <=  1'b0;
            I6d1434907f0292ea2ee47cbc5b52bfb9 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00039 <=  1'b0;
            I938bef7ba7ae1739d8e6a6a7c117a1b1 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00040 <=  1'b0;
            I6384a9416b2d1da01df1b2d7b16c5390 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00041 <=  1'b0;
            I5097a79e7cf7a30d38ba198d1407119c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00042 <=  1'b0;
            Ib113c26c8dcf49c972c41a938059a787 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00043 <=  1'b0;
            I970c4a25a8bce82a9d2846679029fcab <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00044 <=  1'b0;
            Ibe2af096ad2db26e54d8b4b3bb05175c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00045 <=  1'b0;
            Ie48569c467fba0c1291f71d6080ebedc <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00046 <=  1'b0;
            I90e7ded06617b49cdb8b5301fe9c6a20 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00047 <=  1'b0;
            I4920014f5d017f4e840dc3b88526955f <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00048 <=  1'b0;
            I03b70553f1c501609400574ae7cd73f5 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00049 <=  1'b0;
            I63c9bf68b43ed66c51b0f4c0ed92e9ab <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00050 <=  1'b0;
            If408dfead07757878cc878131bc7d6a3 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00051 <=  1'b0;
            Ia0857d63d309807789b6ff4f6028f1b3 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00052 <=  1'b0;
            I53921b825c5e434b63bee0e1ecb7a517 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00053 <=  1'b0;
            I5e68f84e123c37f19a03c13892c77e19 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00054 <=  1'b0;
            Id5270b57c6fb4b18db3bbd0a523e467e <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00055 <=  1'b0;
            I3c18a84617eb21472d53e598700d7f4c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00056 <=  1'b0;
            Id36663e7a01fff3170833ecfecac1321 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00057 <=  1'b0;
            I8d3be15109c7007a79fecaac0d891626 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00058 <=  1'b0;
            I92169cc57291f20d336a479e392ec271 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00059 <=  1'b0;
            I6178b220b469b40dac39168057023a1c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00060 <=  1'b0;
            I55342938216a0ea0889f96c2f6c05ce5 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00061 <=  1'b0;
            Idf28431c76a84a48dd895979d2b11a63 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00062 <=  1'b0;
            I1ef61124c8d62e8f6a82a729fb091694 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00063 <=  1'b0;
            Ib8bb96f0372323e6a8072ca56fb9396d <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00064 <=  1'b0;
            I432f74dda4f6b1cebdf5ad59c659080b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00065 <=  1'b0;
            Idc689442305acd00f0f32416d8fb3773 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00066 <=  1'b0;
            Ida03738adc101c03c2229756bed2469d <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00067 <=  1'b0;
            I4d14c75f28f3e516c259ea288996131b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00068 <=  1'b0;
            I6e6cbbf430d57f347a0d70558af143d8 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00069 <=  1'b0;
            Ib7487df45118e44acec6b9d07bbd5969 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00070 <=  1'b0;
            I492f382fea500462b3d0866240fb91b2 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00071 <=  1'b0;
            I3fb3ebddaf28efb56092d19a1b4695de <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00072 <=  1'b0;
            I22a26b7f0b1c8c16b00597732ce2ab23 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00073 <=  1'b0;
            I2ac08a2d8c917ecb37fbaf5325cb0473 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00074 <=  1'b0;
            I50ff8f51e75fb9ce3db983c2a0f57196 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00075 <=  1'b0;
            I444bc340ffb7ef7b72d4d2e761d58872 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00076 <=  1'b0;
            I039c6cac5830759529595a958b7f65c9 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00077 <=  1'b0;
            I0584de7d919236ab138e288a27d08ff1 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00078 <=  1'b0;
            I086402c82ec67ae09a9e6360c58904b4 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00079 <=  1'b0;
            I1cefdc831c146187c77f861b3e2d1af0 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00080 <=  1'b0;
            Ida9c16ae57d17b6faee8a54838860447 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00081 <=  1'b0;
            Ia3b9fb112f39dd0ccbf7555659369efb <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00082 <=  1'b0;
            Ib1bfcdc0c972aafc99116ed8c0511445 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00083 <=  1'b0;
            I7adff505c50450a04f1717cac1adebe7 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00084 <=  1'b0;
            I699feb4382974a02b21cb387c13f7f3f <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00085 <=  1'b0;
            Idc99c3b23e49aca3c98f0685ea34441c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00086 <=  1'b0;
            Ib67318fa6954ec8f3247927d34e74f8c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00087 <=  1'b0;
            I8774ce3f11362915c4331d1026e452dd <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00088 <=  1'b0;
            I2392b2d17ffed6073875fbe8e92534cf <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00089 <=  1'b0;
            I3a4f0d3e32596ef05477f494768d4266 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00090 <=  1'b0;
            Icd08ff59cf6be3ba97698dd55703339e <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00091 <=  1'b0;
            I985fb7ed22a8476ea322c9e3c2b3851c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00092 <=  1'b0;
            Ib985709316b1b0a9d3fa3c1eaf6c641f <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00093 <=  1'b0;
            I4be898887dff6e2cebe53f135ece131b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00094 <=  1'b0;
            I004db04f61fb57aba81e15cc015442b3 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00095 <=  1'b0;
            I8f7e3dfb2f728d4cd1e79b82b62b0406 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00096 <=  1'b0;
            I991054370345e61638ddaf81785505bd <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00097 <=  1'b0;
            Ifa1f503965270d10e7a5c9a15576069b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00098 <=  1'b0;
            I24f773842a4742fb58d09cae45717b2f <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00099 <=  1'b0;
            I5bac7e0d778a547a0ae764fe259b6f7a <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00100 <=  1'b0;
            I255577ebee6768871df0224fc1db2db3 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00101 <=  1'b0;
            Ia7fb4af3d3529a32f902a52cf5598474 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00102 <=  1'b0;
            I2c98806141f064c9e92935b23a84ede1 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00103 <=  1'b0;
            I5680847bc8d224fa4ed93b2fc0d841e1 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00104 <=  1'b0;
            I365254279ebb10dd7ba0b3482d5e34cd <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00105 <=  1'b0;
            I57bf4ad773cc058ae1bb7b1911dc3174 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00106 <=  1'b0;
            I57072dfb29c4a3d2e2b40e46e62f0d95 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00107 <=  1'b0;
            Id8cafb6f76321bdaba9711133be7be99 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00108 <=  1'b0;
            I6344e71ca2b0fd39d36caedd889c3085 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00109 <=  1'b0;
            I0c99a68e0bed90afce18807acf7d55bb <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00110 <=  1'b0;
            I1c95650979c86310ae2a949961c9db11 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00111 <=  1'b0;
            I04eaefa5d133e53494fc270b07be7043 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00112 <=  1'b0;
            I4a64fa2412eb8058c2dfd9351d7b297d <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00113 <=  1'b0;
            Ie8bb2fcb752c6a33254963d1ebb4130d <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00114 <=  1'b0;
            Iac05b7e3ae18f948b72c356ccfb8000f <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00115 <=  1'b0;
            I27da3f75cca6c49e55db90306aa68e94 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00116 <=  1'b0;
            Idc7fed723190098341225fe01ba65ced <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00117 <=  1'b0;
            Ife9065805598960919ee4f14c3cc6fd4 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00118 <=  1'b0;
            I717c5c2d6a2be61593492ae5f17a112f <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00119 <=  1'b0;
            I4c31fa8e6eb648439cdae1de1afe0d6f <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00120 <=  1'b0;
            Iead549a9af27f1fced7d9c36e7b5c3f5 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00121 <=  1'b0;
            I10422eb79364e7d0e21e1643d9060331 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00122 <=  1'b0;
            I914cb87eba8baa40cd515334e59f26b2 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00123 <=  1'b0;
            I32ed679af4ab759901aee43c9d93eb67 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00124 <=  1'b0;
            Id376dfa5141402f4d41a8858180ed87e <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00125 <=  1'b0;
            I98a384bc62ee03f5ad7df20ef2d9af95 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00126 <=  1'b0;
            Icfed259ca2bb2732d8e0c26ef67cd4cf <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00127 <=  1'b0;
            I20861535c450d6e6bf11c45dac120454 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00128 <=  1'b0;
            I013929385ad819ddfcfcc59c22902ee3 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00129 <=  1'b0;
            I34fffcb07fe82f11fe142f7c37f39155 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00130 <=  1'b0;
            I61ca60fde05ed88cce714dcd8c13b827 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00131 <=  1'b0;
            I4907dd45c158dc7e0041c64f1fb388f6 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00132 <=  1'b0;
            I2c8f6a9b9f655b317bb0af4d60fdbc4b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00133 <=  1'b0;
            Ic7dff631559304ec59f0696c66436d62 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00134 <=  1'b0;
            I6a239d3e55b4a9a3be9989a85bbec545 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00135 <=  1'b0;
            I630f905e55f08e7d1569a08e937ad216 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00136 <=  1'b0;
            I8d13eb3669785c4279c685763d4f3fad <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00137 <=  1'b0;
            I25a6f3de9a9a01cbbdd32ed848561aa4 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00138 <=  1'b0;
            Iba3dd4b2c2c85c4cfe770d9b52ef4634 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00139 <=  1'b0;
            Ie1b744387b5200a504e4874e14d2f282 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00140 <=  1'b0;
            Icf76cb69aedf4db01cd3444f4c4ba471 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00141 <=  1'b0;
            I4857b5b50556c8e7fff4b2d3e08e4b28 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00142 <=  1'b0;
            I0a1e9cf99f1d4725327615f50fcc3ad0 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00143 <=  1'b0;
            Ie844f4c446983ce381b0bc4c0e8ef7d7 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00144 <=  1'b0;
            I6067f47cccceea96ac46ff0d457b25f2 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00145 <=  1'b0;
            Ifd6fd1f3cbf8884ca7f64bc42278e4fa <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00146 <=  1'b0;
            Iaec9fd9e79371676bfa8ff14b4feae52 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00147 <=  1'b0;
            I500757c4eda5d3d899aee47b87da585b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00148 <=  1'b0;
            I47bf091b0fa74ad511a760bad9d2506c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00149 <=  1'b0;
            Ia4c3d0cd9957f678880de5775de76e0d <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00150 <=  1'b0;
            If5f957fa2f055b1c2c28e8d7cfe3e9ad <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00151 <=  1'b0;
            I3608378a5da8c66bef58528d56192530 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00152 <=  1'b0;
            Ie6dead855e00ea0a8e6a9b7503aaebb8 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00153 <=  1'b0;
            I3bae5e6862e003a8b9a476f72cc6858b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00154 <=  1'b0;
            I4431adecba8be9e5f21bc6b3e1f8cb10 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00155 <=  1'b0;
            I21c7a2885126d532d00484376588a469 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00156 <=  1'b0;
            I2c4d7339ff2fe68d060dd8d961dcab8c <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00157 <=  1'b0;
            Iee518b15b067eec58cccfa37f7432ea5 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00158 <=  1'b0;
            I42145be9c2a80288ba4a2edd91f661a3 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00159 <=  1'b0;
            I9dc297ad41fafcda77f5347f331cfc25 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00160 <=  1'b0;
            I846700c79f30ca954cc2933fc94d355b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00161 <=  1'b0;
            I8af96a91457316e49e3f7dd5e57c82da <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00162 <=  1'b0;
            I7d1c247500d7d32e406b2a5f7e2b745b <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00163 <=  1'b0;
            I66d85c030a8864505298919046056305 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00164 <=  1'b0;
            I4841257ae596d9d3e4eb1e6f886956b0 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00165 <=  1'b0;
            Icd6f7ec117f9ab4eda8c5eba41386ffa <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00166 <=  1'b0;
            Ibc0498839d1d9b6dc853b8e5d7a88fa3 <= {MAX_SUM_WDTH_L{1'b0}};
            sgnprod_00167 <=  1'b0;
            I142ebca7f155e287e38ddf45423ab0fd <= {MAX_SUM_WDTH_L{1'b0}};
       end else begin
          sgnprod_00000 <=
            I5b177dd5c14ad082516b47f550875682 ^
            I477326720157df2503149125a43ee987 ^
            I319012bc6fe93d78de57bcace0caaef5 ^
            I174b6c36f2af82f8047cc76543a3b4ee ^
            I8fd5787ebf758919e7cb75d7419441e8 ^
            I413b1c1985a6c9c6f202e85ff901e3a8 ^
            Iea3e35ece9fdb3aff3b9ff5369e9a7e0 ^
            I30c0fcd89e0cc7c5fa348df7b4fa2ccf ^
            exp_syn[0];
          sgnprod_00001 <=
            I77b05a8aa92c66a235195a66dc13c0cc ^
            I876fdba97e755b74532f7ab191fbac14 ^
            I5590d801fd7fb496019d4c31b7c6d898 ^
            I25f1ee9cee4d04bd8fec1fe601d016d7 ^
            Ifebcf64858d5e2d07ad7894d6182eb11 ^
            I163cf58b9a308e0439a8dc7c1526e6b5 ^
            I3347717ba9556e69de30ce7533d4f5a4 ^
            I5f96a68d20e3ebc71dad4b43305baa20 ^
            exp_syn[1];
          sgnprod_00002 <=
            Ie117f6ec475f5d6444998af151ce4e69 ^
            Ia538dadbd6ae3711740595a18c89b65d ^
            I141cda06bae0c5666e3bc61c6fe5ad66 ^
            Ifb70a30f8bade95f402e71f95fe6644b ^
            Ie50aca688b3433fad7565998cb900155 ^
            Ied33f18cbb778d5ba744d249f91c950b ^
            Ibe97860165dc5d9a076ebd935385ae51 ^
            Ie46b71f55aef4d00168202431d47dce0 ^
            exp_syn[2];
          sgnprod_00003 <=
            I92cb615e2c439914e72ce001256518e4 ^
            I7d6a6026eb3c4d06e682523424f9628f ^
            I06ad520cb02e46d34c45f207d42a9243 ^
            Ifa3df8b249467cc1e827c69925ef415f ^
            I4ba41864bb1d2130c6971e0b2903027a ^
            Ia67f9b902a21de0414eb8dda52171991 ^
            Idbbf2ce4a30787c5f07c3b908a73da75 ^
            I71d3a999d88e591e102398409b3adebf ^
            exp_syn[3];
          sgnprod_00004 <=
            If7f3174da35dd39af7f4792aaa649bf1 ^
            I953b975a89adcc88039284970e9b3404 ^
            I5a247475beb737d470f03507e55f5b24 ^
            I93084ccf5b5e4efaee968b497bb2a775 ^
            Ibab55499323660588ec82ebd07ab0572 ^
            If9285bf7611bcc5ea6432215c349e021 ^
            I3566033cf5c9a06977c9182925750707 ^
            I87b10521099179c18652c86d5887c908 ^
            I13a98f98c54b2e412cd88c96f016c41b ^
            I6f7a45fe64ffeda9ed120be3a4519aea ^
            exp_syn[4];
          sgnprod_00005 <=
            Iad799775eb657f8973e6dfcf70a9875c ^
            I5ec1e530b9007a75a778af4d82ab427b ^
            Idd59a5357d4c835379ed180ac0924bf1 ^
            I7a626ec321bf963a5401892a7e3891c7 ^
            I3342fe0c5d3ee5021892d53eb45bde21 ^
            Ia858ff5551286beffd4cf82f876d30ac ^
            I5402fd208dc7ca81dfd2920a9cfa2715 ^
            Ic32c6734132776c290155a80025fe366 ^
            I5d92fdff96b9cd64f3af2b28b13e9956 ^
            I221524a69e18854f029cad30e8f94e8a ^
            exp_syn[5];
          sgnprod_00006 <=
            I55e4ad2d71a29ad63b4999d64ac0dc4f ^
            I592a495aecc800236c3470ff8e6adbb5 ^
            Ifdb5589982db805a0416e1c01276249a ^
            I0c47ccef4b55410286248884a7249703 ^
            Ib68deeb7bec4ca3585d1a4dcbf8793f1 ^
            Ia17906696bd0e095d7a5297da2e049ea ^
            Ic11a6b77b84c44180eb99220a0c4c9f6 ^
            Ie08ad9bd71329858c1742c8f571a1c36 ^
            I8c0c1a0a35f4f7a688f516c567242d39 ^
            Ib105151d91678f81978495ff94b1e651 ^
            exp_syn[6];
          sgnprod_00007 <=
            Ie92110d19f4886cdfcfacd0920c06a4e ^
            Icf3ad912aaeaa0c5cd1ab0edb898d6e8 ^
            I857d3155df0b6dd704514b039c66fa97 ^
            I3bc094d67805664859fdcb66f1360e64 ^
            Id14074d5230885c38b89b09b130ecf68 ^
            Ibf312ae4f51fbc44b43848f9df62a45f ^
            If6ce2fa9f0b8bc74442ed8262b5089cf ^
            Ibabf61085ca7af8dfc7927b3656a76f7 ^
            Iebecd2d19f9174d87deedc1a273e7baa ^
            I94a9de743d5bedbea3876de954f479bd ^
            exp_syn[7];
          sgnprod_00008 <=
            I59c5da6338f431a626c86a065a355c35 ^
            I8edf1a08ef943f06ee28771c6e140e28 ^
            I1c8024aa9d81704d2dcf63e34853f8cf ^
            Idc1b8aa2f81a7fbd87e4f5821d14bf01 ^
            I02812a8a833bb69eb168a1004b6fafdf ^
            Ic44eab478be232721e7a43d14beca32f ^
            Id1dafb7e45b860d506e0c2c91b28142e ^
            I9db50007841762c9a10f6b7e9d40f858 ^
            exp_syn[8];
          sgnprod_00009 <=
            I36ba87b69b5b9dd919319230f697dfad ^
            Ie7d9730b191781c78391141d95d4f8bd ^
            Ib774f380e3d7cfd1f5f064e93d8134b4 ^
            I13b0c9578f7b6b3b7e6704d7b44079c4 ^
            Ia01c82761aeb124cd92fb15ee367ee8b ^
            I2db290170ddae8dc52ce07edaf48b365 ^
            Ied764ee7730ad129b6f62837ef50774a ^
            Idc5dd6caa4ed17a63746d30d381a944e ^
            exp_syn[9];
          sgnprod_00010 <=
            I719a892ad54e63b217c7271741b29cc5 ^
            Ia0c192e590d8c914555b434ce5a634a8 ^
            If2b40d249c531e10cc22d1335f350441 ^
            Ibe7e5c2cb9c50eca34a3859d13e83a92 ^
            If0970d9f7b053fce3ced3521b4885588 ^
            I777ee54ff20d0544af18ad8a870d6915 ^
            I4edd64d1f1da865b1eb886e22726a033 ^
            I4dbabfd592b74aef93b819163130ef5e ^
            exp_syn[10];
          sgnprod_00011 <=
            Ifb064c69c7110c014593149ae69c75fb ^
            I2c741a5fed7d88e9bdd6b7459feac649 ^
            I8a9e516aa824260998d10db758642bb0 ^
            I8bb5522183b65583fda83067990b3e94 ^
            Ib0001d7298ad1f3b1c7603173a70d8b5 ^
            Ibc9a860879ccc58c815b9f6caa23320a ^
            I17c9d8f658dd6b2916b645d103f4702a ^
            Iba283e99a57d0a3b78ad2e309c316b65 ^
            exp_syn[11];
          sgnprod_00012 <=
            Ic98c8641d2022080297c54ff2539e75d ^
            Ia9c273b32d0701c7f185ab2de9e57829 ^
            Ibf5c141c5cc0a6a20c05b52bf8282476 ^
            I2518ccf385b3b677d95983bc550282e8 ^
            I86fefad34d3c864dd0e725133f303b4f ^
            I180d4f3b23b518271d7cb8189fbeadc5 ^
            Ic7ebdc317c978eb275eca41d5b9106a5 ^
            I84057a3b319ab3d6a2ed8f2310f970fc ^
            Ifab075b1437495268b6a3be4cb022e71 ^
            I89c5af1a6176cefa1f77ee69996473cb ^
            exp_syn[12];
          sgnprod_00013 <=
            I17a6511072c7fb4846be5844decf17d6 ^
            I9d18ff3465afd8cae63abba68487542e ^
            I1e77fe6aeaba852aba34ed37dd53add6 ^
            Id38852415486e6989b89a0d85ad6771b ^
            I89af7644c48a80d7d22f50b008d35841 ^
            Icfc03646b36b971b9fa57d04a26dbfc4 ^
            I05e739fc87e962848f265e2c73338cac ^
            I624958486d181501c7a8ec2642cb503c ^
            Idd775d9fe6fa8dbdbfb07d4071b9caa5 ^
            I17086dc5193aa55e5c6f56ecd365cc00 ^
            exp_syn[13];
          sgnprod_00014 <=
            I7e12ad8a8ef857e02f4563b2f3a7f0ca ^
            Ibb35bace971548c9fc98d773d1aff712 ^
            I68b585571699a57bc6ba5e8955467119 ^
            If76f04fe0baf171d7df2c0cd849aea2b ^
            I5134b762ac428bed07ce102d8927a418 ^
            Id277f5f05551eeb5dec1701056330da1 ^
            Ie886c5effc85f1fe0b6411db4a2cde77 ^
            I3c10d579f80bd0106506ad047d75f188 ^
            Id18c5a1d4eaa73a94e699e5f9e3c3d35 ^
            I9ece87047aec25abc02a5eea72f0e647 ^
            exp_syn[14];
          sgnprod_00015 <=
            I12f2f886517647044cc251861721bbb9 ^
            I27e1d2e0e980216b27b90ea48c061025 ^
            I41eff06fe1dea8be4613945de596d3ca ^
            I94e4041b482064334fd0ed92b91bde89 ^
            Ida3d808d100e0bba290f96ed9e744e65 ^
            I4c66570630a650fa7b9bec543f685487 ^
            Ib1a40247057324b0bd810c844bf11f51 ^
            Iddc5b5b4501f9f13bcaf22081e5a70f4 ^
            Ia71cf07b645c58cffe33be1a9a960eb2 ^
            Ifba3e46933049cb093d2c1809f3a8a3e ^
            exp_syn[15];
          sgnprod_00016 <=
            I4acf6d84471cd237f65c9b2391b7a20c ^
            I17b3a9df6752da6cc987e902e6bbad48 ^
            I168afc1863f909dbcb6a9230db9f3e00 ^
            I989dda9add29306d7b3c0f376822763a ^
            exp_syn[16];
          sgnprod_00017 <=
            I7f7b30f2acbb8e31f50b58096b738254 ^
            I615053b36a1851a06125e2ed5ec7f880 ^
            I9890f7fc708c7b8cf460849b4a30025b ^
            Ibc929201e2eeb3e61cc8f0acbade497a ^
            exp_syn[17];
          sgnprod_00018 <=
            Ia098bbeda8b755ece6b88eac83d03e55 ^
            I87f34821cd0b58f8855b25c75f2dd32d ^
            Iab2f643f81921ed8464e1bbd9fa8c68e ^
            Ib0dfbbbca2d3d264065f73b4241caed5 ^
            exp_syn[18];
          sgnprod_00019 <=
            Id20e72ac258d1d1b6cdca1e6c9e3596d ^
            I5ebc3047985651f4b9a957d502a97e95 ^
            I53222c82827cab7c770e057ae91bc10e ^
            I339786aa60d4c71d12c65db27ac420fe ^
            exp_syn[19];
          sgnprod_00020 <=
            I7a387a1f887c32e9d0f8e89912a8618c ^
            Ifa09fc1b009d073d5a9973b430c63469 ^
            Ia9c8cc5e3becf3d48feedec8fa2c93a4 ^
            I4f134c0669b5a6a8c7e03be7eee30c6c ^
            I1c4b29e48d0effac4839037ae5688334 ^
            I3ade020bbdf8f954821f737439513043 ^
            exp_syn[20];
          sgnprod_00021 <=
            Iefe4099ff7e457f6b9fefc83e176c1a0 ^
            I487496233a32f657171b3789590d0522 ^
            I39d3bce4060032a81e6b6a1c1805cfe8 ^
            I9963d0b24763ed8038b1f3922b8f9548 ^
            I5e69e930a318dcb0594a823b3129d650 ^
            Ia50526cd3a3174bebc5a7a0889fda661 ^
            exp_syn[21];
          sgnprod_00022 <=
            Ie7470dd75b54d14038de19e4d3043ba9 ^
            Ifbc6aa14cd448bbe416897a3671ba857 ^
            I7547c56b32513ad45d775b4502596d9d ^
            If10f33385e236eaba56cbab8c2883399 ^
            I17d7f36fdade16dbcf621fe302bd7e57 ^
            Ie9f37dba0791359bc426a73639ce33ad ^
            exp_syn[22];
          sgnprod_00023 <=
            Ifc34f5d6b7a7d0533439794958959856 ^
            I87211ac14d832ad3205d47fb83cf256a ^
            I17cf58ef5326978c62c03c56090a299f ^
            Id79636d195efff260c430978f0bcee9c ^
            I8015717cd36aabbf2cf4aa3a5c234690 ^
            I9518532a8617fc8290eb6a5e981dea94 ^
            exp_syn[23];
          sgnprod_00024 <=
            Ib862ac63c230ccde7fae0e62f9d047fe ^
            I013d84bfd582acc7accf07ec522961fa ^
            I7cb58e4c486e683faa4acad4756815d5 ^
            I67d57e38df8cb35ca686ac2eb44e233e ^
            Ic0c13c9a929c8c46e8702cef74de8955 ^
            If66524125bfde5aa48ac70c4e448b38f ^
            exp_syn[24];
          sgnprod_00025 <=
            Icddb43f9b760a4597a0bb637fb405616 ^
            Ie41ca18c7d11a47e274f9c33f75393ec ^
            Idbf4ad11ab2a27044193448c8739fec6 ^
            I04864c28351edb33b61a103add6fb875 ^
            I431fc2e9533012c8571d8158d4777dea ^
            Ic3ec6375998b05a3e48f6c5fe7b3910b ^
            exp_syn[25];
          sgnprod_00026 <=
            Ie95662d4faf6b5a4cd5ecfa41697b983 ^
            If3b77c41fabcdb283f2c6fdacaa5e9a4 ^
            I6c765e677f42fe600b848698c8a78349 ^
            Ieca2767ac27170058499d83016447aa7 ^
            I403303228c0df825f67436f4a7e64061 ^
            I0ac421af6e311b6005c3e02e93ff94ce ^
            exp_syn[26];
          sgnprod_00027 <=
            I849ee5d34760be03d4285185136aa52e ^
            Ifb422c30663eb4824caa72326b238df6 ^
            Ia98de3691917dfb63bebdc3f8655c8be ^
            I67f87fbb746dd937fffc534c596f36c4 ^
            I23afd747ecece714e32fbb896b5c022a ^
            Ib9db80f43718305a8a8774d8d80c86c9 ^
            exp_syn[27];
          sgnprod_00028 <=
            Ie6212a29c7c6b035cfff4c869f945b68 ^
            I41ab6fb6ec6ef7ffff70e50f25f217b6 ^
            I0bce960fcc58938e6a1e01b912eabbf2 ^
            Ief72606c77113ae37845e4aa4a2ae5e7 ^
            I5ede62333e0f7ddc5446b653ba9a2382 ^
            I3b775b06b5d78fcd7373c966a62f44ad ^
            exp_syn[28];
          sgnprod_00029 <=
            Ie34534dfd435b3d1cf35e82ca71e83ba ^
            I0ec27b590ee6dcdd9c1086105e3b6c23 ^
            I452e51cca9acec44e36e4efd21b43034 ^
            I946246be5b4745508b7d4b578f83aaa2 ^
            Ib2fe0f68044c11f879e512a200f8099e ^
            If2372a5956f21f97eeb9c76281b6675e ^
            exp_syn[29];
          sgnprod_00030 <=
            Ie596289582a73e37f78f4ca4cab21e3c ^
            I7b80b4902fe98c10dd72c9eb082346e5 ^
            I3051f561a5e1131ebf167cb6ccb5adf4 ^
            I388528eaf83566cc56b23485a9c05962 ^
            I3ed6426fbdba8aaf1c948cca7442b3a6 ^
            I7b32c2b108e24750e2a24785668af3ea ^
            exp_syn[30];
          sgnprod_00031 <=
            Ib81431cfb3b281555fa7e5b4582a2524 ^
            Ie5373b01a92f2ff85be8077cfef2175a ^
            I284b23051c85300c2a1e3afe8f25e99e ^
            I71d7f72d83b7410de31e09ea96adb95c ^
            I4af3e2bf2ebc913ac902b48da672c5b6 ^
            I8ec99197a7d823f5745d382c10161430 ^
            exp_syn[31];
          sgnprod_00032 <=
            Ia3559d98eb372b7307f30ad1f7c4c7cd ^
            I0e8679271ba733bb87c44b6b9f0b6ed2 ^
            Ia7c9c24f8e993526e76c6915e56908c4 ^
            Ib895fec0b3756932b85962c1d129a03e ^
            exp_syn[32];
          sgnprod_00033 <=
            I8f1a8a22637d37c3692e808d5eb3d543 ^
            Ifad8c7bacf72583f91be27fbe5b7a1e1 ^
            I384e50fa8daa639124f083dda56fac00 ^
            I76aab345d13c6678fe37a4a7133cfd7d ^
            exp_syn[33];
          sgnprod_00034 <=
            Ic76e72b434b47c10ebac3fac4ea50bde ^
            I835b902949c2c4c09b757d4d35574a76 ^
            I5f1609647f1e71cef4ba2d605c6c8445 ^
            Ib4f368fa3d3ec11d9ffb2ae9a2ae6310 ^
            exp_syn[34];
          sgnprod_00035 <=
            Ia1b617e3d141263b51e58c5ef0bd7a89 ^
            If343015b4815b01dae88bbb6f2017b3d ^
            Ic98f33c6a4613534bcc9b6bc4b4f2d17 ^
            Idd0f3cfc5599481c954a2bfe69f044e5 ^
            exp_syn[35];
          sgnprod_00036 <=
            Ie74c72742807ae4243748fd27d80d626 ^
            Ied8bd4b6fd0e4fbcced6d20eb7435f55 ^
            I6cbc06919b9c695d99621db6f8d768cb ^
            I641539560711ff1824bd90baa0f21f96 ^
            Ie624c4dad5036a25ca314b94cf3c4b95 ^
            exp_syn[36];
          sgnprod_00037 <=
            I8510240df7dc41f85ad58a39868a1fd7 ^
            Ibe3d3e6bc58efc2e9d9eb1f96cdfe424 ^
            I72939e49bf2d9c6a84e404419fc644a1 ^
            I95f0acd4f955058041c035789c3a4d99 ^
            Ibf4b3caa5655cfb6663f9b7e2383bbbf ^
            exp_syn[37];
          sgnprod_00038 <=
            Ia0116a3cebf94318ed5b287960957ad6 ^
            Iaaaf373f7e6f55214915b93da9bd71d3 ^
            I0ceb14ac0187d804f9692e0c55b8e941 ^
            Iea424dd9d8916c4951b8746408b8a521 ^
            I049d1c09c15def12ba7bae95fc1c3d55 ^
            exp_syn[38];
          sgnprod_00039 <=
            Ic14760b65c6fe150c3c48e64389a41d8 ^
            Ibab1d13cd6a4f7b0c79c9f845339e53f ^
            I2919272e9ae3996a3e1d602ff72ba86d ^
            I1db4ea6916125702e7fb09d0f742e60a ^
            Ide06ba186ddb179b489ba6e3e209e3e8 ^
            exp_syn[39];
          sgnprod_00040 <=
            I6f420c64640dfb0c001f57df7e3b4504 ^
            Id75c23e80cdf25d883806ed20d4ae783 ^
            I4d4901ff372f6820ca9c8c29cefa664a ^
            Ice0234f25de4ab1f03a3cb01a2d61dbf ^
            I1b78785ebe2e7f77a3125a6334c4dc54 ^
            exp_syn[40];
          sgnprod_00041 <=
            I9eb87e62d23bc87d7cd82c0f329f247f ^
            Ied6c684cdd280b41ffab93a026d27282 ^
            I1ca188bcdebbf41d84f7a5220bd1d195 ^
            I9322a2a61900943075bbc23c72a3f65d ^
            Ie79c93f1703121713fb9401617f349a8 ^
            exp_syn[41];
          sgnprod_00042 <=
            If9a5d830e3ade0fd96b98f5949f165f0 ^
            Ie7a68c2b368a295f95571bc4a109b9f1 ^
            I0152dc6e6a7acd72a2144623e63998ef ^
            I9b560d9baf8a7422b0dd84720e924ced ^
            Icf25f076eec2bf81c899c66f6cfbebc0 ^
            exp_syn[42];
          sgnprod_00043 <=
            I7332e088bbff69db19c62685e033d26a ^
            I1b6abc8fbab3849b285e9f88a4fe867b ^
            Ic14f948884da19a272a4760ffaab9ea9 ^
            Ice5f7168aeb940d48093cc9df7cba36b ^
            Ic5c837a0556d1cb66edbf0294d08283a ^
            exp_syn[43];
          sgnprod_00044 <=
            I3600031716c2b4e21c9f577d34e033dc ^
            I859d795a7d141eb777c1f3c038203794 ^
            Ib9c194ec16f435a9357cb344cf25bdcc ^
            I69d82ab774d52c219509e993e7cc4deb ^
            I51ff4bda38746682e3cd4c68118c3216 ^
            exp_syn[44];
          sgnprod_00045 <=
            I2eac5b39c6f485c9ae0bd341f894633d ^
            I12a18a1f8d4416e9bc8abee6ac3dacfc ^
            I45bdd0cfe107da0d57cad1333bf95e3b ^
            I768720af835b02a8dab376ef23d17a15 ^
            I1c074a53e6c0f2467bcdd7c952f51670 ^
            exp_syn[45];
          sgnprod_00046 <=
            Id3de87169c440f95d406693ef77cacd6 ^
            Iedc463e359dd3003d9f7e50f3e858e93 ^
            I23955b54e486f0f0d21a2809a9472b86 ^
            I24075f37c6bbd90c83370de1a2e58af2 ^
            I37c49c5a2af240496f5a5706b0d42ea6 ^
            exp_syn[46];
          sgnprod_00047 <=
            I44daa5992b00e7af19adbee70bf01f2b ^
            I457ae11ad90c8478751eb4b42764e158 ^
            Ida3dd5e990ce3c237e9628a9a090901e ^
            Ifbadefd3a7ab50719a703400ddd742c6 ^
            Ia94c439131e1df5c95fc8ad3cfdba473 ^
            exp_syn[47];
          sgnprod_00048 <=
            Id88a7edf897eea1b4a137141789a04f5 ^
            I70dd1350d65155ee7b562f4c79024a3d ^
            Idc445d3f5b3b62562b0ac83e5f17e92a ^
            I723a6fee3b2496f23c48b3584f8bf9ce ^
            exp_syn[48];
          sgnprod_00049 <=
            Ied638fee34f8baed4154b0b72e43a21e ^
            Ief03713f5cf37200373a20d42c7fc9eb ^
            I3ac0799861144b599995318bdade2114 ^
            I648b62fa0bc2185c1756ee531e8e34de ^
            exp_syn[49];
          sgnprod_00050 <=
            I1b43f29e0ddb72467befd6f3a9c1c829 ^
            Ic07c650e6e49892a41cfaf3a37471426 ^
            I4082b3564c1949a19ed35bd5a88e1ef4 ^
            Ife631f9a3c4c64a3d92aa9586ae75f3c ^
            exp_syn[50];
          sgnprod_00051 <=
            Id0f4dbb72da33748d8baf723c5a32567 ^
            I44ccc3ae897109dd51f9afeef93daca4 ^
            I73bbf90b625d56f663ad10f9d21d8e76 ^
            Iaac1d82f0846fce1bd88ebf8e60300ac ^
            exp_syn[51];
          sgnprod_00052 <=
            I002820a37fa7c6c504c487df4368e2cf ^
            Ib0bb71b1f8829347b3a9a7543f9dd964 ^
            I1dd4671765f8826c2fe20c592c5e32c8 ^
            I3175159add7b814df637c2db8feb43f6 ^
            I48cd09f035f668536cd288a23010b07b ^
            exp_syn[52];
          sgnprod_00053 <=
            I76992221b1edff5684c482df7ac4693d ^
            Ib13436ad16a37d656d6b1ee95b9aee20 ^
            I47b0847946b0e00961233ac0101fa2a7 ^
            If2042aede3390bd208a281f0380c95a4 ^
            I119b2e5c2fea5338244c4019884af26f ^
            exp_syn[53];
          sgnprod_00054 <=
            I3751f191f5009322acb7c9be4f8d7129 ^
            I14fa7aebb608d4a3d67176ba27d34d9a ^
            I7b813d83b13bb7bc13940cf5714c06ba ^
            I0eaa22f5eca8f33dd254fe241017a098 ^
            I2bd34b2fd12f12bc301fd0d5d69c0fb6 ^
            exp_syn[54];
          sgnprod_00055 <=
            Ie517386cb5832e406fefc5e85eb2e7d1 ^
            I3fd0fa3b774d30a267d61e9427d09f3f ^
            I4ee312036de8c08300c358edcff1e1e9 ^
            I1d98943b01a6a2d8c4db18b98dd62f5c ^
            Ib715b1e0061b84ce614a30d961a83e7e ^
            exp_syn[55];
          sgnprod_00056 <=
            Idc07dc30c0a957e474546ac7a60df38f ^
            Ifc640243288c9b37b7eb9e00351b23f0 ^
            Ie83fa8157a7cce44c2e25f46ce897dbb ^
            I570c036d0237c53bb069c52d621e539e ^
            Ief8c2838abac83370fd7ec25c06d509b ^
            exp_syn[56];
          sgnprod_00057 <=
            Iad90879acba3fc2101829549264960f3 ^
            I951dedd7af44c3865a8f36888432d0c9 ^
            Ia7606050c683ecefc510ba92ac539a9c ^
            Id3b089fb6edd5bcfdbca142fddd5ff89 ^
            I561d79eb079915c0b1732cbddb119c2d ^
            exp_syn[57];
          sgnprod_00058 <=
            I2eb08ebaa07a1004638cdd61a7209b7d ^
            I46e1047bca2b38e62b4de80d1d2249de ^
            I41796b587316c600bf583edc62649bd8 ^
            I0a569f6536789efb7ad2377c11842830 ^
            I8bb75bf828d5ef337fa6a965808e4638 ^
            exp_syn[58];
          sgnprod_00059 <=
            I47cbb92d2284aef7b9e56e88f0ba6f7e ^
            Ib99e1b93fb7fbda260d93eea3d24c3e9 ^
            Iee6e52d75c093a24eb4e5e0b45feb256 ^
            I19b73c5c93a71e90f620572f23f0e6d2 ^
            I11ba339c8250d07b497c88a39a6df1ac ^
            exp_syn[59];
          sgnprod_00060 <=
            I8a4c1f23212ff846400651b100add502 ^
            Ief18a19d451f05f6051e3cc8de16d73c ^
            I7009c18515dd43d8dd2e5d1ee6779641 ^
            I173aa69cf52114e223ac1410d90b4bfe ^
            exp_syn[60];
          sgnprod_00061 <=
            Iada5bc4a51dc1bf57bb9cca11326bdff ^
            Ib6fbe376477afa58bfcc17a8564f78b2 ^
            Id48fe0672aa98f987162931527e9f9bc ^
            Ia4e89e99acb95f4183474b94798ca35d ^
            exp_syn[61];
          sgnprod_00062 <=
            Ic1927bb3335f6a28c0816eba12d3975e ^
            I5b8a1e1a6b904b0f6822c224ee0486e3 ^
            I8be4711146486fea913843e497065b50 ^
            If4c36727ab1c29bf78f72e8acfc00d7c ^
            exp_syn[62];
          sgnprod_00063 <=
            I9b096ce09467c10f448496fda13987d2 ^
            I57b7b48f13436b19a8d6a47e014eb41f ^
            I5446c1c323774715371c73bd1be66697 ^
            I6426943b4ab66f17c2b7b399ccc7a6a9 ^
            exp_syn[63];
          sgnprod_00064 <=
            I595665d8128bb87ab62741d7ac520a4b ^
            Ic920452d5997a8477724fa78c86c0fba ^
            I3a8e9e7d2cd6751e8500a5567cef5acc ^
            Ib0dadebad37d9ea9d01350054872863c ^
            Iddcffa815489773b3688fd68dba18bd8 ^
            exp_syn[64];
          sgnprod_00065 <=
            Ife0952b85f14a960007b67646b0cd969 ^
            I4d54dd2ee2f32909098d3cc2b6689220 ^
            I797c9cb725f88c07be28f017871d17f8 ^
            Ie165d0729542c81ca89f45d15e0afd3d ^
            Id00642563679fa9a6696f8e7bbdf6576 ^
            exp_syn[65];
          sgnprod_00066 <=
            I258c45897919cec5c6acaddee7f3a41b ^
            I1e11f0088959aa40b4ad1a047b59caf4 ^
            Idce46f6d03376bea1ba361e8c59f8bd1 ^
            If17c0096ce34b88007247bf4c429d5c4 ^
            Ifda1c55899cd3506853cc82b450b3936 ^
            exp_syn[66];
          sgnprod_00067 <=
            Ic69094123b75ae36e3e54f179a9f2cb5 ^
            Id182a776b03f48fb139c28194ae7ab6b ^
            I65171c9ee8449407484e5c82d13c6751 ^
            I92eb6f60c14ee9eecb01718b01ea980f ^
            Ib5d1a7cdbcba0b654c12063d4f1768e1 ^
            exp_syn[67];
          sgnprod_00068 <=
            I07abbbd75d91018ac53f53e64cffafb9 ^
            I4cdc955fa9afc75c2c977de4ec540e1e ^
            Ie79ce8adeef2c3c24a3386f054d0cf5b ^
            Ifc2963762403a00c4f3662b2863c991e ^
            I5e8ed024e2f2548bb375a2ecf1918a5f ^
            exp_syn[68];
          sgnprod_00069 <=
            I256050251d23250854ff337bef28e460 ^
            I20ffba20af04b99954bf719589e90d1a ^
            I7353ebf3a1cde89d2bb3fa667f7f5485 ^
            I97e82e5f6775d1e31537b891597223bd ^
            Id25deba967318f049de8163e67262f4b ^
            exp_syn[69];
          sgnprod_00070 <=
            If876ca6a14ffb4323503ed46666bc25f ^
            I5109afc4dc91780e05704ea5e1399e3e ^
            I621b20d29d3a9a9f41065bc3c3bbd2d8 ^
            I76fd9005abd511c3c5bf6c77de8bf2f3 ^
            I925f6b549a25cdc8f85152eb21ea3b58 ^
            exp_syn[70];
          sgnprod_00071 <=
            Ib42d37576e3aff3d205f1f8822cc58b5 ^
            I3ce10718a2211184999663c3c2493cc1 ^
            I06b48093d4c9b0327c3efc6fa4ca7daf ^
            Ie8e29053f122a9247b0dec291c6ef4f3 ^
            I9b49e1acb81ef5b088b808d2e4ce9954 ^
            exp_syn[71];
          sgnprod_00072 <=
            I364ed3f83c49626bc3b939e53524d9c7 ^
            I8188dd7cb03854c6f709de06ff785d91 ^
            Ie7cfdd25541414ff3f8d6e5d7677fbe5 ^
            I6386a4dd26e7c36165dc265b3a2c93cf ^
            exp_syn[72];
          sgnprod_00073 <=
            Ia659126b51468cfef48c97a135a71500 ^
            I866b30a63b3b5fb708934a1cbb0e1d9a ^
            I2b7822d5d77aaed61eee87570564df76 ^
            Ia20709f08cfff3a51d4af1e81d640400 ^
            exp_syn[73];
          sgnprod_00074 <=
            If1c0a3726041f70e508d68cbf6e40e04 ^
            I019e399a1cef87745e025a7d74e94db0 ^
            I0dccb8eaad52ce4d780696a8485420f1 ^
            I1ff042bdb52aac5d69791e96e2f9706c ^
            exp_syn[74];
          sgnprod_00075 <=
            Ice1ce5b4c30841dd92268559ebadafcf ^
            I3d149293f106ae8680c7f4702daa0bd6 ^
            Id17ada8dae3f9810d1892d34f2288859 ^
            Iaa2cbf59f6f61198b4fcf5a741cd5bc8 ^
            exp_syn[75];
          sgnprod_00076 <=
            I3eeeb1949945032d6c1759875426b733 ^
            If2dfcbf493b761fb5d7c622e739b23f3 ^
            I3f5053e519a928640ae49cf4e5b39d1e ^
            I01c94743a11042e75638ba6618356203 ^
            exp_syn[76];
          sgnprod_00077 <=
            Ic2b000c3b2ca3beff2d427caab04701a ^
            I1c2ee281cd47a8414851c5e1c758ea65 ^
            Ia3ef2f70c5abaa852586a33c505aee0d ^
            I0a0340a0e52145f3597accfe4a4e8624 ^
            exp_syn[77];
          sgnprod_00078 <=
            I3c3c22bf63e55a81ae91b1dd1ef615a0 ^
            Ib02268d5048c7c8e83118070e927453f ^
            I30be0b18e4415ca50f2d8149efaaafe6 ^
            I3bb4d24caaa0882a75125e466070f0b1 ^
            exp_syn[78];
          sgnprod_00079 <=
            Iaf36ce8598a29573979c683a5e2cf9fd ^
            I82f0e5a32d1bcd761a74f1f9ce8c88ba ^
            I659322a9fd0d5eac514437b02e0491b3 ^
            I44ead0ab5ccc53226fccc03024643771 ^
            exp_syn[79];
          sgnprod_00080 <=
            Idc2a9c6dd8d2aa912548c918c8a488f4 ^
            I08f22261d5713c0636d77c7938f592d6 ^
            I04c734eb876aa722e84d6b9edd297978 ^
            Iaded125f7fd5c833e7206dd7071069be ^
            exp_syn[80];
          sgnprod_00081 <=
            I98febac90cccb5fc1f3d966b6e38c4d3 ^
            I0038305f94aaefe2cd1a243580d95932 ^
            I0d41bef808860bde56d48792764612d5 ^
            I373be7c3f9511a2906584e33e5048abf ^
            exp_syn[81];
          sgnprod_00082 <=
            I2c8f4a147b363d9c5ef0e080d9a9ed40 ^
            I9171019227f35760d02d0c8ce786f4d3 ^
            I669d34b955d2991ebbb31c149ad1b6f8 ^
            Ie0b5f51835ebdb508a596eeebf0e4847 ^
            exp_syn[82];
          sgnprod_00083 <=
            Ie644d131c4f2c603e8e64c5581fdf822 ^
            Ib70e99c3acc76286a6811bcacc9284de ^
            I263aad78110a1136eb7012c6983b2a8d ^
            Iddb75e0197b9a76b36a59ac2a7ccdf3a ^
            exp_syn[83];
          sgnprod_00084 <=
            I8e873fb2321eea82bb590a92411e2e2c ^
            I6cde57127c5bd2732e71ecb7738fad6d ^
            Iae6ed7748692f2edf1aa9d73380075f0 ^
            I08c03198b9599b2f4590e3022e398f7c ^
            exp_syn[84];
          sgnprod_00085 <=
            Ia62832d325f86160285c4d1a790a32cb ^
            I2f23d4cdb6f5f827513aa60266936e4f ^
            I4b99891bed4f5c149cd4a5b4f1dde0f0 ^
            Ia4f3cff223e24815ee1d86bf41756f06 ^
            exp_syn[85];
          sgnprod_00086 <=
            Ice82cfe55a5f226746e59e5c8beb46be ^
            I09031235f61238b0e32ff52641aab70e ^
            I9d7614d286377329eb3999213889b707 ^
            I56592e1452c4b559af19465b30230ec0 ^
            exp_syn[86];
          sgnprod_00087 <=
            I384d5377ee6b8f7eb2db23a2e444ddbc ^
            I477a920e2326828bf026b0a6b6a18e2b ^
            I5196382b75d16892d550f17893de15ec ^
            I213ce488e5345fa405a9c5df297d6f74 ^
            exp_syn[87];
          sgnprod_00088 <=
            I5ad7eb9d3ce7c712515254f892d1670d ^
            I914dedc1d5e5e21c9b8d07ec0ecc01f9 ^
            Iefac1e428116a797c2c0803410ac5601 ^
            exp_syn[88];
          sgnprod_00089 <=
            Ib534288c2cf976b6ec85db743bc2a823 ^
            I90023493600924a76d2192080cf6194e ^
            I8b419d5827e5b1af9649d602401c189a ^
            exp_syn[89];
          sgnprod_00090 <=
            I485f9d1104a965d5d035feef912a2ca8 ^
            I474f6bd977f4197742d0bddb3bece684 ^
            Ie989550c9101de382056dd60d5da0e01 ^
            exp_syn[90];
          sgnprod_00091 <=
            I9b76f0121a3f7e887e7121db50024ab4 ^
            Ic3fb524ab434e80b3289c9241b65d224 ^
            I259010e323e1e8dcd9dd719091131f6c ^
            exp_syn[91];
          sgnprod_00092 <=
            I30d615203b697787ead37394953925cc ^
            Ic9146d8b3dd0c612073b70b8a8791e8c ^
            I3e0b41bee4c76eb5f3340ad23bfa01ad ^
            I389ac86954fd70464c9550e3fed4ed33 ^
            exp_syn[92];
          sgnprod_00093 <=
            If4cb744ee52b6ae793431cd038069b57 ^
            Ic3cb34aae74c5f1a870b3635f8a40764 ^
            I877e8d94236c3d8b0a31858a98fba5d6 ^
            I77371f0e55b4684d1af196ed52d3d997 ^
            exp_syn[93];
          sgnprod_00094 <=
            I83c7d177eec2dad0a924557cdc91ba77 ^
            Ib1073489d63ea33d7f3892f4ff875358 ^
            Ieefbb5d6f4ac1e586832c5c0f513c5a2 ^
            I5a21996f5724a2a49fcf8e928c01b062 ^
            exp_syn[94];
          sgnprod_00095 <=
            Iea1297491d1dfe98f395d8c73808a893 ^
            Ie9236599cea94cfb603c6b977fdbb44a ^
            If8fe5af7e5c3c97b5a713f6bcf919f1f ^
            Id46108963921efa50aff64d4dd7d1701 ^
            exp_syn[95];
          sgnprod_00096 <=
            Ife25829fb3c5023b7d69bbaadf9cf77e ^
            I3375fff5ee0d4b4b12c5a70fbdee59fe ^
            I68c35d63dc95baff41b4dc27a86d2342 ^
            I8da50e5093acefb6f809aed64564a53e ^
            exp_syn[96];
          sgnprod_00097 <=
            If988b82b86db1f4ff6d3695f7b0197e4 ^
            Ia9f5ce4603af279bbd9b486b67016482 ^
            I0c5539373b3868d0664a92157b4b4226 ^
            I03b0694777d0160a83cbc82ac1397736 ^
            exp_syn[97];
          sgnprod_00098 <=
            I10fca5f2cbf5e2bc3433c0dda579a051 ^
            Iaa1e981134f5a5c02983c49562683bc5 ^
            I6eea5fde8e2517554ad6ba25018572dc ^
            I85c2bffb93569d9fe1b1bcb10b98bcac ^
            exp_syn[98];
          sgnprod_00099 <=
            I9eaf4e9ebe07717503ff69b51f0e1905 ^
            I23c8b64e433af0bd00cef44e38df99f8 ^
            I7bfb4c5d9e22d1bd8811844d9c74dff8 ^
            Id00274c88b93867a80606343add1cdab ^
            exp_syn[99];
          sgnprod_00100 <=
            I7741e239c16828889d488cc87647c154 ^
            Ic828cdd5dfde844df4c150921af2a443 ^
            I61e829cbf7d6c0ef8ddc11677981e2cf ^
            exp_syn[100];
          sgnprod_00101 <=
            I7050adb9d06f767549b7f35c4679e391 ^
            Idc5fb0f3a04ab32948e249e088a11b11 ^
            I9e8ae2aed048068b01b3bd46f30baae8 ^
            exp_syn[101];
          sgnprod_00102 <=
            If43dd31198c8a0da6fabd194cf13bb70 ^
            Ic0732810fd355d59a3168be896a0f9ac ^
            I7dab71adbe62687846fc027d2789451d ^
            exp_syn[102];
          sgnprod_00103 <=
            Ib16548d471f0a4f4625852ea04335dcc ^
            Iff2f1716cbd73b406d8f07c22dc79fc8 ^
            If1295608bd218ed60922a0b95bf1d098 ^
            exp_syn[103];
          sgnprod_00104 <=
            Ib051eb1091a85f85a1e50007f1b27cab ^
            Ibdad0ab78e4404c852e60a2b04c3a5f6 ^
            I5fdd8e1550feaecd81b82069fe73ed7e ^
            Ib4ae1cedd09d72c235765a6cd7e91366 ^
            Idf04e08c120ed116af14a62659675b44 ^
            exp_syn[104];
          sgnprod_00105 <=
            If6a5dc79c0f6ce348956286737a369d8 ^
            I6d4fc81ced37c159303c243af04d345e ^
            Iba1c0ebd9cefeb0dd7f690bdbbbfec58 ^
            I3472ee8c06644490252e606b62bf9bd5 ^
            Ieb7614ad1b1bfed3e2b0089a72fe214a ^
            exp_syn[105];
          sgnprod_00106 <=
            Ia8e304ca12c82e41cb8e4de7be199394 ^
            Ia2c5fe53cb5b318fa63d09881609655f ^
            Ic124975d36a292816146a2fe61ab3ab9 ^
            I3eab1582cc42db0ac7739386cce2a712 ^
            I589062eca318b25dfe5735da455b6fe1 ^
            exp_syn[106];
          sgnprod_00107 <=
            I05721e06a1acdcc0571907c7d853f18c ^
            I1e93f0470d2818249f1c28ef2a399a0e ^
            I453dd7d7c0a2f003f0b67e909630d641 ^
            I6387919f2426c283e2d70e471cda54a6 ^
            If3db87afb3ea184c9e4020c5e45cb161 ^
            exp_syn[107];
          sgnprod_00108 <=
            I7979161aa1e2262ebea862004c387697 ^
            Iaddc1f2e822fd2fe9d9046d759a82cb4 ^
            Ia14bc1fcd5bbdcb60b8e68298f7d716a ^
            exp_syn[108];
          sgnprod_00109 <=
            I04aacd95d9e44657f616e01c9053f0fb ^
            Ia8974083bfd064f2c27dcd421490fcfd ^
            I268b60cb371b3d46dc3f8b0009f541b1 ^
            exp_syn[109];
          sgnprod_00110 <=
            Ibeb8c72b90b50c6897224ca1a792fa56 ^
            Ie232799bd6c4ec99e24c78f3ad798265 ^
            If2cd93b57cd1c2b91ee7a73a97dd19f2 ^
            exp_syn[110];
          sgnprod_00111 <=
            I0987c561670b7b2b6683303c1be39561 ^
            I3b30b4ab00a49e10a75587aa324d6132 ^
            Id81305359a07db527e49fda05cd2784f ^
            exp_syn[111];
          sgnprod_00112 <=
            I8b2a79aa4ac88e6b4ca8188a7852022e ^
            I6b5645cdde4b35a16fe3e91d90caaa4e ^
            Ibc48fabc172f27ebce18d0a9b5120dc5 ^
            Id8292eca087c1a17dc8b5a572a76f21f ^
            exp_syn[112];
          sgnprod_00113 <=
            I6ef260ef75e47b011a46ba2080ac3684 ^
            I34e6e9d2153e4a70ee36ab85e72d5318 ^
            Idf1ecab26889c4adcb835fda6b1cb368 ^
            Iddb19725b093506e5e521d8d68dcb8e1 ^
            exp_syn[113];
          sgnprod_00114 <=
            If8572800d5d80cc92dd917b60447b63b ^
            I3566f2779e860008b1a5d305366a07c9 ^
            Ia9f1e580e8f441394d719d52a7bad688 ^
            I0b573d3a86a3111451da661e46384876 ^
            exp_syn[114];
          sgnprod_00115 <=
            Icb0841ecf142687c3aa23e68f01c927c ^
            Ibfcfd3151af0d82bfce293ada44059b3 ^
            I220e32641265b46527ca61111f7ebf1b ^
            I0ff479e61d1a0cede88ebffb073c60be ^
            exp_syn[115];
          sgnprod_00116 <=
            I8e87530a131b5a73cad6df68b9e4967f ^
            Iee17ece482d04964d3c21a092ec955a4 ^
            Icd6f8f5df6b4ca4c81855e974db76526 ^
            exp_syn[116];
          sgnprod_00117 <=
            I2bdf4736022e5da7294a0e851006a124 ^
            I1c7e41b9cb1bdb6f649c88c0ed3f4100 ^
            I7ce064a756dad56d37684d5d7d168047 ^
            exp_syn[117];
          sgnprod_00118 <=
            Ic62fc602da3d16fe13d03a49a21269d0 ^
            I5364deb983adc2ae505ed2b8c57f876d ^
            Ied2ea62cfb21602645babc36e27b8218 ^
            exp_syn[118];
          sgnprod_00119 <=
            I2ff317d57f59747c4524ef4278d51092 ^
            I6e92a48aaab94074a555efa9bd1e7243 ^
            I79b85da6e5ce0b02ebd1619115c98e24 ^
            exp_syn[119];
          sgnprod_00120 <=
            Ie68b31360c12a83c6095254b6f14603c ^
            I00d3f14b20e1ea7d726533386e0eba27 ^
            I579c7926e7b78f4ffc606adc10522f53 ^
            I837183265ee22d080e81fea468ab0887 ^
            I8e1ddd7e4185c28caa71d30bc28138f3 ^
            exp_syn[120];
          sgnprod_00121 <=
            I9539fcc40d26b13015a864718b116d5b ^
            I02849282dd1bd663fd39baccf41762f9 ^
            I5d6e576b0fa7e3219aaf9ccc345085b8 ^
            Ic0191941cb968bbd7644c21767423d2e ^
            Iab0bff1633e2f3ea0bfbc291f3ab5d29 ^
            exp_syn[121];
          sgnprod_00122 <=
            I8850ab26807dcd55fefadf6310729ca7 ^
            Ice59d2af73d0b0f2ae91a2ef0c2b7f04 ^
            Ic4efba3932e598784f5b9ad6ad04772d ^
            I9ad2f6fd2d7f68011fc926ec9abd5c34 ^
            I5f0751fceaa008feba5c6867ced453dc ^
            exp_syn[122];
          sgnprod_00123 <=
            Ifdabf743a8cb46b7053000ff48ea0c60 ^
            Ie562ebb336e476a81f20a652d4cb20f1 ^
            Iefdb8bd28839af9413a3906cbfe715e6 ^
            Ib9d58222da98f29fa302b4896594fe26 ^
            I9f6751c15237c20b0cf2175575195ea7 ^
            exp_syn[123];
          sgnprod_00124 <=
            I081e2595b18f306a74d070203447ecf6 ^
            I3b84dad6d0dd8730312b3e20c6d5a2a8 ^
            I6ea50be10bc990a1206cdc9e28e0c4c2 ^
            exp_syn[124];
          sgnprod_00125 <=
            Ifc1da524e7670772834d521a6fc4c96f ^
            Ie2d946edaddd3c87f328e861f3e72c0a ^
            I43c2fab87f70ea883321ab82de85f133 ^
            exp_syn[125];
          sgnprod_00126 <=
            I24645082ef16129eed1c574f5fc601ca ^
            Idb1efe99b5d7fd567a7f82cfd52f7eb8 ^
            I1af02ed6cf00d4cb0704b5e44c83bfa3 ^
            exp_syn[126];
          sgnprod_00127 <=
            Ie8c0fac00a9de74870e59cbf9e87a39b ^
            Ie4827dc0983c1a63053c08de6e36d375 ^
            Ib71611afdd0381cc1884f5ddbbae1acc ^
            exp_syn[127];
          sgnprod_00128 <=
            Idf8d15c7bd7705b9aafbda09c3a5b46c ^
            I7f720a18542528f0c9bfb14f699ff4da ^
            I70a4926e9e6a05fa9ee51a26988862fe ^
            I38fc49afce0298846ae8ed63ae715e81 ^
            exp_syn[128];
          sgnprod_00129 <=
            Ic6fd9592d2ffcb8f4ca83c6f0bd19975 ^
            Ie4cda4648f6ceb76b8fb74f290ab6439 ^
            I5707d30ca29842b6a96cfaeb44ac6668 ^
            Iddc3e44d83e8253e5129b6cbf5082df7 ^
            exp_syn[129];
          sgnprod_00130 <=
            I94009bb7239be96243902ab0f0abea7e ^
            Ic308610ea8bb62ecb6094192e02dbdba ^
            I85654bd3a07b4329aba17d8b27777f4e ^
            I975a87bdda30c5b6be8d2f0e4b107450 ^
            exp_syn[130];
          sgnprod_00131 <=
            I8bd2a9d90074500698b302cb8db7f03a ^
            Ib5ee5a6ffc45ed1fece0822dc4619b57 ^
            I235c3a9fd3e8ea1cee762c10bc8e2c53 ^
            I582bd96afa764ded148202f738b7a1df ^
            exp_syn[131];
          sgnprod_00132 <=
            I5490039998187a1a2efc3549e3dee7d6 ^
            I0615acb0f7cf79b5f6ae8e91cb525dc9 ^
            I7ec15b73b2811b44e1e50c74a9f921e9 ^
            I6fb88d97bc9ed37a06b729020a1df140 ^
            exp_syn[132];
          sgnprod_00133 <=
            Ic5cb81c821716a8aabf8cc2283ff73ba ^
            Iffa06a336949f56f4e5a88a06d8b7e60 ^
            Ic68f500938d80460ffdb33a0adc48298 ^
            I1500943c4a550e78fc169437b0a663b7 ^
            exp_syn[133];
          sgnprod_00134 <=
            I22f5bb821a2571d1764978fd76c8f1d0 ^
            Id962beade26396738ba0e97f67d5e261 ^
            I7c965c047d862c973d09a81abe03a845 ^
            I0b83f4ef8ba9badb27e81b32765ec5b6 ^
            exp_syn[134];
          sgnprod_00135 <=
            I42ae0c42360c977b35429ce290516a6f ^
            Ia03836a4e93d2f36513227d1dfaea0fa ^
            I6d423a7d17e05a3c597ec6ef6c5a7cba ^
            I2c420acf428e44cdd9ca9998e276f258 ^
            exp_syn[135];
          sgnprod_00136 <=
            I14bf11ad80890227e47fda26ae1b9c24 ^
            Idd474d80b50992537d6f527faf279800 ^
            I2eed3d32a27d51036e17c4a21382b4c1 ^
            Ic7b6dae3017b55dd3cd27423d5f1b0ec ^
            exp_syn[136];
          sgnprod_00137 <=
            Iae7b72abf4d3c536330a229e3836b441 ^
            Idc5e98f6958786ccf95d39b922b42ea9 ^
            I2a4bbedf880a9a7b4e1bf946f9f96c0e ^
            I4a91a7c9b2a0f3552b8f2ef4e2398be2 ^
            exp_syn[137];
          sgnprod_00138 <=
            I3b8cdfb1440732ce98cd1676e05a2af1 ^
            I3fbd40faa4c3b78b547b8348c466fd1f ^
            Id6b508145cd21ba088ab8fda34577c35 ^
            I99ff29c7ba68b5d0819f1e1bead51287 ^
            exp_syn[138];
          sgnprod_00139 <=
            I2aea17846a53e2eb2968581ee2c48226 ^
            Ibf2a253afde05c905d0b2404c5a808a0 ^
            I24f82a3f2c0e8df486fe495dd95cf8bc ^
            If06b00be0356a2be5074d958ddcdb2f9 ^
            exp_syn[139];
          sgnprod_00140 <=
            Iae5d6faac1f5685cb1d400ee2b1d85e0 ^
            Ia98a6f01e4eb5bc74d50d350e79be426 ^
            Iabb01dc9980b4879a7356712b51df0d6 ^
            I604283449f13c7b225ea03f99f2e296a ^
            exp_syn[140];
          sgnprod_00141 <=
            I68b152a599887c0039dd9d45c528c219 ^
            I24135210c23b2422a42c90ee25594191 ^
            If4308ed204e33952c9931f8fe257aca4 ^
            I2b600e5f5c146ee97c4044c08e1f5ad5 ^
            exp_syn[141];
          sgnprod_00142 <=
            I852d5295a32984af00c95f6d9389555e ^
            I33ee415d85e2bcd8f975d34b880f6ea7 ^
            Ifb89e7ad8ef661959d82b7c22f187243 ^
            I9fe16403fc21bb1159a5e0305fd1ef69 ^
            exp_syn[142];
          sgnprod_00143 <=
            I207a0f6184a0b3be71766a8b47ea5535 ^
            I86ba73ee348f80e2f9891d2ebc8a02ed ^
            Ib6ae81df8db1dae269437861ee11ec0d ^
            Iabdb9374e5caee281c25b003624b2c4e ^
            exp_syn[143];
          sgnprod_00144 <=
            Ie5d9cc18b2dd300132470f206452ff17 ^
            I1b695aa715615662eff7065c742b0859 ^
            Id0ab747d92288f23cef793567b2363d1 ^
            Ibd12036702fe60b57354b3aac921559d ^
            exp_syn[144];
          sgnprod_00145 <=
            I671de3d408b5b783541663c7f1e3a6fa ^
            Ibe01835305315fab50269c72ef849b61 ^
            I138fb0c48f2d27e3315e237d9e61d653 ^
            Ib1639811de6eb1c38257800c201fb704 ^
            exp_syn[145];
          sgnprod_00146 <=
            I169d8f2bb5fde5b202b4239b7a7f1ed5 ^
            I2b97a79c90f6578c8b2f321f8d598cc8 ^
            Ieed4c810a5bb69de112522dcf00b16ed ^
            If926d98f659e8fe4bbf36ad2c5c852c5 ^
            exp_syn[146];
          sgnprod_00147 <=
            I8ca17b6cf35e1b1f8f601604575d3f27 ^
            I9a6923c6368526a53ef70e16471386ef ^
            Iaf82668eb49248709540f2f529f1b3e4 ^
            I211f8d7f97ebb8eb3e50313513abfb1b ^
            exp_syn[147];
          sgnprod_00148 <=
            I0fd2f706e374a4eb57ee26ab50201e15 ^
            I83ecf12f3b38fc14c3b75e47b71ecc09 ^
            I304ac9f96945546cdf1b6f1fa7136731 ^
            exp_syn[148];
          sgnprod_00149 <=
            If5ae6fbf843fdeee17945bc5ce81aec8 ^
            Ie039ab562e9cf90289047b5425186123 ^
            I7a9800418bd5c195fc47a72370680b56 ^
            exp_syn[149];
          sgnprod_00150 <=
            I9b8023f4dced915cd52c91bc9d4ed78f ^
            I49d35ec6369de10afb15be8e0cf135c3 ^
            I5f6a61c9f0c67510e148e596f553a4d6 ^
            exp_syn[150];
          sgnprod_00151 <=
            I48e3309c61918c3991852b45d9c72ea5 ^
            Ifa6e3541f5e12bf9677ffc51d0392749 ^
            I8e313ceb21359bcc44114ab217b1c394 ^
            exp_syn[151];
          sgnprod_00152 <=
            I3c0a621dbef864fd1f566bc2e47f32c6 ^
            Ie61f299252b8fecfd3e8634b64df5a90 ^
            I33ddee677715877c11a1df45cbfb01ac ^
            I4c9518755c33d725221ad79ee6badba9 ^
            exp_syn[152];
          sgnprod_00153 <=
            I5cac08dabbb6de3b01c821d4db93a8e3 ^
            I1e96d5af3d0e3fdce39530dfd0131a7d ^
            I373841aa2bcbad8232d54ac9035a3ef9 ^
            I3c3cffec9f47c9979cb9503f222f370c ^
            exp_syn[153];
          sgnprod_00154 <=
            Ib62b02ddf0f57bee49838d19783ef6c3 ^
            I182b43872d50de6f7afb700f178b160e ^
            Iddcfab4a7022e0f12fd20cb34e9b9d02 ^
            I68d6769541fdc3df321e192f645c667f ^
            exp_syn[154];
          sgnprod_00155 <=
            Id051f1d5454802e0eb37e22248efe8ca ^
            Ib08897f9216599042f7b97b137e07fe1 ^
            Id1dce2b9eafc35fa71df33ada4aac539 ^
            Ided55428cbb77f454c2607ac783d7548 ^
            exp_syn[155];
          sgnprod_00156 <=
            I275cd09649a750edb8ae8313e4e1e279 ^
            If533578cacb685a95afbb8e1c05d3c07 ^
            I8879df010bbdf6e5fc9370e2fb3289b4 ^
            Ifd3d4f3e2a388b3c70e7704d6351e0ba ^
            exp_syn[156];
          sgnprod_00157 <=
            I7c791c854d0bc28e8dd787545f8fbda0 ^
            I90b3708abdf742370f06cc513ee307e1 ^
            I9a403c511fe2d44472ab319a9477199c ^
            I17d32f292758416fe02527dfd938fa0d ^
            exp_syn[157];
          sgnprod_00158 <=
            I446857735e680cae93a24dccb59b1924 ^
            Ie536879e6fa9be65376d7f00e0fc40d0 ^
            I3ade5535a79ce83857481ac771cd8618 ^
            I9ce3942aba354c1fd7d6b9a39c994d7b ^
            exp_syn[158];
          sgnprod_00159 <=
            I40a223380fb4414a3f26a08cb90025ec ^
            Id0b1c46fa4caa63a4c63a44ba3c5ef8a ^
            I88a89b2d938552458dab9bc34728959b ^
            I2c6c6041c9c69c84f4d64af6458955f5 ^
            exp_syn[159];
          sgnprod_00160 <=
            I0c616f736879c28a5222de3d6f49a587 ^
            I44f170d02bae7fe044456e125a98451d ^
            Iefbdf686d9452a62cb99cf023a4d9fe7 ^
            I830a4fffe1244e071eb82c28ddc4a308 ^
            exp_syn[160];
          sgnprod_00161 <=
            I620b8ecdcaccc1ec80ebcf9fa6af0017 ^
            I94460b6ce7b776bcc5eca149eab80c26 ^
            Ic3ba4531855366e9a060cec1c7694844 ^
            Ifad8e46fc3844bbfaf434a14f6b5869d ^
            exp_syn[161];
          sgnprod_00162 <=
            Iec91b3ca3b54010755d57f8b8ea4a544 ^
            Idc6b6357741c9887a9db1037ccc2d922 ^
            I21e72a7e5870151c3247d15121e5fb4f ^
            I10a6c6a8fdb0003de1f360c148777d0f ^
            exp_syn[162];
          sgnprod_00163 <=
            Id806a2df1c4519bbbe811791cb4072f9 ^
            I472352e7027b9df2fa957d9fd68443ff ^
            I74cbc0ec3bb682e0f927890eef8d7a58 ^
            I4cde586fc28f8d03fc9934d56f7ff7b8 ^
            exp_syn[163];
          sgnprod_00164 <=
            Ibd59d0e5a062f149bd0e91ba76985a13 ^
            I51e14ece9ab6607f83e6ba27f3f046a9 ^
            I433dd5092cf1851cd196feade3cfa6d8 ^
            Ib83a067fb08e118dcf794902beef9405 ^
            exp_syn[164];
          sgnprod_00165 <=
            Ic4c6f707f461cebbc4c93f2ba664ae7b ^
            Icc67656ad2dd3fffae4e5abe02f8fff9 ^
            Ib6124faff821158c6a2c9a9c454ab68c ^
            I358cf9609272a4562423a85f9b2f56bf ^
            exp_syn[165];
          sgnprod_00166 <=
            Ic04828ba2db8239b093043c27476d345 ^
            I38352b363fa37f6f822fbc1a39100968 ^
            I759409e242eaeb144a53e630a8cfd514 ^
            Ic1e9d9113150ad57954c0e369259dc62 ^
            exp_syn[166];
          sgnprod_00167 <=
            Ibe6b8c57d7ff47b6fdad5fadf1f6b841 ^
            Ic9b72b2a91d951cf08cf54ed215ecaa8 ^
            Ied19cb51636bfb029ba8a2c390f97105 ^
            If7fe3f5ccbb5b279e41fd183c8ff3974 ^
            exp_syn[167];



          I5033323484d90d6bfbe03749019fc6dd <=
            flogtanh_00001_00000 +
            flogtanh_00005_00000 +
            flogtanh_00008_00000 +
            flogtanh_00014_00000 +
            flogtanh_00025_00000 +
            flogtanh_00037_00000 +
            flogtanh_00040_00000 +
            flogtanh_00044_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          If5dad13ac41b3034bdb034bc86c9b348 <=
            flogtanh_00002_00000 +
            flogtanh_00006_00000 +
            flogtanh_00009_00000 +
            flogtanh_00015_00000 +
            flogtanh_00026_00000 +
            flogtanh_00038_00000 +
            flogtanh_00041_00000 +
            flogtanh_00045_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Iac428f9f798618e1ef495c626c41892b <=
            flogtanh_00003_00000 +
            flogtanh_00007_00000 +
            flogtanh_00010_00000 +
            flogtanh_00012_00000 +
            flogtanh_00027_00000 +
            flogtanh_00039_00000 +
            flogtanh_00042_00000 +
            flogtanh_00046_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I5a6427c8f18b36d2ea18fe60a0831ef1 <=
            flogtanh_00000_00000 +
            flogtanh_00004_00000 +
            flogtanh_00011_00000 +
            flogtanh_00013_00000 +
            flogtanh_00024_00000 +
            flogtanh_00036_00000 +
            flogtanh_00043_00000 +
            flogtanh_00047_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Icc29441eac6ca7a138d45743d37505e3 <=
            flogtanh_00003_00001 +
            flogtanh_00014_00001 +
            flogtanh_00017_00000 +
            flogtanh_00021_00000 +
            flogtanh_00026_00001 +
            flogtanh_00028_00000 +
            flogtanh_00032_00000 +
            flogtanh_00036_00001 +
            flogtanh_00044_00001 +
            flogtanh_00048_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I0e7754dcbc04a4850e052ae4a2fbe328 <=
            flogtanh_00000_00001 +
            flogtanh_00015_00001 +
            flogtanh_00018_00000 +
            flogtanh_00022_00000 +
            flogtanh_00027_00001 +
            flogtanh_00029_00000 +
            flogtanh_00033_00000 +
            flogtanh_00037_00001 +
            flogtanh_00045_00001 +
            flogtanh_00049_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia30c019ed8ce395556494a92e7b42a92 <=
            flogtanh_00001_00001 +
            flogtanh_00012_00001 +
            flogtanh_00019_00000 +
            flogtanh_00023_00000 +
            flogtanh_00024_00001 +
            flogtanh_00030_00000 +
            flogtanh_00034_00000 +
            flogtanh_00038_00001 +
            flogtanh_00046_00001 +
            flogtanh_00050_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I9799695ea8244992a6694eaf5c8ae64d <=
            flogtanh_00002_00001 +
            flogtanh_00013_00001 +
            flogtanh_00016_00000 +
            flogtanh_00020_00000 +
            flogtanh_00025_00001 +
            flogtanh_00031_00000 +
            flogtanh_00035_00000 +
            flogtanh_00039_00001 +
            flogtanh_00047_00001 +
            flogtanh_00051_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4524cd664b4cb41f642c675fa484c84b <=
            flogtanh_00001_00002 +
            flogtanh_00006_00001 +
            flogtanh_00012_00002 +
            flogtanh_00016_00001 +
            flogtanh_00032_00001 +
            flogtanh_00040_00001 +
            flogtanh_00048_00001 +
            flogtanh_00052_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I64e959d80af111ed2fcd54a5407d21bf <=
            flogtanh_00002_00002 +
            flogtanh_00007_00001 +
            flogtanh_00013_00002 +
            flogtanh_00017_00001 +
            flogtanh_00033_00001 +
            flogtanh_00041_00001 +
            flogtanh_00049_00001 +
            flogtanh_00053_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3e0da4bcbab4804b5397fb3aa2c94f51 <=
            flogtanh_00003_00002 +
            flogtanh_00004_00001 +
            flogtanh_00014_00002 +
            flogtanh_00018_00001 +
            flogtanh_00034_00001 +
            flogtanh_00042_00001 +
            flogtanh_00050_00001 +
            flogtanh_00054_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3740b30d31f3c61d93a14a46e3199c4d <=
            flogtanh_00000_00002 +
            flogtanh_00005_00001 +
            flogtanh_00015_00002 +
            flogtanh_00019_00001 +
            flogtanh_00035_00001 +
            flogtanh_00043_00001 +
            flogtanh_00051_00001 +
            flogtanh_00055_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ibf0a30abfec9031737eada436ac1a0d4 <=
            flogtanh_00004_00002 +
            flogtanh_00010_00001 +
            flogtanh_00018_00002 +
            flogtanh_00020_00001 +
            flogtanh_00025_00002 +
            flogtanh_00030_00001 +
            flogtanh_00034_00002 +
            flogtanh_00036_00002 +
            flogtanh_00040_00002 +
            flogtanh_00052_00001 +
            {MAX_SUM_WDTH_L{1'h0}};
          Id36e8953a02400a5ab1f4dfdb0422e6d <=
            flogtanh_00005_00002 +
            flogtanh_00011_00001 +
            flogtanh_00019_00002 +
            flogtanh_00021_00001 +
            flogtanh_00026_00002 +
            flogtanh_00031_00001 +
            flogtanh_00035_00002 +
            flogtanh_00037_00002 +
            flogtanh_00041_00002 +
            flogtanh_00053_00001 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ica71108a53bfcfd1892b4d03ef68110c <=
            flogtanh_00006_00002 +
            flogtanh_00008_00001 +
            flogtanh_00016_00002 +
            flogtanh_00022_00001 +
            flogtanh_00027_00002 +
            flogtanh_00028_00001 +
            flogtanh_00032_00002 +
            flogtanh_00038_00002 +
            flogtanh_00042_00002 +
            flogtanh_00054_00001 +
            {MAX_SUM_WDTH_L{1'h0}};
          I7c97629ec6e594f9b2160815ddd133cc <=
            flogtanh_00007_00002 +
            flogtanh_00009_00001 +
            flogtanh_00017_00002 +
            flogtanh_00023_00001 +
            flogtanh_00024_00002 +
            flogtanh_00029_00001 +
            flogtanh_00033_00002 +
            flogtanh_00039_00002 +
            flogtanh_00043_00002 +
            flogtanh_00055_00001 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4823c8239ace86dc399e906c1b5a0d74 <=
            flogtanh_00003_00003 +
            flogtanh_00006_00003 +
            flogtanh_00047_00002 +
            flogtanh_00056_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I10ad572ca72c2ea991487c39f7eabd7b <=
            flogtanh_00000_00003 +
            flogtanh_00007_00003 +
            flogtanh_00044_00002 +
            flogtanh_00057_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie9f3fd3a6d16316e55addbe0e336519f <=
            flogtanh_00001_00003 +
            flogtanh_00004_00003 +
            flogtanh_00045_00002 +
            flogtanh_00058_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I07965bca84276dd56da1af98e64b0adc <=
            flogtanh_00002_00003 +
            flogtanh_00005_00003 +
            flogtanh_00046_00002 +
            flogtanh_00059_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ic2ade31b8bcf68c4dcc1a371ff14074b <=
            flogtanh_00003_00004 +
            flogtanh_00005_00004 +
            flogtanh_00022_00002 +
            flogtanh_00031_00002 +
            flogtanh_00047_00003 +
            flogtanh_00060_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ic0edcf240048fbfde4e938c3e4c5e281 <=
            flogtanh_00000_00004 +
            flogtanh_00006_00004 +
            flogtanh_00023_00002 +
            flogtanh_00028_00002 +
            flogtanh_00044_00003 +
            flogtanh_00061_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8b42e89ff5f780d4ef8cd1cd5c99ef61 <=
            flogtanh_00001_00004 +
            flogtanh_00007_00004 +
            flogtanh_00020_00002 +
            flogtanh_00029_00002 +
            flogtanh_00045_00003 +
            flogtanh_00062_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I70b1b8521b36920707e95fc9418eb8a9 <=
            flogtanh_00002_00004 +
            flogtanh_00004_00004 +
            flogtanh_00021_00002 +
            flogtanh_00030_00002 +
            flogtanh_00046_00003 +
            flogtanh_00063_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4fb1c32a62cbbaeb585c6564a3c938f9 <=
            flogtanh_00003_00005 +
            flogtanh_00020_00003 +
            flogtanh_00029_00003 +
            flogtanh_00036_00003 +
            flogtanh_00046_00004 +
            flogtanh_00064_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Iefc37daeec14e14ef2fe0716f73109dc <=
            flogtanh_00000_00005 +
            flogtanh_00021_00003 +
            flogtanh_00030_00003 +
            flogtanh_00037_00003 +
            flogtanh_00047_00004 +
            flogtanh_00065_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ibd15f164f6d2ac9e5721a21464bc2c5c <=
            flogtanh_00001_00005 +
            flogtanh_00022_00003 +
            flogtanh_00031_00003 +
            flogtanh_00038_00003 +
            flogtanh_00044_00004 +
            flogtanh_00066_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I951dfff9507bb70214d48e03a0ebb3a7 <=
            flogtanh_00002_00005 +
            flogtanh_00023_00003 +
            flogtanh_00028_00003 +
            flogtanh_00039_00003 +
            flogtanh_00045_00004 +
            flogtanh_00067_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie78e30b2a2eda75d0df7d10fd67b5e36 <=
            flogtanh_00005_00005 +
            flogtanh_00023_00004 +
            flogtanh_00028_00004 +
            flogtanh_00047_00005 +
            flogtanh_00052_00002 +
            flogtanh_00068_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia0b83a372dd4115dc4d61eb8ff0811b9 <=
            flogtanh_00006_00005 +
            flogtanh_00020_00004 +
            flogtanh_00029_00004 +
            flogtanh_00044_00005 +
            flogtanh_00053_00002 +
            flogtanh_00069_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          If5c5bcbbea01aa22f242b913f0d01929 <=
            flogtanh_00007_00005 +
            flogtanh_00021_00004 +
            flogtanh_00030_00004 +
            flogtanh_00045_00005 +
            flogtanh_00054_00002 +
            flogtanh_00070_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Iccba58cd3519fb4cc75a61b50da1d562 <=
            flogtanh_00004_00005 +
            flogtanh_00022_00004 +
            flogtanh_00031_00004 +
            flogtanh_00046_00005 +
            flogtanh_00055_00002 +
            flogtanh_00071_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ibc0999e4d0b3cc2650f9348b8c204b14 <=
            flogtanh_00002_00006 +
            flogtanh_00006_00006 +
            flogtanh_00050_00002 +
            flogtanh_00072_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I2aeff1fb4b839a581acaf26f90f9113c <=
            flogtanh_00003_00006 +
            flogtanh_00007_00006 +
            flogtanh_00051_00002 +
            flogtanh_00073_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I7d60d53f883f8187700c4e78b4c22f1c <=
            flogtanh_00000_00006 +
            flogtanh_00004_00006 +
            flogtanh_00048_00002 +
            flogtanh_00074_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Id6fcf4b7af4a37c854a12e2ae80851fa <=
            flogtanh_00001_00006 +
            flogtanh_00005_00006 +
            flogtanh_00049_00002 +
            flogtanh_00075_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ifa5e5f7d753964f14f0f16dbe552fd85 <=
            flogtanh_00007_00007 +
            flogtanh_00033_00003 +
            flogtanh_00041_00003 +
            flogtanh_00047_00006 +
            flogtanh_00076_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I900d471b087cf5a436c2ad66a84d8280 <=
            flogtanh_00004_00007 +
            flogtanh_00034_00003 +
            flogtanh_00042_00003 +
            flogtanh_00044_00006 +
            flogtanh_00077_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6d1434907f0292ea2ee47cbc5b52bfb9 <=
            flogtanh_00005_00007 +
            flogtanh_00035_00003 +
            flogtanh_00043_00003 +
            flogtanh_00045_00006 +
            flogtanh_00078_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I938bef7ba7ae1739d8e6a6a7c117a1b1 <=
            flogtanh_00006_00007 +
            flogtanh_00032_00003 +
            flogtanh_00040_00003 +
            flogtanh_00046_00006 +
            flogtanh_00079_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6384a9416b2d1da01df1b2d7b16c5390 <=
            flogtanh_00003_00007 +
            flogtanh_00005_00008 +
            flogtanh_00024_00003 +
            flogtanh_00029_00005 +
            flogtanh_00080_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I5097a79e7cf7a30d38ba198d1407119c <=
            flogtanh_00000_00007 +
            flogtanh_00006_00008 +
            flogtanh_00025_00003 +
            flogtanh_00030_00005 +
            flogtanh_00081_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib113c26c8dcf49c972c41a938059a787 <=
            flogtanh_00001_00007 +
            flogtanh_00007_00008 +
            flogtanh_00026_00003 +
            flogtanh_00031_00005 +
            flogtanh_00082_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I970c4a25a8bce82a9d2846679029fcab <=
            flogtanh_00002_00007 +
            flogtanh_00004_00008 +
            flogtanh_00027_00003 +
            flogtanh_00028_00005 +
            flogtanh_00083_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ibe2af096ad2db26e54d8b4b3bb05175c <=
            flogtanh_00003_00008 +
            flogtanh_00028_00006 +
            flogtanh_00038_00004 +
            flogtanh_00052_00003 +
            flogtanh_00084_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie48569c467fba0c1291f71d6080ebedc <=
            flogtanh_00000_00008 +
            flogtanh_00029_00006 +
            flogtanh_00039_00004 +
            flogtanh_00053_00003 +
            flogtanh_00085_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I90e7ded06617b49cdb8b5301fe9c6a20 <=
            flogtanh_00001_00008 +
            flogtanh_00030_00006 +
            flogtanh_00036_00004 +
            flogtanh_00054_00003 +
            flogtanh_00086_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4920014f5d017f4e840dc3b88526955f <=
            flogtanh_00002_00008 +
            flogtanh_00031_00006 +
            flogtanh_00037_00004 +
            flogtanh_00055_00003 +
            flogtanh_00087_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I03b70553f1c501609400574ae7cd73f5 <=
            flogtanh_00007_00009 +
            flogtanh_00015_00003 +
            flogtanh_00046_00007 +
            flogtanh_00088_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I63c9bf68b43ed66c51b0f4c0ed92e9ab <=
            flogtanh_00004_00009 +
            flogtanh_00012_00003 +
            flogtanh_00047_00007 +
            flogtanh_00089_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          If408dfead07757878cc878131bc7d6a3 <=
            flogtanh_00005_00009 +
            flogtanh_00013_00003 +
            flogtanh_00044_00007 +
            flogtanh_00090_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia0857d63d309807789b6ff4f6028f1b3 <=
            flogtanh_00006_00009 +
            flogtanh_00014_00003 +
            flogtanh_00045_00007 +
            flogtanh_00091_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I53921b825c5e434b63bee0e1ecb7a517 <=
            flogtanh_00003_00009 +
            flogtanh_00006_00010 +
            flogtanh_00034_00004 +
            flogtanh_00054_00004 +
            flogtanh_00092_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I5e68f84e123c37f19a03c13892c77e19 <=
            flogtanh_00000_00009 +
            flogtanh_00007_00010 +
            flogtanh_00035_00004 +
            flogtanh_00055_00004 +
            flogtanh_00093_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Id5270b57c6fb4b18db3bbd0a523e467e <=
            flogtanh_00001_00009 +
            flogtanh_00004_00010 +
            flogtanh_00032_00004 +
            flogtanh_00052_00004 +
            flogtanh_00094_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3c18a84617eb21472d53e598700d7f4c <=
            flogtanh_00002_00009 +
            flogtanh_00005_00010 +
            flogtanh_00033_00004 +
            flogtanh_00053_00004 +
            flogtanh_00095_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Id36663e7a01fff3170833ecfecac1321 <=
            flogtanh_00007_00011 +
            flogtanh_00025_00004 +
            flogtanh_00047_00008 +
            flogtanh_00052_00005 +
            flogtanh_00096_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8d3be15109c7007a79fecaac0d891626 <=
            flogtanh_00004_00011 +
            flogtanh_00026_00004 +
            flogtanh_00044_00008 +
            flogtanh_00053_00005 +
            flogtanh_00097_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I92169cc57291f20d336a479e392ec271 <=
            flogtanh_00005_00011 +
            flogtanh_00027_00004 +
            flogtanh_00045_00008 +
            flogtanh_00054_00005 +
            flogtanh_00098_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6178b220b469b40dac39168057023a1c <=
            flogtanh_00006_00011 +
            flogtanh_00024_00004 +
            flogtanh_00046_00008 +
            flogtanh_00055_00005 +
            flogtanh_00099_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I55342938216a0ea0889f96c2f6c05ce5 <=
            flogtanh_00003_00010 +
            flogtanh_00043_00004 +
            flogtanh_00045_00009 +
            flogtanh_00100_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Idf28431c76a84a48dd895979d2b11a63 <=
            flogtanh_00000_00010 +
            flogtanh_00040_00004 +
            flogtanh_00046_00009 +
            flogtanh_00101_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I1ef61124c8d62e8f6a82a729fb091694 <=
            flogtanh_00001_00010 +
            flogtanh_00041_00004 +
            flogtanh_00047_00009 +
            flogtanh_00102_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib8bb96f0372323e6a8072ca56fb9396d <=
            flogtanh_00002_00010 +
            flogtanh_00042_00004 +
            flogtanh_00044_00009 +
            flogtanh_00103_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I432f74dda4f6b1cebdf5ad59c659080b <=
            flogtanh_00007_00012 +
            flogtanh_00038_00005 +
            flogtanh_00044_00010 +
            flogtanh_00050_00003 +
            flogtanh_00104_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Idc689442305acd00f0f32416d8fb3773 <=
            flogtanh_00004_00012 +
            flogtanh_00039_00005 +
            flogtanh_00045_00010 +
            flogtanh_00051_00003 +
            flogtanh_00105_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ida03738adc101c03c2229756bed2469d <=
            flogtanh_00005_00012 +
            flogtanh_00036_00005 +
            flogtanh_00046_00010 +
            flogtanh_00048_00003 +
            flogtanh_00106_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4d14c75f28f3e516c259ea288996131b <=
            flogtanh_00006_00012 +
            flogtanh_00037_00005 +
            flogtanh_00047_00010 +
            flogtanh_00049_00003 +
            flogtanh_00107_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6e6cbbf430d57f347a0d70558af143d8 <=
            flogtanh_00006_00013 +
            flogtanh_00020_00005 +
            flogtanh_00046_00011 +
            flogtanh_00048_00004 +
            flogtanh_00108_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib7487df45118e44acec6b9d07bbd5969 <=
            flogtanh_00007_00013 +
            flogtanh_00021_00005 +
            flogtanh_00047_00011 +
            flogtanh_00049_00004 +
            flogtanh_00109_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I492f382fea500462b3d0866240fb91b2 <=
            flogtanh_00004_00013 +
            flogtanh_00022_00005 +
            flogtanh_00044_00011 +
            flogtanh_00050_00004 +
            flogtanh_00110_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3fb3ebddaf28efb56092d19a1b4695de <=
            flogtanh_00005_00013 +
            flogtanh_00023_00005 +
            flogtanh_00045_00011 +
            flogtanh_00051_00004 +
            flogtanh_00111_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I22a26b7f0b1c8c16b00597732ce2ab23 <=
            flogtanh_00000_00011 +
            flogtanh_00026_00005 +
            flogtanh_00030_00007 +
            flogtanh_00112_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I2ac08a2d8c917ecb37fbaf5325cb0473 <=
            flogtanh_00001_00011 +
            flogtanh_00027_00005 +
            flogtanh_00031_00007 +
            flogtanh_00113_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I50ff8f51e75fb9ce3db983c2a0f57196 <=
            flogtanh_00002_00011 +
            flogtanh_00024_00005 +
            flogtanh_00028_00007 +
            flogtanh_00114_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I444bc340ffb7ef7b72d4d2e761d58872 <=
            flogtanh_00003_00011 +
            flogtanh_00025_00005 +
            flogtanh_00029_00007 +
            flogtanh_00115_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I039c6cac5830759529595a958b7f65c9 <=
            flogtanh_00003_00012 +
            flogtanh_00004_00014 +
            flogtanh_00041_00005 +
            flogtanh_00116_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I0584de7d919236ab138e288a27d08ff1 <=
            flogtanh_00000_00012 +
            flogtanh_00005_00014 +
            flogtanh_00042_00005 +
            flogtanh_00117_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I086402c82ec67ae09a9e6360c58904b4 <=
            flogtanh_00001_00012 +
            flogtanh_00006_00014 +
            flogtanh_00043_00005 +
            flogtanh_00118_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I1cefdc831c146187c77f861b3e2d1af0 <=
            flogtanh_00002_00012 +
            flogtanh_00007_00014 +
            flogtanh_00040_00005 +
            flogtanh_00119_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ida9c16ae57d17b6faee8a54838860447 <=
            flogtanh_00006_00015 +
            flogtanh_00017_00003 +
            flogtanh_00045_00012 +
            flogtanh_00120_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia3b9fb112f39dd0ccbf7555659369efb <=
            flogtanh_00007_00015 +
            flogtanh_00018_00003 +
            flogtanh_00046_00012 +
            flogtanh_00121_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib1bfcdc0c972aafc99116ed8c0511445 <=
            flogtanh_00004_00015 +
            flogtanh_00019_00003 +
            flogtanh_00047_00012 +
            flogtanh_00122_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I7adff505c50450a04f1717cac1adebe7 <=
            flogtanh_00005_00015 +
            flogtanh_00016_00003 +
            flogtanh_00044_00012 +
            flogtanh_00123_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I699feb4382974a02b21cb387c13f7f3f <=
            flogtanh_00000_00013 +
            flogtanh_00034_00005 +
            flogtanh_00054_00006 +
            flogtanh_00124_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Idc99c3b23e49aca3c98f0685ea34441c <=
            flogtanh_00001_00013 +
            flogtanh_00035_00005 +
            flogtanh_00055_00006 +
            flogtanh_00125_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib67318fa6954ec8f3247927d34e74f8c <=
            flogtanh_00002_00013 +
            flogtanh_00032_00005 +
            flogtanh_00052_00006 +
            flogtanh_00126_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8774ce3f11362915c4331d1026e452dd <=
            flogtanh_00003_00013 +
            flogtanh_00033_00005 +
            flogtanh_00053_00006 +
            flogtanh_00127_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I2392b2d17ffed6073875fbe8e92534cf <=
            flogtanh_00006_00016 +
            flogtanh_00011_00002 +
            flogtanh_00128_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3a4f0d3e32596ef05477f494768d4266 <=
            flogtanh_00007_00016 +
            flogtanh_00008_00002 +
            flogtanh_00129_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Icd08ff59cf6be3ba97698dd55703339e <=
            flogtanh_00004_00016 +
            flogtanh_00009_00002 +
            flogtanh_00130_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I985fb7ed22a8476ea322c9e3c2b3851c <=
            flogtanh_00005_00016 +
            flogtanh_00010_00002 +
            flogtanh_00131_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib985709316b1b0a9d3fa3c1eaf6c641f <=
            flogtanh_00003_00014 +
            flogtanh_00015_00004 +
            flogtanh_00022_00006 +
            flogtanh_00132_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4be898887dff6e2cebe53f135ece131b <=
            flogtanh_00000_00014 +
            flogtanh_00012_00004 +
            flogtanh_00023_00006 +
            flogtanh_00133_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I004db04f61fb57aba81e15cc015442b3 <=
            flogtanh_00001_00014 +
            flogtanh_00013_00004 +
            flogtanh_00020_00006 +
            flogtanh_00134_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8f7e3dfb2f728d4cd1e79b82b62b0406 <=
            flogtanh_00002_00014 +
            flogtanh_00014_00004 +
            flogtanh_00021_00006 +
            flogtanh_00135_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I991054370345e61638ddaf81785505bd <=
            flogtanh_00006_00017 +
            flogtanh_00011_00003 +
            flogtanh_00036_00006 +
            flogtanh_00136_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ifa1f503965270d10e7a5c9a15576069b <=
            flogtanh_00007_00017 +
            flogtanh_00008_00003 +
            flogtanh_00037_00006 +
            flogtanh_00137_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I24f773842a4742fb58d09cae45717b2f <=
            flogtanh_00004_00017 +
            flogtanh_00009_00003 +
            flogtanh_00038_00006 +
            flogtanh_00138_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I5bac7e0d778a547a0ae764fe259b6f7a <=
            flogtanh_00005_00017 +
            flogtanh_00010_00003 +
            flogtanh_00039_00006 +
            flogtanh_00139_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I255577ebee6768871df0224fc1db2db3 <=
            flogtanh_00000_00015 +
            flogtanh_00020_00007 +
            flogtanh_00140_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia7fb4af3d3529a32f902a52cf5598474 <=
            flogtanh_00001_00015 +
            flogtanh_00021_00007 +
            flogtanh_00141_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I2c98806141f064c9e92935b23a84ede1 <=
            flogtanh_00002_00015 +
            flogtanh_00022_00007 +
            flogtanh_00142_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I5680847bc8d224fa4ed93b2fc0d841e1 <=
            flogtanh_00003_00015 +
            flogtanh_00023_00007 +
            flogtanh_00143_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I365254279ebb10dd7ba0b3482d5e34cd <=
            flogtanh_00009_00004 +
            flogtanh_00031_00008 +
            flogtanh_00048_00005 +
            flogtanh_00054_00007 +
            flogtanh_00144_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I57bf4ad773cc058ae1bb7b1911dc3174 <=
            flogtanh_00010_00004 +
            flogtanh_00028_00008 +
            flogtanh_00049_00005 +
            flogtanh_00055_00007 +
            flogtanh_00145_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I57072dfb29c4a3d2e2b40e46e62f0d95 <=
            flogtanh_00011_00004 +
            flogtanh_00029_00008 +
            flogtanh_00050_00005 +
            flogtanh_00052_00007 +
            flogtanh_00146_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Id8cafb6f76321bdaba9711133be7be99 <=
            flogtanh_00008_00004 +
            flogtanh_00030_00008 +
            flogtanh_00051_00005 +
            flogtanh_00053_00007 +
            flogtanh_00147_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6344e71ca2b0fd39d36caedd889c3085 <=
            flogtanh_00000_00016 +
            flogtanh_00027_00006 +
            flogtanh_00148_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I0c99a68e0bed90afce18807acf7d55bb <=
            flogtanh_00001_00016 +
            flogtanh_00024_00006 +
            flogtanh_00149_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I1c95650979c86310ae2a949961c9db11 <=
            flogtanh_00002_00016 +
            flogtanh_00025_00006 +
            flogtanh_00150_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I04eaefa5d133e53494fc270b07be7043 <=
            flogtanh_00003_00016 +
            flogtanh_00026_00006 +
            flogtanh_00151_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4a64fa2412eb8058c2dfd9351d7b297d <=
            flogtanh_00006_00018 +
            flogtanh_00009_00005 +
            flogtanh_00023_00008 +
            flogtanh_00152_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie8bb2fcb752c6a33254963d1ebb4130d <=
            flogtanh_00007_00018 +
            flogtanh_00010_00005 +
            flogtanh_00020_00008 +
            flogtanh_00153_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Iac05b7e3ae18f948b72c356ccfb8000f <=
            flogtanh_00004_00018 +
            flogtanh_00011_00005 +
            flogtanh_00021_00008 +
            flogtanh_00154_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I27da3f75cca6c49e55db90306aa68e94 <=
            flogtanh_00005_00018 +
            flogtanh_00008_00005 +
            flogtanh_00022_00008 +
            flogtanh_00155_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Idc7fed723190098341225fe01ba65ced <=
            flogtanh_00002_00017 +
            flogtanh_00016_00004 +
            flogtanh_00156_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ife9065805598960919ee4f14c3cc6fd4 <=
            flogtanh_00003_00017 +
            flogtanh_00017_00004 +
            flogtanh_00157_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I717c5c2d6a2be61593492ae5f17a112f <=
            flogtanh_00000_00017 +
            flogtanh_00018_00004 +
            flogtanh_00158_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4c31fa8e6eb648439cdae1de1afe0d6f <=
            flogtanh_00001_00017 +
            flogtanh_00019_00004 +
            flogtanh_00159_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Iead549a9af27f1fced7d9c36e7b5c3f5 <=
            flogtanh_00011_00006 +
            flogtanh_00020_00009 +
            flogtanh_00029_00009 +
            flogtanh_00036_00007 +
            flogtanh_00160_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I10422eb79364e7d0e21e1643d9060331 <=
            flogtanh_00008_00006 +
            flogtanh_00021_00009 +
            flogtanh_00030_00009 +
            flogtanh_00037_00007 +
            flogtanh_00161_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I914cb87eba8baa40cd515334e59f26b2 <=
            flogtanh_00009_00006 +
            flogtanh_00022_00009 +
            flogtanh_00031_00009 +
            flogtanh_00038_00007 +
            flogtanh_00162_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I32ed679af4ab759901aee43c9d93eb67 <=
            flogtanh_00010_00006 +
            flogtanh_00023_00009 +
            flogtanh_00028_00009 +
            flogtanh_00039_00007 +
            flogtanh_00163_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Id376dfa5141402f4d41a8858180ed87e <=
            flogtanh_00006_00019 +
            flogtanh_00053_00008 +
            flogtanh_00164_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I98a384bc62ee03f5ad7df20ef2d9af95 <=
            flogtanh_00007_00019 +
            flogtanh_00054_00008 +
            flogtanh_00165_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Icfed259ca2bb2732d8e0c26ef67cd4cf <=
            flogtanh_00004_00019 +
            flogtanh_00055_00008 +
            flogtanh_00166_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I20861535c450d6e6bf11c45dac120454 <=
            flogtanh_00005_00019 +
            flogtanh_00052_00008 +
            flogtanh_00167_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I013929385ad819ddfcfcc59c22902ee3 <=
            flogtanh_00002_00018 +
            flogtanh_00020_00010 +
            flogtanh_00050_00006 +
            flogtanh_00168_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I34fffcb07fe82f11fe142f7c37f39155 <=
            flogtanh_00003_00018 +
            flogtanh_00021_00010 +
            flogtanh_00051_00006 +
            flogtanh_00169_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I61ca60fde05ed88cce714dcd8c13b827 <=
            flogtanh_00000_00018 +
            flogtanh_00022_00010 +
            flogtanh_00048_00006 +
            flogtanh_00170_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4907dd45c158dc7e0041c64f1fb388f6 <=
            flogtanh_00001_00018 +
            flogtanh_00023_00010 +
            flogtanh_00049_00006 +
            flogtanh_00171_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I2c8f6a9b9f655b317bb0af4d60fdbc4b <=
            flogtanh_00008_00007 +
            flogtanh_00028_00010 +
            flogtanh_00043_00006 +
            flogtanh_00172_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ic7dff631559304ec59f0696c66436d62 <=
            flogtanh_00009_00007 +
            flogtanh_00029_00010 +
            flogtanh_00040_00006 +
            flogtanh_00173_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6a239d3e55b4a9a3be9989a85bbec545 <=
            flogtanh_00010_00007 +
            flogtanh_00030_00010 +
            flogtanh_00041_00006 +
            flogtanh_00174_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I630f905e55f08e7d1569a08e937ad216 <=
            flogtanh_00011_00007 +
            flogtanh_00031_00010 +
            flogtanh_00042_00006 +
            flogtanh_00175_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8d13eb3669785c4279c685763d4f3fad <=
            flogtanh_00003_00019 +
            flogtanh_00049_00007 +
            flogtanh_00052_00009 +
            flogtanh_00176_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I25a6f3de9a9a01cbbdd32ed848561aa4 <=
            flogtanh_00000_00019 +
            flogtanh_00050_00007 +
            flogtanh_00053_00009 +
            flogtanh_00177_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Iba3dd4b2c2c85c4cfe770d9b52ef4634 <=
            flogtanh_00001_00019 +
            flogtanh_00051_00007 +
            flogtanh_00054_00009 +
            flogtanh_00178_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie1b744387b5200a504e4874e14d2f282 <=
            flogtanh_00002_00019 +
            flogtanh_00048_00007 +
            flogtanh_00055_00009 +
            flogtanh_00179_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Icf76cb69aedf4db01cd3444f4c4ba471 <=
            flogtanh_00005_00020 +
            flogtanh_00020_00011 +
            flogtanh_00047_00013 +
            flogtanh_00180_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4857b5b50556c8e7fff4b2d3e08e4b28 <=
            flogtanh_00006_00020 +
            flogtanh_00021_00011 +
            flogtanh_00044_00013 +
            flogtanh_00181_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I0a1e9cf99f1d4725327615f50fcc3ad0 <=
            flogtanh_00007_00020 +
            flogtanh_00022_00011 +
            flogtanh_00045_00013 +
            flogtanh_00182_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie844f4c446983ce381b0bc4c0e8ef7d7 <=
            flogtanh_00004_00020 +
            flogtanh_00023_00011 +
            flogtanh_00046_00013 +
            flogtanh_00183_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6067f47cccceea96ac46ff0d457b25f2 <=
            flogtanh_00000_00020 +
            flogtanh_00010_00008 +
            flogtanh_00030_00011 +
            flogtanh_00184_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ifd6fd1f3cbf8884ca7f64bc42278e4fa <=
            flogtanh_00001_00020 +
            flogtanh_00011_00008 +
            flogtanh_00031_00011 +
            flogtanh_00185_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Iaec9fd9e79371676bfa8ff14b4feae52 <=
            flogtanh_00002_00020 +
            flogtanh_00008_00008 +
            flogtanh_00028_00011 +
            flogtanh_00186_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I500757c4eda5d3d899aee47b87da585b <=
            flogtanh_00003_00020 +
            flogtanh_00009_00008 +
            flogtanh_00029_00011 +
            flogtanh_00187_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I47bf091b0fa74ad511a760bad9d2506c <=
            flogtanh_00043_00007 +
            flogtanh_00055_00010 +
            flogtanh_00188_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia4c3d0cd9957f678880de5775de76e0d <=
            flogtanh_00040_00007 +
            flogtanh_00052_00010 +
            flogtanh_00189_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          If5f957fa2f055b1c2c28e8d7cfe3e9ad <=
            flogtanh_00041_00007 +
            flogtanh_00053_00010 +
            flogtanh_00190_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3608378a5da8c66bef58528d56192530 <=
            flogtanh_00042_00007 +
            flogtanh_00054_00010 +
            flogtanh_00191_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie6dead855e00ea0a8e6a9b7503aaebb8 <=
            flogtanh_00007_00021 +
            flogtanh_00022_00012 +
            flogtanh_00046_00014 +
            flogtanh_00192_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3bae5e6862e003a8b9a476f72cc6858b <=
            flogtanh_00004_00021 +
            flogtanh_00023_00012 +
            flogtanh_00047_00014 +
            flogtanh_00193_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4431adecba8be9e5f21bc6b3e1f8cb10 <=
            flogtanh_00005_00021 +
            flogtanh_00020_00012 +
            flogtanh_00044_00014 +
            flogtanh_00194_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I21c7a2885126d532d00484376588a469 <=
            flogtanh_00006_00021 +
            flogtanh_00021_00012 +
            flogtanh_00045_00014 +
            flogtanh_00195_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I2c4d7339ff2fe68d060dd8d961dcab8c <=
            flogtanh_00003_00021 +
            flogtanh_00028_00012 +
            flogtanh_00050_00008 +
            flogtanh_00196_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Iee518b15b067eec58cccfa37f7432ea5 <=
            flogtanh_00000_00021 +
            flogtanh_00029_00012 +
            flogtanh_00051_00008 +
            flogtanh_00197_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I42145be9c2a80288ba4a2edd91f661a3 <=
            flogtanh_00001_00021 +
            flogtanh_00030_00012 +
            flogtanh_00048_00008 +
            flogtanh_00198_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I9dc297ad41fafcda77f5347f331cfc25 <=
            flogtanh_00002_00021 +
            flogtanh_00031_00012 +
            flogtanh_00049_00008 +
            flogtanh_00199_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I846700c79f30ca954cc2933fc94d355b <=
            flogtanh_00008_00009 +
            flogtanh_00043_00008 +
            flogtanh_00052_00011 +
            flogtanh_00200_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8af96a91457316e49e3f7dd5e57c82da <=
            flogtanh_00009_00009 +
            flogtanh_00040_00008 +
            flogtanh_00053_00011 +
            flogtanh_00201_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I7d1c247500d7d32e406b2a5f7e2b745b <=
            flogtanh_00010_00009 +
            flogtanh_00041_00008 +
            flogtanh_00054_00011 +
            flogtanh_00202_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I66d85c030a8864505298919046056305 <=
            flogtanh_00011_00009 +
            flogtanh_00042_00008 +
            flogtanh_00055_00011 +
            flogtanh_00203_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4841257ae596d9d3e4eb1e6f886956b0 <=
            flogtanh_00005_00022 +
            flogtanh_00021_00013 +
            flogtanh_00046_00015 +
            flogtanh_00204_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Icd6f7ec117f9ab4eda8c5eba41386ffa <=
            flogtanh_00006_00022 +
            flogtanh_00022_00013 +
            flogtanh_00047_00015 +
            flogtanh_00205_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ibc0498839d1d9b6dc853b8e5d7a88fa3 <=
            flogtanh_00007_00022 +
            flogtanh_00023_00013 +
            flogtanh_00044_00015 +
            flogtanh_00206_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
          I142ebca7f155e287e38ddf45423ab0fd <=
            flogtanh_00004_00022 +
            flogtanh_00020_00013 +
            flogtanh_00045_00015 +
            flogtanh_00207_00000 +
            {MAX_SUM_WDTH_L{1'h0}};
       end
   end







always_comb begin

            I5deafec6e5f32da1bcf8f7018cf794d8= I5033323484d90d6bfbe03749019fc6dd + I8cab6f6faf0758f26d1a8851fae43896;
            tout_00000_00000    = fgallag_final_00000_00000;

            I35b3fb2670f3a60d165c1fd10f02c00c= I5033323484d90d6bfbe03749019fc6dd + Ia3f7f07ddb09ea33218afe14281ac3c6;
            tout_00000_00001    = fgallag_final_00000_00001;

            I68925439e233444a4da44871f31de94a= I5033323484d90d6bfbe03749019fc6dd + Ie23ed3ee61f468f59f2baf661cb7f85d;
            tout_00000_00002    = fgallag_final_00000_00002;

            I3108702b5ca506422c1ba6174619f193= I5033323484d90d6bfbe03749019fc6dd + I79458089b042e181e37cc44c06d08681;
            tout_00000_00003    = fgallag_final_00000_00003;

            Icc8e8f6446ac64350a05f5e1e0541bb9= I5033323484d90d6bfbe03749019fc6dd + I856eada207c5006beb8f83f01d5d74c9;
            tout_00000_00004    = fgallag_final_00000_00004;

            Iadebaf3f6cca1ba78feab50ce70c8aef= I5033323484d90d6bfbe03749019fc6dd + I1ddfd31bbf062aa5c3c71d61e492e3a2;
            tout_00000_00005    = fgallag_final_00000_00005;

            I8681cf376dbeceab29279a7637249e7d= I5033323484d90d6bfbe03749019fc6dd + Ic5e0a84cf1a2ef907b2456559ea26c75;
            tout_00000_00006    = fgallag_final_00000_00006;

            Ie850a07565bed90389bb125ddcd39658= I5033323484d90d6bfbe03749019fc6dd + If367d63311c96726517240de13bd2a4b;
            tout_00000_00007    = fgallag_final_00000_00007;

            I97b77743c2311ec629ea24c933b60053= If5dad13ac41b3034bdb034bc86c9b348 + If49f97cc0c42b23ce393b534015559a0;
            tout_00001_00000    = fgallag_final_00001_00000;

            I07a0a8d41ed8176e92380f2c89c2afdd= If5dad13ac41b3034bdb034bc86c9b348 + I6c4ba0863ab4c8d1a56324a4d89ccbeb;
            tout_00001_00001    = fgallag_final_00001_00001;

            I021842328f948a94159b32903c8bcb68= If5dad13ac41b3034bdb034bc86c9b348 + I5a3297f48e1045273db6522744582b05;
            tout_00001_00002    = fgallag_final_00001_00002;

            Icaf3bd685005a05c8fb334266ea4e4b9= If5dad13ac41b3034bdb034bc86c9b348 + I326660e98f61bb2ced4c23c7bcc9324a;
            tout_00001_00003    = fgallag_final_00001_00003;

            I92d9e1d7dcf45a4d738c546e959687c3= If5dad13ac41b3034bdb034bc86c9b348 + Icdb143a4ce96029c2441758bf2edd7b0;
            tout_00001_00004    = fgallag_final_00001_00004;

            I39ca3a8ca714a9726114326ae6bfab0a= If5dad13ac41b3034bdb034bc86c9b348 + I3c6fb0df5846a19228a4e6cf9f9106ac;
            tout_00001_00005    = fgallag_final_00001_00005;

            Ie9ae20ed5b2a0cad2c37c5bb2ea05ff4= If5dad13ac41b3034bdb034bc86c9b348 + I6a3854ed571e8c262aa3ec377c247778;
            tout_00001_00006    = fgallag_final_00001_00006;

            I8f131eb6138c23fdcb35195703131e64= If5dad13ac41b3034bdb034bc86c9b348 + If19dc22d45cc4664c85a043ec4c00617;
            tout_00001_00007    = fgallag_final_00001_00007;

            Iff77e08da4bcbb85b95fa277b69653a9= Iac428f9f798618e1ef495c626c41892b + Ia7f53f0cd86055da72c13ac474f052a1;
            tout_00002_00000    = fgallag_final_00002_00000;

            I703e0a4879a39b3b8b0a49de86ca4ff4= Iac428f9f798618e1ef495c626c41892b + I0cbdfae6f75a639eb591d9c0022f5838;
            tout_00002_00001    = fgallag_final_00002_00001;

            I3da217f6f2d0f515bb9036673d753a88= Iac428f9f798618e1ef495c626c41892b + I1d0f031e8ae9c0335d501d1565118220;
            tout_00002_00002    = fgallag_final_00002_00002;

            Ifcc06d5a010e01a781ae8a9e9e2b31a0= Iac428f9f798618e1ef495c626c41892b + I4b66c202450986ef0df05e979cc8bc7f;
            tout_00002_00003    = fgallag_final_00002_00003;

            I42fd611fec087113ba6e35f281bced9c= Iac428f9f798618e1ef495c626c41892b + I972bee4216f8e532e8fa4bd25fbb9c57;
            tout_00002_00004    = fgallag_final_00002_00004;

            I5bb626e7347bb9ae4219cc72244b38f8= Iac428f9f798618e1ef495c626c41892b + I1182655739d7ab5bbe4a6546a5ca36fd;
            tout_00002_00005    = fgallag_final_00002_00005;

            I47e2dac0068652338f94ddffd2dbe88a= Iac428f9f798618e1ef495c626c41892b + I195c3a82123142d509886ee37dc6fc98;
            tout_00002_00006    = fgallag_final_00002_00006;

            I59a3f06de2984078a4d4c430a2980fe3= Iac428f9f798618e1ef495c626c41892b + I96ef4b631a7f63e19f67f3920685f0e6;
            tout_00002_00007    = fgallag_final_00002_00007;

            I857b7fd58279b1063a06a4f33b880ba6= I5a6427c8f18b36d2ea18fe60a0831ef1 + I5f68368511b59d2e365cc91b806b334e;
            tout_00003_00000    = fgallag_final_00003_00000;

            I3901bbda029cd0a41640001c1efd400f= I5a6427c8f18b36d2ea18fe60a0831ef1 + Ia6255a136d5f36ea6cba654bd5823850;
            tout_00003_00001    = fgallag_final_00003_00001;

            Ifceeccf10f1d85a32f70c04654a1a1b4= I5a6427c8f18b36d2ea18fe60a0831ef1 + I21594c8b0169efd7c2aa6cbc31f4a901;
            tout_00003_00002    = fgallag_final_00003_00002;

            I2d810c1d1304658edff74921e8d0f388= I5a6427c8f18b36d2ea18fe60a0831ef1 + Ife123bf57fe693dabe6aeaa236c4e058;
            tout_00003_00003    = fgallag_final_00003_00003;

            I575b0201be445388607ab83465eab8d6= I5a6427c8f18b36d2ea18fe60a0831ef1 + I518a2736384c14c02f27bfa3d8ea7aff;
            tout_00003_00004    = fgallag_final_00003_00004;

            I7928c5ce0f821df1cb6271d15e19fa22= I5a6427c8f18b36d2ea18fe60a0831ef1 + I2dcc0d17b9fcac35693bf32b5c5540fd;
            tout_00003_00005    = fgallag_final_00003_00005;

            I12695a21c942d02a432cf6382d7d7452= I5a6427c8f18b36d2ea18fe60a0831ef1 + Ic0819ccefe784a6379716b3633ae0196;
            tout_00003_00006    = fgallag_final_00003_00006;

            I00d03f0f71b008dad8035bbf251f41bf= I5a6427c8f18b36d2ea18fe60a0831ef1 + Ia540866403683bc30504bace19bdda7b;
            tout_00003_00007    = fgallag_final_00003_00007;

            I41afedcbc0f492e3243436cbefdaf609= Icc29441eac6ca7a138d45743d37505e3 + I915054f2fbb8b93516d8748a3e3e29e2;
            tout_00004_00000    = fgallag_final_00004_00000;

            I638c4c2708e437a050ed7cbbac516a59= Icc29441eac6ca7a138d45743d37505e3 + I42460fae0acff25fa2b829e39ddcc4fd;
            tout_00004_00001    = fgallag_final_00004_00001;

            I6877d3306b1f08c236b5d1b59f0de259= Icc29441eac6ca7a138d45743d37505e3 + I77a94cd9186ca546ca9664942ea3537f;
            tout_00004_00002    = fgallag_final_00004_00002;

            Ib3e66aa460f39d32110ea6f115785b3d= Icc29441eac6ca7a138d45743d37505e3 + I9a5388f8aa6e9924a309aa8db4c1983b;
            tout_00004_00003    = fgallag_final_00004_00003;

            I5e603e8392a5322951b3225b65b19446= Icc29441eac6ca7a138d45743d37505e3 + I3a76f70ca3bfbcacc6f3342aa71f1912;
            tout_00004_00004    = fgallag_final_00004_00004;

            If5da7fa1a615e1122445460e33487772= Icc29441eac6ca7a138d45743d37505e3 + I46e9c76b19ed1ff21f102efe6ee5c732;
            tout_00004_00005    = fgallag_final_00004_00005;

            Ic4153dafafaf7d047478c5d81109437f= Icc29441eac6ca7a138d45743d37505e3 + I3096d11098113da669ee0a94686e600d;
            tout_00004_00006    = fgallag_final_00004_00006;

            I7b5476007f04e81afc0125e6a8930303= Icc29441eac6ca7a138d45743d37505e3 + Ie6764a631310e312ba5c2c1e601d828f;
            tout_00004_00007    = fgallag_final_00004_00007;

            I3521a18022925249caddb8e37d2c1262= Icc29441eac6ca7a138d45743d37505e3 + Icc6d895d943e14f2801c22e79ce190e8;
            tout_00004_00008    = fgallag_final_00004_00008;

            Ifd0f52d4f814e2bb4c3bd34c1e09bda7= Icc29441eac6ca7a138d45743d37505e3 + I9b09b800a9dcd8ac36f25cb0324e748d;
            tout_00004_00009    = fgallag_final_00004_00009;

            I8945f6d420c8b373225451defcd2c805= I0e7754dcbc04a4850e052ae4a2fbe328 + I71e4d98dca37256fcc84248a26d703e2;
            tout_00005_00000    = fgallag_final_00005_00000;

            Ieec6cb6518cc0d9300de0c4f2d32487d= I0e7754dcbc04a4850e052ae4a2fbe328 + Ic6fa98631d742b27f252fe7c95caef55;
            tout_00005_00001    = fgallag_final_00005_00001;

            Ic62eb7e90d703ef994e68587345a4293= I0e7754dcbc04a4850e052ae4a2fbe328 + I20c65000bbc10299168af7390776a03c;
            tout_00005_00002    = fgallag_final_00005_00002;

            Id3efd8419da986aa89b8ad8e75848cfa= I0e7754dcbc04a4850e052ae4a2fbe328 + I66a304016a9adfd85a2abb6f8fd39afc;
            tout_00005_00003    = fgallag_final_00005_00003;

            I40803f10b7c4dc9ae4969739349b0265= I0e7754dcbc04a4850e052ae4a2fbe328 + Ib303ea0240e7ab5f000dd10e975b2274;
            tout_00005_00004    = fgallag_final_00005_00004;

            I7d961743fdeaf1e72e4b25c12a1d4c46= I0e7754dcbc04a4850e052ae4a2fbe328 + I5dfc71255cba279420b7545df4d35c40;
            tout_00005_00005    = fgallag_final_00005_00005;

            Ifea156f33eb61fece272efe379327f6e= I0e7754dcbc04a4850e052ae4a2fbe328 + I02330ade2eed926076cc071e45eed82c;
            tout_00005_00006    = fgallag_final_00005_00006;

            Ifc99169b3399f3d14121c1a9bce3fc21= I0e7754dcbc04a4850e052ae4a2fbe328 + Iae9e023628eb6686708b2656f15616cc;
            tout_00005_00007    = fgallag_final_00005_00007;

            I6536144383cbda6f3b3c564391866906= I0e7754dcbc04a4850e052ae4a2fbe328 + Ibf482db0f5058be72061267c42ebc292;
            tout_00005_00008    = fgallag_final_00005_00008;

            Ic21bf9a8a4cd85ec123d7fe142ed49c0= I0e7754dcbc04a4850e052ae4a2fbe328 + Iebdf938a28594624f4d4a337356485cb;
            tout_00005_00009    = fgallag_final_00005_00009;

            I1f31fe6a0ca8510bcadbc2069403150b= Ia30c019ed8ce395556494a92e7b42a92 + I6ecf7249e6151477fe74a79d0b126b21;
            tout_00006_00000    = fgallag_final_00006_00000;

            I0e40933d00f4a7d9b53b2764aa0da700= Ia30c019ed8ce395556494a92e7b42a92 + I737daf208eccf95feb3192897586cdce;
            tout_00006_00001    = fgallag_final_00006_00001;

            Ic41a6e00bc84bfc1b8194d15bb899c93= Ia30c019ed8ce395556494a92e7b42a92 + Icfc1c6d96a3598af73e99a350c387d72;
            tout_00006_00002    = fgallag_final_00006_00002;

            I2832571f2b0a7fbb41d2e8ca7f64e003= Ia30c019ed8ce395556494a92e7b42a92 + Ie3e0c0e40c7a67ce7f957e74bd2a895d;
            tout_00006_00003    = fgallag_final_00006_00003;

            I9593c853e41952e408a809cb24efa4fd= Ia30c019ed8ce395556494a92e7b42a92 + I847cf7ff866f8a666872c12d6b67b1b1;
            tout_00006_00004    = fgallag_final_00006_00004;

            I6edffbf4136e193dca0fcec3a74e8e9c= Ia30c019ed8ce395556494a92e7b42a92 + I954ff0f9ee871a31774a3d786128fa13;
            tout_00006_00005    = fgallag_final_00006_00005;

            Ibaed50cc2e36ae58945887d11a6ec9e4= Ia30c019ed8ce395556494a92e7b42a92 + If8b0b96a659183e3651c691a2848b86b;
            tout_00006_00006    = fgallag_final_00006_00006;

            Ie4570cac44f59e6ff46f73a703026479= Ia30c019ed8ce395556494a92e7b42a92 + I7168b0efdd2fae57292379c9d15c62eb;
            tout_00006_00007    = fgallag_final_00006_00007;

            Ibaa136d37936687e9dbe4222749d19c3= Ia30c019ed8ce395556494a92e7b42a92 + I9e2de71442b8f504358e582087a6d19f;
            tout_00006_00008    = fgallag_final_00006_00008;

            If85de3225f45478827b43b89089cd29e= Ia30c019ed8ce395556494a92e7b42a92 + I3e265a7dcf29687248b9275df49771fb;
            tout_00006_00009    = fgallag_final_00006_00009;

            I0344b86a6e9c036e103a9c1f3651175f= I9799695ea8244992a6694eaf5c8ae64d + Ie932a22a7f1fa37087cbc9e8d73efef4;
            tout_00007_00000    = fgallag_final_00007_00000;

            I5463d13575e0b9fb8a0f6cc8b35d0ce9= I9799695ea8244992a6694eaf5c8ae64d + I0c0d844fe3b7d35c1ed6bd7cc4e0dc24;
            tout_00007_00001    = fgallag_final_00007_00001;

            I8a3c63ef122001a29e5abe93c4e1a48f= I9799695ea8244992a6694eaf5c8ae64d + Idc77c7d5123717fc2596a51d904c6d82;
            tout_00007_00002    = fgallag_final_00007_00002;

            I6a79108484fcb192f6d93bfb98e271c4= I9799695ea8244992a6694eaf5c8ae64d + I07048dc5cbe24ff72d24902d572face0;
            tout_00007_00003    = fgallag_final_00007_00003;

            I9001e95b71457a2bd09a9846af370b16= I9799695ea8244992a6694eaf5c8ae64d + I79a46279070c53678a5af54f661c5821;
            tout_00007_00004    = fgallag_final_00007_00004;

            I51620de618db6327358a5cac97e1e97f= I9799695ea8244992a6694eaf5c8ae64d + I5e8ecdbb018402b2fbc0049ee44bae8c;
            tout_00007_00005    = fgallag_final_00007_00005;

            Ib9c58818059af5c5a03e77a5dcef4654= I9799695ea8244992a6694eaf5c8ae64d + I9aab16e89f1b64117caece8ca8af5940;
            tout_00007_00006    = fgallag_final_00007_00006;

            I8081c71aa01a8d575bfea6ea7f2f595f= I9799695ea8244992a6694eaf5c8ae64d + I8110a5a62607093b21b7cd088b1d9ee0;
            tout_00007_00007    = fgallag_final_00007_00007;

            Iad999607ad8d7da0f3b341f83ea030a6= I9799695ea8244992a6694eaf5c8ae64d + I05fb1982415bd3fa78dd9a00af7a3d4a;
            tout_00007_00008    = fgallag_final_00007_00008;

            Ie7291c914d2cb66f547b0a7717f71311= I9799695ea8244992a6694eaf5c8ae64d + Ia9f375709014a9d553d46cff2799b59f;
            tout_00007_00009    = fgallag_final_00007_00009;

            Ic01018a5f1bc392bbd267016f6612a83= I4524cd664b4cb41f642c675fa484c84b + I3753b2c4ba8f1bee70def390a96586b0;
            tout_00008_00000    = fgallag_final_00008_00000;

            Ib11dff839e7e532657b32f29fd9b1651= I4524cd664b4cb41f642c675fa484c84b + I4dbd1bb8f1641f15e3a4f1e309962811;
            tout_00008_00001    = fgallag_final_00008_00001;

            I251d7ea16dd5407d22a6846ddcfe12d8= I4524cd664b4cb41f642c675fa484c84b + I29c8133231cfda17668bbe7b692bdfe2;
            tout_00008_00002    = fgallag_final_00008_00002;

            I773797f81f73b9b6e844441142a1bb48= I4524cd664b4cb41f642c675fa484c84b + I779da979707d9712c1626d6025f97599;
            tout_00008_00003    = fgallag_final_00008_00003;

            I853ecadf30fc10a13dd1ffb1f2dfb5d6= I4524cd664b4cb41f642c675fa484c84b + I09a1d04c307fcb8a0e30925d86df3fe9;
            tout_00008_00004    = fgallag_final_00008_00004;

            Ibb8b3c91e1d3b890cfe58f32f8ec3ae3= I4524cd664b4cb41f642c675fa484c84b + I2cefbf897bb7f6f67ca500727e85c683;
            tout_00008_00005    = fgallag_final_00008_00005;

            I3485d69de942d64e56925da522175b51= I4524cd664b4cb41f642c675fa484c84b + I74ac0327175f50f508a5013df298df02;
            tout_00008_00006    = fgallag_final_00008_00006;

            Iae42f12bc0475c8b58341d80027a57cb= I4524cd664b4cb41f642c675fa484c84b + Ifebfa58419ecd22a334ed4b67f5c3581;
            tout_00008_00007    = fgallag_final_00008_00007;

            I22fe2af25463f87ee7315a9aac32854e= I64e959d80af111ed2fcd54a5407d21bf + I2956687a5fc2fba7149889624ef85647;
            tout_00009_00000    = fgallag_final_00009_00000;

            Idf44ad78c338c39699721ce511691dfd= I64e959d80af111ed2fcd54a5407d21bf + I088898ee932a96c14f2f0f568f5455b6;
            tout_00009_00001    = fgallag_final_00009_00001;

            I984a657f9265d41318c0290e249e9712= I64e959d80af111ed2fcd54a5407d21bf + I2d9632ae6a0f3ba44c3da8f56ba3fedf;
            tout_00009_00002    = fgallag_final_00009_00002;

            I915fccfb1d1ada9aa7c8e24c2eebd04c= I64e959d80af111ed2fcd54a5407d21bf + I3c0ddec25c53c166d30eb78d4518840e;
            tout_00009_00003    = fgallag_final_00009_00003;

            I2bdf58ecd0974720631be830efb48dc8= I64e959d80af111ed2fcd54a5407d21bf + I296bc392d4223cbdd6f77be6523df819;
            tout_00009_00004    = fgallag_final_00009_00004;

            Ibaedf6246fa43acc8accb5a24d49cc2f= I64e959d80af111ed2fcd54a5407d21bf + I05028975b49ec0c089bd981696f85a8b;
            tout_00009_00005    = fgallag_final_00009_00005;

            I904d13524dcdf55478a5266d50e53ff7= I64e959d80af111ed2fcd54a5407d21bf + I3fd068d55154441ffd005999ea823fd0;
            tout_00009_00006    = fgallag_final_00009_00006;

            I22d8e5d57c1bc082169437a654d22bba= I64e959d80af111ed2fcd54a5407d21bf + I066cd52173ec5dbce9a3f470d73325af;
            tout_00009_00007    = fgallag_final_00009_00007;

            I719cdaa2a2e61a0df7f1fd5efe517426= I3e0da4bcbab4804b5397fb3aa2c94f51 + If257757fa31c2f4cc9ec322e4ecccf83;
            tout_00010_00000    = fgallag_final_00010_00000;

            I8e92a61eb73c41680652936cfcc614ff= I3e0da4bcbab4804b5397fb3aa2c94f51 + I2b9584392ef9a7828ff57bd4c522a302;
            tout_00010_00001    = fgallag_final_00010_00001;

            I7ad5af8319f6da469858300f0777b580= I3e0da4bcbab4804b5397fb3aa2c94f51 + Id3670a6f05d40ab69624544de92b9c64;
            tout_00010_00002    = fgallag_final_00010_00002;

            I32be72eaf04e79120a57ea94296a4e56= I3e0da4bcbab4804b5397fb3aa2c94f51 + Ia840e19ca36795a50ab1a6e6a1729edb;
            tout_00010_00003    = fgallag_final_00010_00003;

            Ie756f6a87d85adb40479ce7cf3545556= I3e0da4bcbab4804b5397fb3aa2c94f51 + I87d958c00fc6209d901147831b0c951c;
            tout_00010_00004    = fgallag_final_00010_00004;

            I8794c6ce0a3f2e6697372e2c911ba420= I3e0da4bcbab4804b5397fb3aa2c94f51 + I1abb512ca0383c9e7104418e07281841;
            tout_00010_00005    = fgallag_final_00010_00005;

            Ic82b1a29b5e63bcc3686a0d4bf1f5c24= I3e0da4bcbab4804b5397fb3aa2c94f51 + Iffd94cf3a8a4681ff3327c90bf89bd8b;
            tout_00010_00006    = fgallag_final_00010_00006;

            I253ef976058080beab79646af18e2d5b= I3e0da4bcbab4804b5397fb3aa2c94f51 + Ifb8b3586a5b69b20cf03eabf51344ab6;
            tout_00010_00007    = fgallag_final_00010_00007;

            I930dd54c36540d75dc870eef89960163= I3740b30d31f3c61d93a14a46e3199c4d + Ib8380902ac4082f834744ddef6d0cc6a;
            tout_00011_00000    = fgallag_final_00011_00000;

            Iaf7554cd4e8b5ea6155ec61a8d589b86= I3740b30d31f3c61d93a14a46e3199c4d + I25aefb53f59a00abe88b9dcf6be6907a;
            tout_00011_00001    = fgallag_final_00011_00001;

            I50907c7d1efa0038d81efed82b192891= I3740b30d31f3c61d93a14a46e3199c4d + Iab6d0f72579687407e029c630b107f7d;
            tout_00011_00002    = fgallag_final_00011_00002;

            If3e9486d2960d164d94641d4f1917416= I3740b30d31f3c61d93a14a46e3199c4d + I523e9b6f828ec7f166750112f8a3f676;
            tout_00011_00003    = fgallag_final_00011_00003;

            I2bec61db45dd79b98d6ebff6c5a4899e= I3740b30d31f3c61d93a14a46e3199c4d + I343df614f97cf732e57cf2ad3f95dc9e;
            tout_00011_00004    = fgallag_final_00011_00004;

            I7f31647f3ea6ce7bbd211c25cf4828fb= I3740b30d31f3c61d93a14a46e3199c4d + I0c4bbd1827b1859caabb067e864ce4b3;
            tout_00011_00005    = fgallag_final_00011_00005;

            Ice65387e606faf9c7b884475b489abba= I3740b30d31f3c61d93a14a46e3199c4d + I34d428a56bd0142a9be9f627f1c3c87f;
            tout_00011_00006    = fgallag_final_00011_00006;

            I63f914927dcf49552e9f3fe0180a30e8= I3740b30d31f3c61d93a14a46e3199c4d + Ice66c108aa66981051df71e226cb0e4d;
            tout_00011_00007    = fgallag_final_00011_00007;

            I742ff5725e3a18acd03454cf9f313f4b= Ibf0a30abfec9031737eada436ac1a0d4 + I6c1235e88ae444a96ea64fd1bfd04d8f;
            tout_00012_00000    = fgallag_final_00012_00000;

            I84e4b3bc63ec0b0bff7f98f433c1fd67= Ibf0a30abfec9031737eada436ac1a0d4 + Ie2c801b2de066c3218d7312615b7bfda;
            tout_00012_00001    = fgallag_final_00012_00001;

            I78c6a1428a1f211c5e89b8c76b3dc033= Ibf0a30abfec9031737eada436ac1a0d4 + I7d98d1e5f07fccff5f20eaca6363c700;
            tout_00012_00002    = fgallag_final_00012_00002;

            I9897cbf9d7cab759f99f5f8f4bc125d0= Ibf0a30abfec9031737eada436ac1a0d4 + Iab3876e5107e3a56b1fafe41e16d9482;
            tout_00012_00003    = fgallag_final_00012_00003;

            I9a6c1ff6dde5141849e4aa925140ebb8= Ibf0a30abfec9031737eada436ac1a0d4 + Ica807adc510a2e32580ca77c18ea0b45;
            tout_00012_00004    = fgallag_final_00012_00004;

            Icc1c25b229393361f1245c40f573b423= Ibf0a30abfec9031737eada436ac1a0d4 + I31f6bbfbbbd4c20d0c5c71663da1d4c1;
            tout_00012_00005    = fgallag_final_00012_00005;

            I53b5a72e41ee53037ee3ae040799f401= Ibf0a30abfec9031737eada436ac1a0d4 + Ie4e4eaf3e5d2f581210af8054df71c6c;
            tout_00012_00006    = fgallag_final_00012_00006;

            I3cc25fb583118f45babf457fe78d5434= Ibf0a30abfec9031737eada436ac1a0d4 + I220f8e45e5fe6e69f02cded87f12e1e5;
            tout_00012_00007    = fgallag_final_00012_00007;

            I20c046dd8a1265e12e902275b73417da= Ibf0a30abfec9031737eada436ac1a0d4 + If47be2ca4617a426258c51f8d977ba3f;
            tout_00012_00008    = fgallag_final_00012_00008;

            I1b184c9a34aeb6eda813d86556e235d9= Ibf0a30abfec9031737eada436ac1a0d4 + I71a28e8525f07dabeabe4b4f45f353d0;
            tout_00012_00009    = fgallag_final_00012_00009;

            I70e03db993e1d26d5814ff5fcd38ada1= Id36e8953a02400a5ab1f4dfdb0422e6d + I22c3140a8db02352d2e2a2a11eeba117;
            tout_00013_00000    = fgallag_final_00013_00000;

            I119dc168a44950d215af877eb81152fe= Id36e8953a02400a5ab1f4dfdb0422e6d + I15022e1b349eee259d3567837283dbf6;
            tout_00013_00001    = fgallag_final_00013_00001;

            Id717ed42457eb1d3f4e3edbf0dd72c41= Id36e8953a02400a5ab1f4dfdb0422e6d + I79259217f63b2f6263552c434d0e5c93;
            tout_00013_00002    = fgallag_final_00013_00002;

            I79d1f852a03bcc11d6121a12d8c5b86d= Id36e8953a02400a5ab1f4dfdb0422e6d + Ief76663994991118b1899ea4ddf4527d;
            tout_00013_00003    = fgallag_final_00013_00003;

            I769e650e49f152c0803b06232740691c= Id36e8953a02400a5ab1f4dfdb0422e6d + I9470c7ab9634c01bb832c9e4ff5496bf;
            tout_00013_00004    = fgallag_final_00013_00004;

            I1ef3c09b8481f14c3526224430a5f4b9= Id36e8953a02400a5ab1f4dfdb0422e6d + I06d859184884c07a14c83d2f06587ad5;
            tout_00013_00005    = fgallag_final_00013_00005;

            I2a38d43a7e25050aa672cbf84a409aa8= Id36e8953a02400a5ab1f4dfdb0422e6d + Ie02de90d8eb06b16314946d21299500c;
            tout_00013_00006    = fgallag_final_00013_00006;

            I1c2be5e13c462a8a6b07bca311582ce4= Id36e8953a02400a5ab1f4dfdb0422e6d + If4b100d26126e460c41b8c1bc8fbbb96;
            tout_00013_00007    = fgallag_final_00013_00007;

            Ie8fd61caf16aa0e504cc7dc8cec6f0b8= Id36e8953a02400a5ab1f4dfdb0422e6d + Ife732309efcc740cfff5c747aab2e3d6;
            tout_00013_00008    = fgallag_final_00013_00008;

            Icd0fe98ca873ad6dacdf80dfdfc450ec= Id36e8953a02400a5ab1f4dfdb0422e6d + Ic7ad59f6a232a997706d17b4098e0324;
            tout_00013_00009    = fgallag_final_00013_00009;

            I94e1ab698dc93ff0764dc5c1e62179fe= Ica71108a53bfcfd1892b4d03ef68110c + I26781ef851ed43c6f88ff1215cddca6b;
            tout_00014_00000    = fgallag_final_00014_00000;

            Ifd48363af9abb390a72991fbdd6f7877= Ica71108a53bfcfd1892b4d03ef68110c + I68e58664be09261e5a80d6f8ecdd1b60;
            tout_00014_00001    = fgallag_final_00014_00001;

            I44f79397a010088e4ecdcb9669f2efbd= Ica71108a53bfcfd1892b4d03ef68110c + I97aede8502e443f98938487a5a5c072c;
            tout_00014_00002    = fgallag_final_00014_00002;

            I124b0b7d91cfb42b0d9722f3229c2d53= Ica71108a53bfcfd1892b4d03ef68110c + I177be24718c59688752097fe2a4085c4;
            tout_00014_00003    = fgallag_final_00014_00003;

            Iadf1875c584adc34f7586a146184a763= Ica71108a53bfcfd1892b4d03ef68110c + I5971253546899e9a82f387d5eabcc7b3;
            tout_00014_00004    = fgallag_final_00014_00004;

            I02d3f9982f02ea85f996bf5b5975b930= Ica71108a53bfcfd1892b4d03ef68110c + Ic75b8bbb1b80001ec188a0cd25623420;
            tout_00014_00005    = fgallag_final_00014_00005;

            Ia6e1b39d83ddce053518c5ae9a5ca33e= Ica71108a53bfcfd1892b4d03ef68110c + Idb0a98cea3ee6cd4308bfc2414a003e1;
            tout_00014_00006    = fgallag_final_00014_00006;

            I3308663053f4307d43ac66f43266f706= Ica71108a53bfcfd1892b4d03ef68110c + Ibe502ebbb366f54a8f8fda4e361308e3;
            tout_00014_00007    = fgallag_final_00014_00007;

            I87ad25dff6c0c9ac46b7a129cb575537= Ica71108a53bfcfd1892b4d03ef68110c + I00ff1331b1900bb031ee81d2a58c1bd5;
            tout_00014_00008    = fgallag_final_00014_00008;

            Ibf5d40b7c46b50866f58f6fa23e1861b= Ica71108a53bfcfd1892b4d03ef68110c + I9ea09f27ce4484f2e7fc3a6b6d6ecb7c;
            tout_00014_00009    = fgallag_final_00014_00009;

            I0e3a9a3b38875156d15f697adaf95410= I7c97629ec6e594f9b2160815ddd133cc + Ide0abde3644a4fafb436aa59768d016e;
            tout_00015_00000    = fgallag_final_00015_00000;

            Ie3f87d094e71e4a82f60e8d91cdd768b= I7c97629ec6e594f9b2160815ddd133cc + I9858bb2a3cc458aca5bf7eb077ee55dd;
            tout_00015_00001    = fgallag_final_00015_00001;

            I793f52d174cd09fe000e8d0351753592= I7c97629ec6e594f9b2160815ddd133cc + I98bbe3b75958f10195dee6460cf2aca6;
            tout_00015_00002    = fgallag_final_00015_00002;

            I89ea3da7db40e7e6705020462b2d1df1= I7c97629ec6e594f9b2160815ddd133cc + I491f2373b2df19a4c22e1787ef034179;
            tout_00015_00003    = fgallag_final_00015_00003;

            Ib2af2f1a928dd824f25b99f0b602753f= I7c97629ec6e594f9b2160815ddd133cc + I9e45e3d7117ce48cdbfc5db8c0ccfcf4;
            tout_00015_00004    = fgallag_final_00015_00004;

            Ie3e887f5f1a64c37a10404d636212b45= I7c97629ec6e594f9b2160815ddd133cc + Ibadcb205c7e9a0f3345cac7eb41b5985;
            tout_00015_00005    = fgallag_final_00015_00005;

            I5c6a004278f155d33d0cc1b576c3b25f= I7c97629ec6e594f9b2160815ddd133cc + I31b0f2fe98cfddbc05dbd14be8be394b;
            tout_00015_00006    = fgallag_final_00015_00006;

            I6a03a4a548a0906d1a3e9ce47f3454c6= I7c97629ec6e594f9b2160815ddd133cc + I8b611f7c12ddd81de403ba74e212857f;
            tout_00015_00007    = fgallag_final_00015_00007;

            I542e525074d049197ac3904e6102f0bd= I7c97629ec6e594f9b2160815ddd133cc + I004c98da87996b77b5761d366210f782;
            tout_00015_00008    = fgallag_final_00015_00008;

            Ie0307a43ce71ba73d4c8e5ad556bd341= I7c97629ec6e594f9b2160815ddd133cc + I645ff0d8c0a87ba7f792fc83f342b958;
            tout_00015_00009    = fgallag_final_00015_00009;

            Ib03e1d3a1f27721e4ea32629c2e86f85= I4823c8239ace86dc399e906c1b5a0d74 + If91268e2b84df18785cd6a53e53eb4e9;
            tout_00016_00000    = fgallag_final_00016_00000;

            I782f4ab4666c9f550a2cfc943cedbe77= I4823c8239ace86dc399e906c1b5a0d74 + Ia349e1f7c10a63ddccb3f300c73b4572;
            tout_00016_00001    = fgallag_final_00016_00001;

            Ib991e16161d5c8b3b655e3c7c08b93c4= I4823c8239ace86dc399e906c1b5a0d74 + I977864efb0d94149cce7dc4d165f11de;
            tout_00016_00002    = fgallag_final_00016_00002;

            I72f8c6bad4bff3b00055aa8824479931= I4823c8239ace86dc399e906c1b5a0d74 + I5f3ff7fa8686f7a380302d71b88cfb4b;
            tout_00016_00003    = fgallag_final_00016_00003;

            I58e5100cc1e9b809e93125fe5d08a9d8= I10ad572ca72c2ea991487c39f7eabd7b + I9570f8498d95bee230bb3c5e720bb857;
            tout_00017_00000    = fgallag_final_00017_00000;

            I0aa7056fdacd6022f328a3be49048856= I10ad572ca72c2ea991487c39f7eabd7b + I08581dc8d42be712cfb36d744f2786e0;
            tout_00017_00001    = fgallag_final_00017_00001;

            Ia2f40b5c49a2284fb6a234bf7472130f= I10ad572ca72c2ea991487c39f7eabd7b + Ieb664ac9be65fba2e25960141f7fb4b6;
            tout_00017_00002    = fgallag_final_00017_00002;

            I8da184aee7953890f2c89e40744402f4= I10ad572ca72c2ea991487c39f7eabd7b + Ic01904f7c518990eff2dc1de127676c4;
            tout_00017_00003    = fgallag_final_00017_00003;

            I613ccfc7dad5627cde02fa1720244d01= Ie9f3fd3a6d16316e55addbe0e336519f + I9b919f3d4ee3f33506b87bcdaf2d43a3;
            tout_00018_00000    = fgallag_final_00018_00000;

            I080fc6c99e506e569b97433f3fdc3e60= Ie9f3fd3a6d16316e55addbe0e336519f + Id09b8242c22851fb960d55222fe733d4;
            tout_00018_00001    = fgallag_final_00018_00001;

            I79aa118ef8ac0d9b13723fb1f5a7e4ad= Ie9f3fd3a6d16316e55addbe0e336519f + I6d2dbb953a58b91dafa7f0d34d41bdc3;
            tout_00018_00002    = fgallag_final_00018_00002;

            I7e6e7601245ca5b3a58b91848e25a6d3= Ie9f3fd3a6d16316e55addbe0e336519f + I43f2ddd9780f86af489f8deae51168ec;
            tout_00018_00003    = fgallag_final_00018_00003;

            I2792edda66743635b837aa3bec0c58b9= I07965bca84276dd56da1af98e64b0adc + Iebf28886bd39c2540c90e808a9c20d3d;
            tout_00019_00000    = fgallag_final_00019_00000;

            I085cc29465c945957d00cbcf804e3ae4= I07965bca84276dd56da1af98e64b0adc + I954dd66f60316803a8f13a39c460a39a;
            tout_00019_00001    = fgallag_final_00019_00001;

            I74a8e879666bb216a331fd2ab723e37c= I07965bca84276dd56da1af98e64b0adc + I1fb13d7500f5ac3821c424bd3688cf4e;
            tout_00019_00002    = fgallag_final_00019_00002;

            I7a90a43ed71e82862457d9fa40bd005c= I07965bca84276dd56da1af98e64b0adc + I0a013fff6c792363bd7feb03d9691db8;
            tout_00019_00003    = fgallag_final_00019_00003;

            Ie1e7b4bd6201baa02b8d59cb0f6ffb8e= Ic2ade31b8bcf68c4dcc1a371ff14074b + Ia072f1d679429d3c3180f8eb67fc7dd7;
            tout_00020_00000    = fgallag_final_00020_00000;

            Ib7b7cdc22b22f276b1c021abaa8fb443= Ic2ade31b8bcf68c4dcc1a371ff14074b + I37b3988d699a1ed42923e3fd1584ecc0;
            tout_00020_00001    = fgallag_final_00020_00001;

            Ib58e33f31be36b28997ba05ef1004573= Ic2ade31b8bcf68c4dcc1a371ff14074b + I7e66a42eb7cdb820cd1297c39f0625e8;
            tout_00020_00002    = fgallag_final_00020_00002;

            Ibec394e82f499e8d2d5a9524f943d6ac= Ic2ade31b8bcf68c4dcc1a371ff14074b + I79e3e49f57d47231c0fe6aaafdbc57f1;
            tout_00020_00003    = fgallag_final_00020_00003;

            Ie06ad127e475dc131859992bb5f350a0= Ic2ade31b8bcf68c4dcc1a371ff14074b + I9362b615a612599239e3b752a9334e8c;
            tout_00020_00004    = fgallag_final_00020_00004;

            Ic494a58468b6a7dda76923a9475bf173= Ic2ade31b8bcf68c4dcc1a371ff14074b + I7cf8401bf6893eab0b9f33a0f91ddd05;
            tout_00020_00005    = fgallag_final_00020_00005;

            Ib82a2db86d03fe8538fa19d06e501dae= Ic0edcf240048fbfde4e938c3e4c5e281 + I55c425102db0a6838012a165c0597680;
            tout_00021_00000    = fgallag_final_00021_00000;

            I5b64727fee9d0825a4ea83261992e489= Ic0edcf240048fbfde4e938c3e4c5e281 + I50c4e1d3a3f63b93bc36b5141226fb3c;
            tout_00021_00001    = fgallag_final_00021_00001;

            Ice7e502b9c2b797719448fde8376087a= Ic0edcf240048fbfde4e938c3e4c5e281 + Ief96603d41b4f670d2bbfa3d3875c903;
            tout_00021_00002    = fgallag_final_00021_00002;

            I792b4f73ed7139b8761443cbc0833e39= Ic0edcf240048fbfde4e938c3e4c5e281 + Idc7df6877bdb7e7d392307d78183d31c;
            tout_00021_00003    = fgallag_final_00021_00003;

            I278d57d1964cbf3339db450926ef4782= Ic0edcf240048fbfde4e938c3e4c5e281 + I66071f20991b414140869a2e3b750471;
            tout_00021_00004    = fgallag_final_00021_00004;

            I9c1a08b61782ef6c72545504693ac54e= Ic0edcf240048fbfde4e938c3e4c5e281 + Ic7ccbeaf4ab94d0660eb7a0533723e24;
            tout_00021_00005    = fgallag_final_00021_00005;

            I363594fb91d01abca7a2b7402e352fd0= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + Ib3be128b6704cc04c61e0fc9814dcf20;
            tout_00022_00000    = fgallag_final_00022_00000;

            Idd284c75a230f4b97d5acb98a8e38b2d= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + I29fb3830a5fc5922f1ec687a38941e97;
            tout_00022_00001    = fgallag_final_00022_00001;

            If040df53a6410b263f5b3dc3090631c4= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + I511a55c2f4d6d3727dff5825597f55a9;
            tout_00022_00002    = fgallag_final_00022_00002;

            I31df60ffcaea9cee63b920478cb058f1= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + I762b2abb876381eff6de97cef0798405;
            tout_00022_00003    = fgallag_final_00022_00003;

            Icdd2f6ce69b389fbf712e45bdc0a0257= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + Ib393146d81d3cf031466543311cee2ad;
            tout_00022_00004    = fgallag_final_00022_00004;

            I8971b250393b397b94db38b9fd0fe501= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + I08043393cb7f2558c145a698ea6652c9;
            tout_00022_00005    = fgallag_final_00022_00005;

            I9199e5e8fdc0e2c62ad1d62fc4d873cb= I70b1b8521b36920707e95fc9418eb8a9 + I8d4f3e64c8e3b0710a4a6b30d27c8be8;
            tout_00023_00000    = fgallag_final_00023_00000;

            I6e03f71fdf20db836c5772658a050e9c= I70b1b8521b36920707e95fc9418eb8a9 + Ie355fa27abbc41291eaf08f2cf9a6ff7;
            tout_00023_00001    = fgallag_final_00023_00001;

            I2ef49f893dbc8581725ca0f6d1c3305c= I70b1b8521b36920707e95fc9418eb8a9 + I6fb63ea54e492bdbc6d1145affc683e9;
            tout_00023_00002    = fgallag_final_00023_00002;

            I8796f168c892ac60c38a0a7f1e18035e= I70b1b8521b36920707e95fc9418eb8a9 + I1898bc3cc6a8b6f71d65c758d1f08366;
            tout_00023_00003    = fgallag_final_00023_00003;

            I64a26e5117c8f3ab95bf0dfa97427243= I70b1b8521b36920707e95fc9418eb8a9 + I2aabda12ff89e708d04b4399472b5203;
            tout_00023_00004    = fgallag_final_00023_00004;

            Id7946a0299ced3ba00f6c3e6e664931f= I70b1b8521b36920707e95fc9418eb8a9 + I84865c4f872c0845124b78fabf695c2c;
            tout_00023_00005    = fgallag_final_00023_00005;

            I5243b90640ea4680de83021601c85c39= I4fb1c32a62cbbaeb585c6564a3c938f9 + I91a8168d3b087ab3891cd6d479427b95;
            tout_00024_00000    = fgallag_final_00024_00000;

            Ic8301fceed328cc031640ecc4ff34803= I4fb1c32a62cbbaeb585c6564a3c938f9 + I2493237a24acdcab8b5bda10e804a5cf;
            tout_00024_00001    = fgallag_final_00024_00001;

            I6e852c94b6105af62ee85f8adf77fa55= I4fb1c32a62cbbaeb585c6564a3c938f9 + Ib3e7633767b6e09e4ee54f6feaddd31e;
            tout_00024_00002    = fgallag_final_00024_00002;

            I7d98c5c2a54832b6368ce60009208eb0= I4fb1c32a62cbbaeb585c6564a3c938f9 + I896cd566a3d078b0f697a788efd223f2;
            tout_00024_00003    = fgallag_final_00024_00003;

            I7e42f2281518bead81a6d18d2dcbd1a3= I4fb1c32a62cbbaeb585c6564a3c938f9 + I8c733a5d394e6b8d045eede5cc7451f6;
            tout_00024_00004    = fgallag_final_00024_00004;

            I63c126c978154f2d68b11f08a938dcb4= I4fb1c32a62cbbaeb585c6564a3c938f9 + I57b9dd7a7deea6695dcd03439c9723cf;
            tout_00024_00005    = fgallag_final_00024_00005;

            I2ff7719c35578b47720cacd9ddfd92eb= Iefc37daeec14e14ef2fe0716f73109dc + Ic970a88c435a85d21ed71c6060b8a8e4;
            tout_00025_00000    = fgallag_final_00025_00000;

            I480599aef36967a670155dd77120a37d= Iefc37daeec14e14ef2fe0716f73109dc + If83ce1cbe3a73472419520c225b288a6;
            tout_00025_00001    = fgallag_final_00025_00001;

            Ic000b2c844de484b8f30b7b84dd6234d= Iefc37daeec14e14ef2fe0716f73109dc + If86532f849bd392dbf599eeb2fae0545;
            tout_00025_00002    = fgallag_final_00025_00002;

            If0e25df151db991185f992eab5d5be99= Iefc37daeec14e14ef2fe0716f73109dc + I85a7fede715578be0634d71e9c7951cd;
            tout_00025_00003    = fgallag_final_00025_00003;

            I2f533699abb7a997160bf4ee4cda3efb= Iefc37daeec14e14ef2fe0716f73109dc + I5d4fb4b5a5ad3dc48beebfa0e0cebbed;
            tout_00025_00004    = fgallag_final_00025_00004;

            If6b33cfc6d34e33fbb18e08fb4d8a5ed= Iefc37daeec14e14ef2fe0716f73109dc + I1cd6b35bcdfd461db69a4c1bdb1d387f;
            tout_00025_00005    = fgallag_final_00025_00005;

            I2ea5423dc8726fc0217899e0f406a1e9= Ibd15f164f6d2ac9e5721a21464bc2c5c + If365a3c3ef86dca7c7315b91298c2db8;
            tout_00026_00000    = fgallag_final_00026_00000;

            Ibf3f4f8a04cbacc9624ca5cc73bf7069= Ibd15f164f6d2ac9e5721a21464bc2c5c + If2021f0735c6c5649ebac0d230fda87c;
            tout_00026_00001    = fgallag_final_00026_00001;

            I9ba53c36934ab1c7f498241a79cfbae8= Ibd15f164f6d2ac9e5721a21464bc2c5c + I12c07042202f66db926861c9ce7c2b25;
            tout_00026_00002    = fgallag_final_00026_00002;

            I106a25f18536f96782927bf3bc2ccd72= Ibd15f164f6d2ac9e5721a21464bc2c5c + Ifce70fefde8f5ea4d2c1857236f66d65;
            tout_00026_00003    = fgallag_final_00026_00003;

            Ie5cdad65e918679607cc5f816987b736= Ibd15f164f6d2ac9e5721a21464bc2c5c + Iffeefa89a2ba7d032db5db64cbf05e20;
            tout_00026_00004    = fgallag_final_00026_00004;

            Ica6dc9ded8756fd6f82eec4271e246c3= Ibd15f164f6d2ac9e5721a21464bc2c5c + I40a1ecabded8add5bffe316f2d8beda9;
            tout_00026_00005    = fgallag_final_00026_00005;

            Ica42ac6ca5813d0d1a67f14d1248437a= I951dfff9507bb70214d48e03a0ebb3a7 + I16e3f3a6802fd206654bb622fa1393fe;
            tout_00027_00000    = fgallag_final_00027_00000;

            I13dc6cfc75ef846c30e5dc1dc5305d59= I951dfff9507bb70214d48e03a0ebb3a7 + I7a029c27d92754041eb6d605837238dd;
            tout_00027_00001    = fgallag_final_00027_00001;

            I33e784182dfb4af39715788b1ae98af6= I951dfff9507bb70214d48e03a0ebb3a7 + Ib8b95ece5da3877b261a06e6d0571921;
            tout_00027_00002    = fgallag_final_00027_00002;

            I9e1a66805348d2e5bbf5e2316187444b= I951dfff9507bb70214d48e03a0ebb3a7 + I84a62a133dbceb5a32a7c907f371663d;
            tout_00027_00003    = fgallag_final_00027_00003;

            Ie9619916a96d218cf5eb5f3a4995d0e7= I951dfff9507bb70214d48e03a0ebb3a7 + I42564ec6a794ea803795f0b5b3523a93;
            tout_00027_00004    = fgallag_final_00027_00004;

            I02ce7969c51ad141df227ed7d18e74b1= I951dfff9507bb70214d48e03a0ebb3a7 + I7c52ae4af926267b5e27a530202fcce0;
            tout_00027_00005    = fgallag_final_00027_00005;

            Idd73461af0d75c4d820f7f8f0f419e0f= Ie78e30b2a2eda75d0df7d10fd67b5e36 + If79bc5a35cb55036a367efb88c7d5510;
            tout_00028_00000    = fgallag_final_00028_00000;

            I3df6c2cdccb2a82c58c1d81b00af7786= Ie78e30b2a2eda75d0df7d10fd67b5e36 + I00dad36628d2fa923120fdaa79bf0045;
            tout_00028_00001    = fgallag_final_00028_00001;

            I97f441fc5ffb88efeb5ed66b60f07a7c= Ie78e30b2a2eda75d0df7d10fd67b5e36 + Ic99654bf4833c9132912eeb4c0dc92fa;
            tout_00028_00002    = fgallag_final_00028_00002;

            I3194a235eb652c8d0e4307cd056e5e72= Ie78e30b2a2eda75d0df7d10fd67b5e36 + Ifb9b29c43f435452cc761218c509f5df;
            tout_00028_00003    = fgallag_final_00028_00003;

            Ibc315f6c79ba2bf336ee57f2e5f7d776= Ie78e30b2a2eda75d0df7d10fd67b5e36 + I514830acdad20c4ff3d078477e939b4b;
            tout_00028_00004    = fgallag_final_00028_00004;

            I937a54f5cda99a7079c7fa46b4ea26f6= Ie78e30b2a2eda75d0df7d10fd67b5e36 + I1a5c6c50817db8bde279d5f0b5095d76;
            tout_00028_00005    = fgallag_final_00028_00005;

            I49c99afecc613656cd1469d8c1e98936= Ia0b83a372dd4115dc4d61eb8ff0811b9 + I12334038c2be8634c47869f397503019;
            tout_00029_00000    = fgallag_final_00029_00000;

            Id76ce0333f43bf7bccf1ce48e25ca69c= Ia0b83a372dd4115dc4d61eb8ff0811b9 + I03829256e357ac17c7ca7cae2f980f41;
            tout_00029_00001    = fgallag_final_00029_00001;

            I2c77f9644145219005751f7a4eb71aaa= Ia0b83a372dd4115dc4d61eb8ff0811b9 + I3f193e9c265c1dfaeada63d59db5b79f;
            tout_00029_00002    = fgallag_final_00029_00002;

            I5cecc266272eef88cda88c1df9bcc37e= Ia0b83a372dd4115dc4d61eb8ff0811b9 + I9ab3cea6ee8d8473221da21bae06066b;
            tout_00029_00003    = fgallag_final_00029_00003;

            I776a0b1b5c14afa21b7fda3c2cacafed= Ia0b83a372dd4115dc4d61eb8ff0811b9 + Icf8cfc800f0a2aa5140a7f83f035b0cc;
            tout_00029_00004    = fgallag_final_00029_00004;

            I84860b1f933339e0f90beeb3d666393b= Ia0b83a372dd4115dc4d61eb8ff0811b9 + Idf0c1b85712fcbbbcc12915158ebff62;
            tout_00029_00005    = fgallag_final_00029_00005;

            Id24581713f1ecb767db39d5154c2f5f4= If5c5bcbbea01aa22f242b913f0d01929 + I715d59fb27e519a9b76bdd8b5139a619;
            tout_00030_00000    = fgallag_final_00030_00000;

            Idb0eae2f0e1dae1d56251d64e2c51f9f= If5c5bcbbea01aa22f242b913f0d01929 + Id1df78ab32daf524b77c0431c782f2bf;
            tout_00030_00001    = fgallag_final_00030_00001;

            I2e3ca4b130e6d3d92385928a28644452= If5c5bcbbea01aa22f242b913f0d01929 + Ia344734d285ac29b53cf401c08a0f987;
            tout_00030_00002    = fgallag_final_00030_00002;

            I7922d80ae333dcfafde31d294f0eb4d8= If5c5bcbbea01aa22f242b913f0d01929 + I4a0033a180d7edce81fcfef603532e28;
            tout_00030_00003    = fgallag_final_00030_00003;

            I82de04cd2dfef5616efca4af26d7c561= If5c5bcbbea01aa22f242b913f0d01929 + If0b9225e759438be175c4128c78605ea;
            tout_00030_00004    = fgallag_final_00030_00004;

            I7ce384520525b15d24c2ef6f161213a5= If5c5bcbbea01aa22f242b913f0d01929 + I6b32298e8c61e75d0a38bca3084c0528;
            tout_00030_00005    = fgallag_final_00030_00005;

            I56aeea71c7bd19d47620cf36adf3f115= Iccba58cd3519fb4cc75a61b50da1d562 + I566224393f6bb27bfd8b0b0d6b8e53d6;
            tout_00031_00000    = fgallag_final_00031_00000;

            I138e1a6db0c6649bc023cc36d81d5b47= Iccba58cd3519fb4cc75a61b50da1d562 + Ie1bf5d97b8f679095d2442bbf9f95608;
            tout_00031_00001    = fgallag_final_00031_00001;

            Ib5e8b1c4dd9b5dad56b59cc11c87a258= Iccba58cd3519fb4cc75a61b50da1d562 + I9d0fdb45b9e86bd409740e538a690320;
            tout_00031_00002    = fgallag_final_00031_00002;

            I86f785e2d5e8d6c08fad1d334c7d244e= Iccba58cd3519fb4cc75a61b50da1d562 + I4f45dd50d2825ab338b8a2a8264096c0;
            tout_00031_00003    = fgallag_final_00031_00003;

            I9a6c8efca218c724da4ee4c1087d58bc= Iccba58cd3519fb4cc75a61b50da1d562 + Ica94017f26e96fb22a47add326ee126e;
            tout_00031_00004    = fgallag_final_00031_00004;

            Ia30e8dbc6974ea94b763842e8dffa633= Iccba58cd3519fb4cc75a61b50da1d562 + I5b0d72cedc120406402076148e2d30b0;
            tout_00031_00005    = fgallag_final_00031_00005;

            Ifa60f45f4d8848eb0b89f5644ec69668= Ibc0999e4d0b3cc2650f9348b8c204b14 + I4b5713aee09999592256c407d4b8a95a;
            tout_00032_00000    = fgallag_final_00032_00000;

            I0aeb4b93cfa6d62ec41b7e6dd0287dd0= Ibc0999e4d0b3cc2650f9348b8c204b14 + I64692d5168554dfd7ce1c7a046aecf72;
            tout_00032_00001    = fgallag_final_00032_00001;

            Ifce1fc978fb5b0187593f46f53c3b469= Ibc0999e4d0b3cc2650f9348b8c204b14 + Iea71417e738c6ca54c50aa014cc38627;
            tout_00032_00002    = fgallag_final_00032_00002;

            If3b6de7c919c5d53a0e191a75bd7e574= Ibc0999e4d0b3cc2650f9348b8c204b14 + Iaf624549f73b0d13c1a73c850b99f810;
            tout_00032_00003    = fgallag_final_00032_00003;

            Iecce594e6e99b0c05fc845144a664b07= I2aeff1fb4b839a581acaf26f90f9113c + Id1dce8c1542f1279badb381aca3c9b51;
            tout_00033_00000    = fgallag_final_00033_00000;

            I2c8431500ecb25619d2884a2fb4260c0= I2aeff1fb4b839a581acaf26f90f9113c + Ibe6a876a041198a581c95457a7d1fcf8;
            tout_00033_00001    = fgallag_final_00033_00001;

            I217c710f7ef39035546efcbb043f63f3= I2aeff1fb4b839a581acaf26f90f9113c + I57db98eb439d59a895dabe029c6a3a8b;
            tout_00033_00002    = fgallag_final_00033_00002;

            I1b4236130cb1879d885653fdd9eeab4e= I2aeff1fb4b839a581acaf26f90f9113c + Iaaf7efeae9f6dc9e8222dc2b10122000;
            tout_00033_00003    = fgallag_final_00033_00003;

            Iae0f7c13f1564d63b4bfdc152ddf4111= I7d60d53f883f8187700c4e78b4c22f1c + Iec8dc328edd6cbaa2d697e05ed222746;
            tout_00034_00000    = fgallag_final_00034_00000;

            I010592496030d138a3a4245d00069957= I7d60d53f883f8187700c4e78b4c22f1c + I8fcad6e7d5ffc9f79eaaf634f6fe8cda;
            tout_00034_00001    = fgallag_final_00034_00001;

            I9d7f47a6289a16448221d61f301586aa= I7d60d53f883f8187700c4e78b4c22f1c + Ica26f542586d50c56ce0f3c00f36b388;
            tout_00034_00002    = fgallag_final_00034_00002;

            I7b8ed2953170c4deadaeb33a6ba165d4= I7d60d53f883f8187700c4e78b4c22f1c + Iea1cd2321d2ac9b891b344e2ba2363d3;
            tout_00034_00003    = fgallag_final_00034_00003;

            I4efe9eef6a48aeb0a9ba4e0ffd9906c3= Id6fcf4b7af4a37c854a12e2ae80851fa + I83560e8d0f8cd37815cca6336fb2208d;
            tout_00035_00000    = fgallag_final_00035_00000;

            I5a8466bbd83c39dfbeaa6399e3fb3337= Id6fcf4b7af4a37c854a12e2ae80851fa + Ideab06dc2448a6950cd1a06a0c90c2c6;
            tout_00035_00001    = fgallag_final_00035_00001;

            I1ab96ffa948dd09bcc4f748c6c2575d2= Id6fcf4b7af4a37c854a12e2ae80851fa + Ic5ca74b66763c6e5591c7c2bfeeb0663;
            tout_00035_00002    = fgallag_final_00035_00002;

            I016f57568eaf00b26f8a22100858c158= Id6fcf4b7af4a37c854a12e2ae80851fa + Ia544fa24b953fe91800978895e3e610e;
            tout_00035_00003    = fgallag_final_00035_00003;

            I1fb995e302f4f1ba493ff85f39938175= Ifa5e5f7d753964f14f0f16dbe552fd85 + Iec078a95a69b081cfb5e987ba9c5a613;
            tout_00036_00000    = fgallag_final_00036_00000;

            Ie643ad235307c60f1ee96dfdcbc8c2a8= Ifa5e5f7d753964f14f0f16dbe552fd85 + Ia71663e8f563041c27cd21a0c9c27a28;
            tout_00036_00001    = fgallag_final_00036_00001;

            I8dafdf2c780082d8dfc2961b3447f104= Ifa5e5f7d753964f14f0f16dbe552fd85 + Idcef10a0465614cf38e0d6f503b5174a;
            tout_00036_00002    = fgallag_final_00036_00002;

            I3a2841a0f5e1b42556f384231ab0717b= Ifa5e5f7d753964f14f0f16dbe552fd85 + If2143db72bf9a02b64eb45b3a4faa39d;
            tout_00036_00003    = fgallag_final_00036_00003;

            I2b00d0e6facf01274c0c3446bb0e1599= Ifa5e5f7d753964f14f0f16dbe552fd85 + I7fa710c37f5f96c3cdc35612a702a71c;
            tout_00036_00004    = fgallag_final_00036_00004;

            I2c645d25871b70dae5b2c283695d5130= I900d471b087cf5a436c2ad66a84d8280 + I6f0f74dcc830fdcb0af9df75a2b722f7;
            tout_00037_00000    = fgallag_final_00037_00000;

            I540a0e8968a6a82aca775a81ef82b520= I900d471b087cf5a436c2ad66a84d8280 + I0b557cf102da41afd26936cbdb64b6e8;
            tout_00037_00001    = fgallag_final_00037_00001;

            I5b95bbc82e6d8d87421efe3f17b97ea5= I900d471b087cf5a436c2ad66a84d8280 + If65eb5e743a7b1878fb232ef2fe13cb0;
            tout_00037_00002    = fgallag_final_00037_00002;

            Iad81f5e5e728ffdec6296b2aff668d75= I900d471b087cf5a436c2ad66a84d8280 + I3403ce6e697b523a9f441d8fd5e2d420;
            tout_00037_00003    = fgallag_final_00037_00003;

            I960a618f63372da74581b8c352f3e618= I900d471b087cf5a436c2ad66a84d8280 + I98fd105696fca11c1075f9bd30013747;
            tout_00037_00004    = fgallag_final_00037_00004;

            I4f5325f1601acde10018d1fd0aff4d35= I6d1434907f0292ea2ee47cbc5b52bfb9 + I1d7d7a68fc53b8be89c4637ac8f29380;
            tout_00038_00000    = fgallag_final_00038_00000;

            Ib297101fe456520e72cd9d208af44eea= I6d1434907f0292ea2ee47cbc5b52bfb9 + I3353a7916b569f2c0ca122180608dccc;
            tout_00038_00001    = fgallag_final_00038_00001;

            I73a21342321a9d81a0fa5308149d72b0= I6d1434907f0292ea2ee47cbc5b52bfb9 + Ia457938da4efe847cb06f645f2a54a52;
            tout_00038_00002    = fgallag_final_00038_00002;

            I2a486524f4f53b3454ee02a8892d4fa3= I6d1434907f0292ea2ee47cbc5b52bfb9 + Ic7a21921e2716fba55aad2e351f4498a;
            tout_00038_00003    = fgallag_final_00038_00003;

            Ic6c4e4e6a9ba43a3354f9f3192ab069e= I6d1434907f0292ea2ee47cbc5b52bfb9 + I61345963ceabdaa0f25f8a463fc9fe5d;
            tout_00038_00004    = fgallag_final_00038_00004;

            Ie3cdee3560bd06aed84dac5fcd2a259a= I938bef7ba7ae1739d8e6a6a7c117a1b1 + Ia4b438844530fff602ea04e72b07db8d;
            tout_00039_00000    = fgallag_final_00039_00000;

            I584febaa4c440fd9353108af36d3a5c6= I938bef7ba7ae1739d8e6a6a7c117a1b1 + Id4788855f9a503e8b506d012aaeea445;
            tout_00039_00001    = fgallag_final_00039_00001;

            I515e78507d7419ca14d77b6d52f75a78= I938bef7ba7ae1739d8e6a6a7c117a1b1 + I7c68e0ae30efc4ca4d68b6047119c6c3;
            tout_00039_00002    = fgallag_final_00039_00002;

            Ie9578453a57d2b3b9c3b98844044b5f0= I938bef7ba7ae1739d8e6a6a7c117a1b1 + Ib45caf6b563d22144be3e9225a99a1cd;
            tout_00039_00003    = fgallag_final_00039_00003;

            I1e58b3062097a46d8d590232b40278cf= I938bef7ba7ae1739d8e6a6a7c117a1b1 + I9e8375af6af10f4bac3e87e416d430ee;
            tout_00039_00004    = fgallag_final_00039_00004;

            I3af126eb28c67797ce625b0d82943833= I6384a9416b2d1da01df1b2d7b16c5390 + I8983f003c30a218543f39f5bbcd9a25c;
            tout_00040_00000    = fgallag_final_00040_00000;

            I130ee1a8acacf4cae8818cd8320d050d= I6384a9416b2d1da01df1b2d7b16c5390 + Ib34ad1d14978608d1440f59998a31672;
            tout_00040_00001    = fgallag_final_00040_00001;

            Idf92dd09c29ce8e921b2b34089550586= I6384a9416b2d1da01df1b2d7b16c5390 + I380ff8528cdba4026fac3c4eda8b2c52;
            tout_00040_00002    = fgallag_final_00040_00002;

            Iba74a64cc1d2ec3c83a4061db298ad37= I6384a9416b2d1da01df1b2d7b16c5390 + Ie72268e979cf069b88f6eadde789e5ab;
            tout_00040_00003    = fgallag_final_00040_00003;

            I01364c233ca541914d790354515aa5c1= I6384a9416b2d1da01df1b2d7b16c5390 + Ida1cd844022bbf1b8431225e66b2b78f;
            tout_00040_00004    = fgallag_final_00040_00004;

            Ic6a8297308a63ed3113008a3cdc76358= I5097a79e7cf7a30d38ba198d1407119c + I16d2084ccfb102c3bafc701872f5ef2d;
            tout_00041_00000    = fgallag_final_00041_00000;

            I6c7ee9d0bd684a7f54bed3d52452219d= I5097a79e7cf7a30d38ba198d1407119c + I9574759e112f27778f3645d5d49126b7;
            tout_00041_00001    = fgallag_final_00041_00001;

            I985ea87550ec8a222e6af621589e186d= I5097a79e7cf7a30d38ba198d1407119c + Ia8094903aed8dd0ce8e9ff459a5287b0;
            tout_00041_00002    = fgallag_final_00041_00002;

            I6836a7d1e006d7f7556edf8b31aea32e= I5097a79e7cf7a30d38ba198d1407119c + I502a8e382aa0881dc86f3c13e0566ca3;
            tout_00041_00003    = fgallag_final_00041_00003;

            Ia7a356a18af18ec131b9df46019f3e58= I5097a79e7cf7a30d38ba198d1407119c + I30e9ab592e97dbc5fb6ab58d2ffbf8d4;
            tout_00041_00004    = fgallag_final_00041_00004;

            If3a7e111247232c47ceccb5e05338312= Ib113c26c8dcf49c972c41a938059a787 + I099441ae3d3dffe49b18bc578af54dc7;
            tout_00042_00000    = fgallag_final_00042_00000;

            I5f38d1665294b2d3c18f9cd888ff60f1= Ib113c26c8dcf49c972c41a938059a787 + I0e8f3f56bce3be1ee4d5f780a2f2a9fe;
            tout_00042_00001    = fgallag_final_00042_00001;

            I10290b9576bf3d8caf90583a388226b7= Ib113c26c8dcf49c972c41a938059a787 + I218ee96418a4f5d734d3d71685bc09c7;
            tout_00042_00002    = fgallag_final_00042_00002;

            Ief36236305fc1521c5bb4c60753a676a= Ib113c26c8dcf49c972c41a938059a787 + Id5fd6f25dc3df22a322434ae3c90dea6;
            tout_00042_00003    = fgallag_final_00042_00003;

            Ibaa0539fbf5ccc979511c09c061cf494= Ib113c26c8dcf49c972c41a938059a787 + I2ec2a6de2be39b1bc259b0be72e35a0f;
            tout_00042_00004    = fgallag_final_00042_00004;

            I95664ffd0ff13c2893421032149f24d2= I970c4a25a8bce82a9d2846679029fcab + Ieb1dbb98d5e5bda5b9ce803857f2ca26;
            tout_00043_00000    = fgallag_final_00043_00000;

            Ie390153b3b7985dc63d65913de215377= I970c4a25a8bce82a9d2846679029fcab + Idd95fd099dd2b53c46d02f09575b8032;
            tout_00043_00001    = fgallag_final_00043_00001;

            I704147dda658f4a03627dacc1c91dd48= I970c4a25a8bce82a9d2846679029fcab + I1fc36e6f738fab96df356979e1e3a612;
            tout_00043_00002    = fgallag_final_00043_00002;

            Ifb09672d505898f081aa13c95fcb88b5= I970c4a25a8bce82a9d2846679029fcab + I2461055ef9b1aa2ffca0f5cac3300e71;
            tout_00043_00003    = fgallag_final_00043_00003;

            Ibb5cb89097dd11bf292d5b5a2422175b= I970c4a25a8bce82a9d2846679029fcab + Ic32e349efae2ca419e095ee5e15a501d;
            tout_00043_00004    = fgallag_final_00043_00004;

            I4a305956b18d6ad6901d2c17e99f2bab= Ibe2af096ad2db26e54d8b4b3bb05175c + Id1b5c33bc63f75561b7cce6fc0981c69;
            tout_00044_00000    = fgallag_final_00044_00000;

            Ibf5bb3b9eb1812383db9634fa9a27ad3= Ibe2af096ad2db26e54d8b4b3bb05175c + I2bc3ffbe5b42b0833206437d3863278e;
            tout_00044_00001    = fgallag_final_00044_00001;

            I66b37d055c3735f011095ee4b1ad02ed= Ibe2af096ad2db26e54d8b4b3bb05175c + Ice2c390d296e09b117d60905343e9098;
            tout_00044_00002    = fgallag_final_00044_00002;

            I43e71dd694d97217e242f267248cd594= Ibe2af096ad2db26e54d8b4b3bb05175c + I036342f6be0f2e2f1f4927099a5c4a78;
            tout_00044_00003    = fgallag_final_00044_00003;

            I4baa925db1ec733bd4bd25d9dc873e23= Ibe2af096ad2db26e54d8b4b3bb05175c + I1befb935ee9cb871c9a7476c1fc0da3f;
            tout_00044_00004    = fgallag_final_00044_00004;

            I547928c9db7acc531af251264d576ffb= Ie48569c467fba0c1291f71d6080ebedc + Id680a9affed622577164b3a8380494f5;
            tout_00045_00000    = fgallag_final_00045_00000;

            Ie4ce634b2fb62a20781f8a2e8fddc762= Ie48569c467fba0c1291f71d6080ebedc + I5732fdb805258fc13c8ba4aaf56574ca;
            tout_00045_00001    = fgallag_final_00045_00001;

            I0e90e96ffa64c2874d79110b622994bf= Ie48569c467fba0c1291f71d6080ebedc + Ia2fc8a1bbc3cb0dd7d89a7f05b04909c;
            tout_00045_00002    = fgallag_final_00045_00002;

            I767e37e3c6f4224eb07adeda480ce253= Ie48569c467fba0c1291f71d6080ebedc + I6bfbf7ff79ff0a6facc9ba5031239644;
            tout_00045_00003    = fgallag_final_00045_00003;

            I75fcaf2c65b7e63adac834054850c6d6= Ie48569c467fba0c1291f71d6080ebedc + I01c57f697f2af7d2c6ae904319f10725;
            tout_00045_00004    = fgallag_final_00045_00004;

            I5f1de2dfbd79204ab2db9b686d6a6862= I90e7ded06617b49cdb8b5301fe9c6a20 + I58f89947eead94b5054a0fea3520ae33;
            tout_00046_00000    = fgallag_final_00046_00000;

            I8d01de6be4091dca2589cef625c05229= I90e7ded06617b49cdb8b5301fe9c6a20 + Ic462cebbfc39190b22d20013259e39eb;
            tout_00046_00001    = fgallag_final_00046_00001;

            Ic09e773899fdd208c0fdd874933b2cec= I90e7ded06617b49cdb8b5301fe9c6a20 + I7caa41076a293edf18c7c4309fdcfc91;
            tout_00046_00002    = fgallag_final_00046_00002;

            I24a3f9fd851c4af70ef66bfcee44af65= I90e7ded06617b49cdb8b5301fe9c6a20 + I33d941ad9d4858fcfb77f0f6cf99d2ec;
            tout_00046_00003    = fgallag_final_00046_00003;

            Idd31807ecd603db8c719349a2be1be40= I90e7ded06617b49cdb8b5301fe9c6a20 + Id580f8a2748efff9b6b747c497c16e9c;
            tout_00046_00004    = fgallag_final_00046_00004;

            Iaf680cae40d1adf7649da12b31a2be0d= I4920014f5d017f4e840dc3b88526955f + Ife1c8d014675240a94f1133a78703ed5;
            tout_00047_00000    = fgallag_final_00047_00000;

            I22d948171c1a66f7a28d5e51007700ea= I4920014f5d017f4e840dc3b88526955f + Id812a8ea2a3b4a912d151be582833fcf;
            tout_00047_00001    = fgallag_final_00047_00001;

            I3954318b2392a82f2da71a0ca1504497= I4920014f5d017f4e840dc3b88526955f + I2d7715a3af03d9664729fa6df85034a2;
            tout_00047_00002    = fgallag_final_00047_00002;

            I15c78b909cbd04fe25820d777655d829= I4920014f5d017f4e840dc3b88526955f + Id32e7ad5b1aa825732d9b26d0fa02ca1;
            tout_00047_00003    = fgallag_final_00047_00003;

            Ia529c5ec88a9f6c14ceda5cad56b346d= I4920014f5d017f4e840dc3b88526955f + I77b54488bd26318f14b4364035cd1836;
            tout_00047_00004    = fgallag_final_00047_00004;

            I5b73c81f28901705f6ee26d63847db0a= I03b70553f1c501609400574ae7cd73f5 + Ia73cacadbf80c0701a5b5b430c0d5c98;
            tout_00048_00000    = fgallag_final_00048_00000;

            I1a9bd3f728db23b679639e5657ced179= I03b70553f1c501609400574ae7cd73f5 + I19eae741ef89baa1a64c403fb29f14f4;
            tout_00048_00001    = fgallag_final_00048_00001;

            I57ca72784a7c91cecbd694ddd08bcb98= I03b70553f1c501609400574ae7cd73f5 + I9d6730140c690037b5ca58aa30103f5b;
            tout_00048_00002    = fgallag_final_00048_00002;

            I50f31ecd3f2b498cc7b759efa057f12f= I03b70553f1c501609400574ae7cd73f5 + I786338397f55073dce91e1c8c5f8e298;
            tout_00048_00003    = fgallag_final_00048_00003;

            I8ccaf29848defdd264f522642968fa29= I63c9bf68b43ed66c51b0f4c0ed92e9ab + I0f277bc88d46a4e6e9f1f2c410b503fd;
            tout_00049_00000    = fgallag_final_00049_00000;

            I808ea92ee1340876cf1d2c47255dc2fe= I63c9bf68b43ed66c51b0f4c0ed92e9ab + Id9d56f09595e80d66c2ac300f7d1d972;
            tout_00049_00001    = fgallag_final_00049_00001;

            I3da806790125328b626be1949f71267a= I63c9bf68b43ed66c51b0f4c0ed92e9ab + Ice780b1695a8e80607a03dee3c426ffe;
            tout_00049_00002    = fgallag_final_00049_00002;

            I55e59bc1daeb8b2be3d7a1e4b272df93= I63c9bf68b43ed66c51b0f4c0ed92e9ab + I0e5931219d94c8e8e1f4af081404dcab;
            tout_00049_00003    = fgallag_final_00049_00003;

            Ib0ffadc6a0091ceff91ad1fa435413a6= If408dfead07757878cc878131bc7d6a3 + Id081512cd113e4d09df0fb13e443d76b;
            tout_00050_00000    = fgallag_final_00050_00000;

            Ic863f139e6bed2d06789a07c6dedf6f8= If408dfead07757878cc878131bc7d6a3 + I38cc7b117c0bcd5e3060cd370d710d7e;
            tout_00050_00001    = fgallag_final_00050_00001;

            Id0e8f6ada5060a911090f76cfaa3c6bf= If408dfead07757878cc878131bc7d6a3 + Ia98a70144e466b356d2998948dc4b602;
            tout_00050_00002    = fgallag_final_00050_00002;

            Ibb8c9b8fc9b58f5f8a6ad342934804a8= If408dfead07757878cc878131bc7d6a3 + I8d96b419b010f8076311420d7b9c8a18;
            tout_00050_00003    = fgallag_final_00050_00003;

            I9323a188737ca54c2dd553cd99bd416c= Ia0857d63d309807789b6ff4f6028f1b3 + I2ffb7c2ad09bac694ef13ec41e5de327;
            tout_00051_00000    = fgallag_final_00051_00000;

            I2694cef38855f496e7ca12f42dfdb9fc= Ia0857d63d309807789b6ff4f6028f1b3 + I81800fb49855a4fd2737faa07ff15d29;
            tout_00051_00001    = fgallag_final_00051_00001;

            I75790b4c0b1f6c7935f5cfbea26407d1= Ia0857d63d309807789b6ff4f6028f1b3 + I9a3f0b4867087790c78f674b719dbf7b;
            tout_00051_00002    = fgallag_final_00051_00002;

            Ib8b366c47e56a49fc53ea4a9e1ebbd99= Ia0857d63d309807789b6ff4f6028f1b3 + Ife13f962c7a8df3845cde104a959f678;
            tout_00051_00003    = fgallag_final_00051_00003;

            Ie1c86256df2bc6c4dad41237eca41986= I53921b825c5e434b63bee0e1ecb7a517 + I003f95fb8f2027efa41a1936e8b53986;
            tout_00052_00000    = fgallag_final_00052_00000;

            I7c9e3f97a94f9a078c209a1b84ff916d= I53921b825c5e434b63bee0e1ecb7a517 + Ib190f589f4d663dbc0a3c166a8dcf5fa;
            tout_00052_00001    = fgallag_final_00052_00001;

            Idde839d34403fdbba62671b83801ea8d= I53921b825c5e434b63bee0e1ecb7a517 + I49eb064043f91112c854e31e4eb9b885;
            tout_00052_00002    = fgallag_final_00052_00002;

            I824e23c3e43434e0a7bf8c8b8e0de597= I53921b825c5e434b63bee0e1ecb7a517 + Ia0868eee7e7e0640ce1a4d3ca9c001cb;
            tout_00052_00003    = fgallag_final_00052_00003;

            I0f83a2c488c229e971030fc66ce212f5= I53921b825c5e434b63bee0e1ecb7a517 + I7f701ff37ad3fc34d2f4efafe5ff5351;
            tout_00052_00004    = fgallag_final_00052_00004;

            I8fdda3dea7a63fd6e57f70365d7b6571= I5e68f84e123c37f19a03c13892c77e19 + Ifcd68be4bea38622d2d57d3a4e6fc5bb;
            tout_00053_00000    = fgallag_final_00053_00000;

            Ifa2fc30c14c549339edc65c3670d90a0= I5e68f84e123c37f19a03c13892c77e19 + Ic634d26fc09589a29a160e4efb5613a8;
            tout_00053_00001    = fgallag_final_00053_00001;

            If69bb1bfa10ca7dd37ba57485c3429e7= I5e68f84e123c37f19a03c13892c77e19 + Ibfe760474fcac99f1e5ffa2e008fef99;
            tout_00053_00002    = fgallag_final_00053_00002;

            I2ab0738fa2d5916d77a81b9da2315376= I5e68f84e123c37f19a03c13892c77e19 + I51b5e641856239367cf43f9b5679b268;
            tout_00053_00003    = fgallag_final_00053_00003;

            I50a9ce776ad2ccd8048b56ce101c80d2= I5e68f84e123c37f19a03c13892c77e19 + I43c815a8ce0b2df9744a525328969691;
            tout_00053_00004    = fgallag_final_00053_00004;

            I9c9d0332ee7ad6a3488b7e39bcb06ca2= Id5270b57c6fb4b18db3bbd0a523e467e + Ibf565bf1803ed43120fa54b80f6f1f29;
            tout_00054_00000    = fgallag_final_00054_00000;

            Idc155814976f0aef9b56b2bb3d52b3a5= Id5270b57c6fb4b18db3bbd0a523e467e + I66b92f1de2cf408c3af53b161a6ffa60;
            tout_00054_00001    = fgallag_final_00054_00001;

            I2e02fbd496d08acb3ad3359b49b9f680= Id5270b57c6fb4b18db3bbd0a523e467e + I5b937934e7aae1f916c2848889f12685;
            tout_00054_00002    = fgallag_final_00054_00002;

            If0f8b3dfce99a5a75c2105d45ccad985= Id5270b57c6fb4b18db3bbd0a523e467e + Iedb655aa25e5f0e35137ec6c3acdc527;
            tout_00054_00003    = fgallag_final_00054_00003;

            I6790223e6a7cf136a7e2b261ba4fdb0a= Id5270b57c6fb4b18db3bbd0a523e467e + I6c4a1ded9bf39091cf302ebe0103e2f0;
            tout_00054_00004    = fgallag_final_00054_00004;

            I6a9643afea7a6cc9b94806ccc8e84c0f= I3c18a84617eb21472d53e598700d7f4c + I94d9412a7b43fa0bd4b9a6d32d313fc7;
            tout_00055_00000    = fgallag_final_00055_00000;

            Id3d19d7c2b941930478a7ab01049e390= I3c18a84617eb21472d53e598700d7f4c + I57a0f8c3710cf8e216d6dc2420f7621c;
            tout_00055_00001    = fgallag_final_00055_00001;

            Ib0a25312d51cb6aa1741f7e425bc5cd8= I3c18a84617eb21472d53e598700d7f4c + Ib46b13498ec14ceaa56719f26f18febb;
            tout_00055_00002    = fgallag_final_00055_00002;

            I44dd1b66f5a9a6b0b976d3d61d6c5cbe= I3c18a84617eb21472d53e598700d7f4c + I78ade92efd265027807c861be44a10af;
            tout_00055_00003    = fgallag_final_00055_00003;

            I3ee456f2f0e7f447ae92b7523136adb5= I3c18a84617eb21472d53e598700d7f4c + Icd4ff8d14af2699db2b5168027894ebb;
            tout_00055_00004    = fgallag_final_00055_00004;

            Ic110e2a08b550acd3c8bda4a1bc2bbae= Id36663e7a01fff3170833ecfecac1321 + Ie1374cac341cf353b1863dae9f544e8b;
            tout_00056_00000    = fgallag_final_00056_00000;

            I3f87162d2874effd66a82f821aa6c73a= Id36663e7a01fff3170833ecfecac1321 + Ie018f3003c5f124bddd13c359257bf35;
            tout_00056_00001    = fgallag_final_00056_00001;

            I660ea6d341fcb38f108270c08d82473b= Id36663e7a01fff3170833ecfecac1321 + I90b0296f5ef87dfaa6110fc2e9d6ed9d;
            tout_00056_00002    = fgallag_final_00056_00002;

            Ic128d603fc08affd2f3d0ab3425710e5= Id36663e7a01fff3170833ecfecac1321 + I0c59e8c82a31aacbf5977ff778a7ff49;
            tout_00056_00003    = fgallag_final_00056_00003;

            Id5372641727970383a59e08f550814b4= Id36663e7a01fff3170833ecfecac1321 + Ia79d52fe2130426c07890fcaa50137db;
            tout_00056_00004    = fgallag_final_00056_00004;

            Ie99ad992d66880542dcd330ef6ccee04= I8d3be15109c7007a79fecaac0d891626 + Id28d9545e8d20ac080fbac5e345692da;
            tout_00057_00000    = fgallag_final_00057_00000;

            I9ed0b194f7d210d57c54b289e01c75e6= I8d3be15109c7007a79fecaac0d891626 + I924514226fdb5bac110a2650bcb2e85f;
            tout_00057_00001    = fgallag_final_00057_00001;

            I227828831c4ad21b06ed00fb5781b0e3= I8d3be15109c7007a79fecaac0d891626 + Ie4ca0836695d951ee09622892ee35928;
            tout_00057_00002    = fgallag_final_00057_00002;

            I09d5ad12cb836adfbb4833ee80fad2c9= I8d3be15109c7007a79fecaac0d891626 + I2bc5a10c587d89d10021aa5eaafb490a;
            tout_00057_00003    = fgallag_final_00057_00003;

            Ifa9c94ee94e4beb2e7c8d2d57150df41= I8d3be15109c7007a79fecaac0d891626 + I308aaa8ac500b5589aa4af533a9062bf;
            tout_00057_00004    = fgallag_final_00057_00004;

            Icb88e59e194db215382e8e949603a9be= I92169cc57291f20d336a479e392ec271 + Iaa164a078c8cdaad694a053c9c1e0313;
            tout_00058_00000    = fgallag_final_00058_00000;

            Id4ebd28aaf1076acec266666f88a02ad= I92169cc57291f20d336a479e392ec271 + Ie2d8c84d8c9a4c8f637068a2ae39fdde;
            tout_00058_00001    = fgallag_final_00058_00001;

            Idf0a0bd862167392357501b3233a8d8c= I92169cc57291f20d336a479e392ec271 + I138f008a6206a1067bb0e22ce3d90990;
            tout_00058_00002    = fgallag_final_00058_00002;

            If94cdb867ea0fc2c5578b16aacb1acfc= I92169cc57291f20d336a479e392ec271 + Icb3ab2c67a87b2ee158e0021b72fc186;
            tout_00058_00003    = fgallag_final_00058_00003;

            Ib8c066b0700941a4fa739820ff12b948= I92169cc57291f20d336a479e392ec271 + Iac91f4037e542d9fda30fadafe7e79ac;
            tout_00058_00004    = fgallag_final_00058_00004;

            I11e0f8dc46b286bafb05f901f968e1ad= I6178b220b469b40dac39168057023a1c + I459c59ac61179d74170db53bf45ba89e;
            tout_00059_00000    = fgallag_final_00059_00000;

            I608537f5639d5e0cd3e80453e21f6f85= I6178b220b469b40dac39168057023a1c + Iee8f9b0654f6f6797f11cae0947e454e;
            tout_00059_00001    = fgallag_final_00059_00001;

            I0e9d8db1bb6347c9507b645132308b3a= I6178b220b469b40dac39168057023a1c + I9df5b63f66c162d517daa69f5d0e6095;
            tout_00059_00002    = fgallag_final_00059_00002;

            I17033b417fa383a2db41d157df33d9de= I6178b220b469b40dac39168057023a1c + I2d1a5645b126761fc7fb70d24e37189a;
            tout_00059_00003    = fgallag_final_00059_00003;

            Ib7f45dbcad513b4dafee60f33622b0c3= I6178b220b469b40dac39168057023a1c + I8cd5970682bc84881489c12ff073212c;
            tout_00059_00004    = fgallag_final_00059_00004;

            Ibfbd8e00e00272f32428c7b4a3c53050= I55342938216a0ea0889f96c2f6c05ce5 + Ie16dc913f571ae73ce03d755077345a9;
            tout_00060_00000    = fgallag_final_00060_00000;

            I27973d1d4e07eaa49608d6f6975d0a93= I55342938216a0ea0889f96c2f6c05ce5 + I7e0474089ebc1c34747be1bc17a81d72;
            tout_00060_00001    = fgallag_final_00060_00001;

            If77fcedbcf99f89045de87e5cae45d8a= I55342938216a0ea0889f96c2f6c05ce5 + I48ad9b737892d7c49340ed679f46e034;
            tout_00060_00002    = fgallag_final_00060_00002;

            Ie8f8691820e7a560db8116f38dae5d49= I55342938216a0ea0889f96c2f6c05ce5 + I1ee27be7e1a38aff0039b21c45f406d1;
            tout_00060_00003    = fgallag_final_00060_00003;

            If0b19af59ad851aded19970494514034= Idf28431c76a84a48dd895979d2b11a63 + I16deb9107193a3536979e4b5e5654b9c;
            tout_00061_00000    = fgallag_final_00061_00000;

            I98b8e05818925a4b65082fa57affde83= Idf28431c76a84a48dd895979d2b11a63 + Iccca1936f4c1c9496205e77b588e9985;
            tout_00061_00001    = fgallag_final_00061_00001;

            I69317e8c556ed67630829c990f8b74db= Idf28431c76a84a48dd895979d2b11a63 + I1b40adfd6fa6c943dfa8d230d9e65514;
            tout_00061_00002    = fgallag_final_00061_00002;

            I9147d103cf235310393f9339f1cbb376= Idf28431c76a84a48dd895979d2b11a63 + Idf90f01353ad1057e11fd060442f4e53;
            tout_00061_00003    = fgallag_final_00061_00003;

            Ibe0b2cab6e2d3f3cc8baf3623ff50988= I1ef61124c8d62e8f6a82a729fb091694 + I619957528c630e7f64924a25127c93fb;
            tout_00062_00000    = fgallag_final_00062_00000;

            Idc64f1443dd2497dfaa223cda3fbd682= I1ef61124c8d62e8f6a82a729fb091694 + Ibd4aaf02982068ffbfd1b8b3795d9217;
            tout_00062_00001    = fgallag_final_00062_00001;

            I6e37e92b812099985436851da8a6ccb2= I1ef61124c8d62e8f6a82a729fb091694 + Icd37da8ea84a606529e32b2db4eb7f5f;
            tout_00062_00002    = fgallag_final_00062_00002;

            I057df2bf67d5580275654bdc28b40027= I1ef61124c8d62e8f6a82a729fb091694 + Id45f4e0f142b6c3925f24a37dcf7c0ae;
            tout_00062_00003    = fgallag_final_00062_00003;

            Ie87a151c8b90942a899b8167bcb34afb= Ib8bb96f0372323e6a8072ca56fb9396d + If13e359e530823319046ce20027445dd;
            tout_00063_00000    = fgallag_final_00063_00000;

            I735752035af159b48f53d8302bb33c21= Ib8bb96f0372323e6a8072ca56fb9396d + I24ae7de3549a84f4f88f561b6017b7a8;
            tout_00063_00001    = fgallag_final_00063_00001;

            I1f26bc7cb30a9659a638e2ab65e1f187= Ib8bb96f0372323e6a8072ca56fb9396d + I485a48b4ff4da08f977425fd10e6d392;
            tout_00063_00002    = fgallag_final_00063_00002;

            If39a50e88c4a7c43428c1d15b0bfbbcc= Ib8bb96f0372323e6a8072ca56fb9396d + I52a9bcfbd2d3a763671f19cfeaf7bb8b;
            tout_00063_00003    = fgallag_final_00063_00003;

            Ibf966c12f049d603361ad32f55b0a2c8= I432f74dda4f6b1cebdf5ad59c659080b + Ia07447985347e9a7f3739bd98867cdfb;
            tout_00064_00000    = fgallag_final_00064_00000;

            Ie1b3ed6d3fdae47669d3c4cb8af8d969= I432f74dda4f6b1cebdf5ad59c659080b + I4b94402a53d981e953c21ef316c709b7;
            tout_00064_00001    = fgallag_final_00064_00001;

            I4ec6c8d9e87224ecbe7c69d92f9419c8= I432f74dda4f6b1cebdf5ad59c659080b + Ie8c79e6a5378808c0ead5a4b24319ce9;
            tout_00064_00002    = fgallag_final_00064_00002;

            I2acb34de8c3fc53117a7ea4f9ce7dd2b= I432f74dda4f6b1cebdf5ad59c659080b + Ic8df04756f67e6dd29f3374c5f86d451;
            tout_00064_00003    = fgallag_final_00064_00003;

            I7fa4009267e80ea7eb71194843c3b22b= I432f74dda4f6b1cebdf5ad59c659080b + Ia3cc6acf2cae41e560e09993007ffd2b;
            tout_00064_00004    = fgallag_final_00064_00004;

            I6854329daadea2734e52180a41f56bcc= Idc689442305acd00f0f32416d8fb3773 + I4a5cfd6ebd47cda4fa2e06ba9ad6e5b2;
            tout_00065_00000    = fgallag_final_00065_00000;

            Ifca16aebaf75b2990188de201e4536fd= Idc689442305acd00f0f32416d8fb3773 + I2a3eb42a4402e873d081f94a14a99c20;
            tout_00065_00001    = fgallag_final_00065_00001;

            I46cc26afc8475f2fb290eefc95a542eb= Idc689442305acd00f0f32416d8fb3773 + I04a9c9765fd468a7e841577f09fc287b;
            tout_00065_00002    = fgallag_final_00065_00002;

            Id746d6515cec9e60e7478898a09787e5= Idc689442305acd00f0f32416d8fb3773 + I9937af6fcf9d834f308bc3683d524981;
            tout_00065_00003    = fgallag_final_00065_00003;

            I09a3ad636db96e00adac78c3c94bdaaa= Idc689442305acd00f0f32416d8fb3773 + Iba0d2f08788f2208a648ae7b5414195d;
            tout_00065_00004    = fgallag_final_00065_00004;

            I28b3baa225a5fd602c9fee9c948ae58b= Ida03738adc101c03c2229756bed2469d + I7eb76b3d17296fdae702d8f820f1428d;
            tout_00066_00000    = fgallag_final_00066_00000;

            Ibe12ef0f56d875c7a44030882deb0e29= Ida03738adc101c03c2229756bed2469d + I928a0e4951208aab170656596f456209;
            tout_00066_00001    = fgallag_final_00066_00001;

            I9bd9979e4acc4944227a4bd62b910c1d= Ida03738adc101c03c2229756bed2469d + I0eb3df4d4094e09e6c4b3c788baed61f;
            tout_00066_00002    = fgallag_final_00066_00002;

            Idcfa802f458499150055dbe4b1ce8146= Ida03738adc101c03c2229756bed2469d + I7c6862830daffc98cb2c1fc121d82c38;
            tout_00066_00003    = fgallag_final_00066_00003;

            Iee010958cc3e9389cb8ecacff84fccee= Ida03738adc101c03c2229756bed2469d + I9f7df6ad60284c812aeb522974578e0b;
            tout_00066_00004    = fgallag_final_00066_00004;

            I3d74b31096917c53757c829a67cf06df= I4d14c75f28f3e516c259ea288996131b + Ie5e432a991aff25577639f1b4ffd594f;
            tout_00067_00000    = fgallag_final_00067_00000;

            Ic27031a9654db9459815fe0ca35408db= I4d14c75f28f3e516c259ea288996131b + I571ddcb0a10938e4c0816c965214b4a8;
            tout_00067_00001    = fgallag_final_00067_00001;

            Idf6ead2c37f75f3cde1d4b40cd73db00= I4d14c75f28f3e516c259ea288996131b + Ie626a24e3680f7d3995dd0c2ce60cbcc;
            tout_00067_00002    = fgallag_final_00067_00002;

            I66a56161cd0ed67f65834b9eb0e94d17= I4d14c75f28f3e516c259ea288996131b + I5ab556386d2973354a5551ba9823e4ba;
            tout_00067_00003    = fgallag_final_00067_00003;

            If6de990e26ca9e8efc009188f8a5a4d9= I4d14c75f28f3e516c259ea288996131b + Iab1fb7006598181bd8749ed90c519b13;
            tout_00067_00004    = fgallag_final_00067_00004;

            I8d866786bb2dea06f5b30f6ea80cff17= I6e6cbbf430d57f347a0d70558af143d8 + I72064a6a84ff956d76a5aa590bbc05a9;
            tout_00068_00000    = fgallag_final_00068_00000;

            I01ca9a1d4901ec9b2a64300617ce4cd1= I6e6cbbf430d57f347a0d70558af143d8 + Iae32c44b88fe7ddb5d4f19cf8fff3ba6;
            tout_00068_00001    = fgallag_final_00068_00001;

            I2dbead35e15afb9affaa6ad4edd3829e= I6e6cbbf430d57f347a0d70558af143d8 + Id6f7923a16cc5adc96a730083153ca6d;
            tout_00068_00002    = fgallag_final_00068_00002;

            I83c57653e24cc09214075b04b06bad83= I6e6cbbf430d57f347a0d70558af143d8 + Icf19dd665616a8c96146b3ab9f46c741;
            tout_00068_00003    = fgallag_final_00068_00003;

            I56b9c1f555b24c2dc197168decfdb8d1= I6e6cbbf430d57f347a0d70558af143d8 + Ieef3b299ec35075c71ef9fb10525bfc4;
            tout_00068_00004    = fgallag_final_00068_00004;

            Id5c48111f1b93de2cfe89f92fd182b43= Ib7487df45118e44acec6b9d07bbd5969 + I2121318f589878b4a9260625f97de518;
            tout_00069_00000    = fgallag_final_00069_00000;

            I32908c3c90ed6488357ce4869e8a1721= Ib7487df45118e44acec6b9d07bbd5969 + Iff142b88493149045fc0de355b767c16;
            tout_00069_00001    = fgallag_final_00069_00001;

            I16b4601f2e07e6cecdb5a030178e75c0= Ib7487df45118e44acec6b9d07bbd5969 + Iebee55168fb47664095b11c9f6641124;
            tout_00069_00002    = fgallag_final_00069_00002;

            I0ae08a41ebd0e6b402a4980478087bb5= Ib7487df45118e44acec6b9d07bbd5969 + I64f65df774d29696425ba460dda09b68;
            tout_00069_00003    = fgallag_final_00069_00003;

            Icb57267a66f117943e964dd6420d7a58= Ib7487df45118e44acec6b9d07bbd5969 + I58a7c08adf48d0737c5803e2a818c045;
            tout_00069_00004    = fgallag_final_00069_00004;

            Icfa47fb87b74106cd3814adfce909424= I492f382fea500462b3d0866240fb91b2 + I62bda8dc70e0b5eb38abe094bbe92fc6;
            tout_00070_00000    = fgallag_final_00070_00000;

            I63067cef0e1a348a3e6d8cd9bd88b907= I492f382fea500462b3d0866240fb91b2 + I632469889d6bb1c268b45fb805467ebd;
            tout_00070_00001    = fgallag_final_00070_00001;

            I10aa5ba0f53632578c0e1cefa4bf4fde= I492f382fea500462b3d0866240fb91b2 + I9ca81c841a75a9ac242835956509e0fe;
            tout_00070_00002    = fgallag_final_00070_00002;

            I427c0215d0ac047e8402c20610676752= I492f382fea500462b3d0866240fb91b2 + I546122346a22ad64a6ab2b4978cde095;
            tout_00070_00003    = fgallag_final_00070_00003;

            Icf4efa87688bd1b80437686eb0126057= I492f382fea500462b3d0866240fb91b2 + I30a1c8fcd9a510a6ed559f07dd809b90;
            tout_00070_00004    = fgallag_final_00070_00004;

            Ic373f785ddd1bf8eccce263df5a82c87= I3fb3ebddaf28efb56092d19a1b4695de + I00ecb5e329390023b318a2ceba0df231;
            tout_00071_00000    = fgallag_final_00071_00000;

            I56f8e8d2d7052af26528530d389b6dc1= I3fb3ebddaf28efb56092d19a1b4695de + I3707f68de059df0af5c652fc0478e543;
            tout_00071_00001    = fgallag_final_00071_00001;

            Ifb145bc18d435fb66779e7415417bc0f= I3fb3ebddaf28efb56092d19a1b4695de + I7b929c228c865112f00bc6b4dcc95b52;
            tout_00071_00002    = fgallag_final_00071_00002;

            I62a6e0c9952d6c6e6095e2364df93078= I3fb3ebddaf28efb56092d19a1b4695de + I463f4f370e1ecad71de44780eff10df4;
            tout_00071_00003    = fgallag_final_00071_00003;

            Id6405c2b2b9aea6bc457f1064d5f3ffa= I3fb3ebddaf28efb56092d19a1b4695de + Ic4f5e9d49419e1c57cfa387761ab643d;
            tout_00071_00004    = fgallag_final_00071_00004;

            I079df9611bd81f672f2ae028bf267995= I22a26b7f0b1c8c16b00597732ce2ab23 + I28cac65a4db3f708cc90a1b023bfe894;
            tout_00072_00000    = fgallag_final_00072_00000;

            I096b226cc511363946a39307a7d97867= I22a26b7f0b1c8c16b00597732ce2ab23 + Idc57f37015a48393608e2b026bc7065c;
            tout_00072_00001    = fgallag_final_00072_00001;

            I4cc42c5a75ef339510ee0e86fb44e16a= I22a26b7f0b1c8c16b00597732ce2ab23 + I385d03def4cfb49f54867687ebd710ed;
            tout_00072_00002    = fgallag_final_00072_00002;

            I680c01c3327cb9372a42c1ec5b4193e3= I22a26b7f0b1c8c16b00597732ce2ab23 + Id3dd71ea0bf0f2996fbe42b8c3318762;
            tout_00072_00003    = fgallag_final_00072_00003;

            I83451a072082194ecb3f9419edd728b3= I2ac08a2d8c917ecb37fbaf5325cb0473 + If3cc31fd16469339470702045fc6d0da;
            tout_00073_00000    = fgallag_final_00073_00000;

            I52ad85b6a1c822ca8c2459bde8fbd510= I2ac08a2d8c917ecb37fbaf5325cb0473 + I114c595caa67a3f777f087a634130a6d;
            tout_00073_00001    = fgallag_final_00073_00001;

            I1c44d2ef638825862061a8ee1a0a2f95= I2ac08a2d8c917ecb37fbaf5325cb0473 + Ifd3638d44e1ba2285891fac152dee327;
            tout_00073_00002    = fgallag_final_00073_00002;

            I8fa1fd425809cc39cd8e2785773c1d7a= I2ac08a2d8c917ecb37fbaf5325cb0473 + Ib834b91bf81067e8efa9d470023e8b9d;
            tout_00073_00003    = fgallag_final_00073_00003;

            Ifa22335f04d35680eb8cfec8f862f357= I50ff8f51e75fb9ce3db983c2a0f57196 + I221777352b48c4e228c6637410113854;
            tout_00074_00000    = fgallag_final_00074_00000;

            I6aff673c27811b81530453906312aa9c= I50ff8f51e75fb9ce3db983c2a0f57196 + Ie3e54a4700d8d0f6478187e06cb6f85d;
            tout_00074_00001    = fgallag_final_00074_00001;

            If674ac0540f457a21235664c213d4923= I50ff8f51e75fb9ce3db983c2a0f57196 + Id5e02d4c48fa6c3b0d45a9e66f09448f;
            tout_00074_00002    = fgallag_final_00074_00002;

            Iac223ac498bdcf2cb2514582aeaf76f3= I50ff8f51e75fb9ce3db983c2a0f57196 + Ic6ead78ed741442f17a15a157cd6ef9c;
            tout_00074_00003    = fgallag_final_00074_00003;

            I7f40931ab78ededfcb52ccaac9b81282= I444bc340ffb7ef7b72d4d2e761d58872 + I86e53eed5b857c439039238bb486067c;
            tout_00075_00000    = fgallag_final_00075_00000;

            Iab7c8dad0ca20eb0988fbd99f25591a8= I444bc340ffb7ef7b72d4d2e761d58872 + Ice18bceb10fec484ffc96155e14c4974;
            tout_00075_00001    = fgallag_final_00075_00001;

            I3cb5f890a5bd3daaae34c8dfb6ecfc49= I444bc340ffb7ef7b72d4d2e761d58872 + I3afe987d8f2c93cc19534a3221d1939c;
            tout_00075_00002    = fgallag_final_00075_00002;

            Id80e145586d7e539a6514dd67ebabf6a= I444bc340ffb7ef7b72d4d2e761d58872 + I4e257dbd6f196a02dc0f5a2e5f6047d7;
            tout_00075_00003    = fgallag_final_00075_00003;

            I01e09bc554768f30dc490041d19b4da2= I039c6cac5830759529595a958b7f65c9 + I89433799cfa534afd66e8d6b9f1b62b9;
            tout_00076_00000    = fgallag_final_00076_00000;

            I0196f7df6f834ae20c4fdd127e66104d= I039c6cac5830759529595a958b7f65c9 + I223b05d94c09b095d1988df121aa5e37;
            tout_00076_00001    = fgallag_final_00076_00001;

            I4669c4f256c123a0fcceb55c1e72193a= I039c6cac5830759529595a958b7f65c9 + I788c64785b992c675fe348a1fa181525;
            tout_00076_00002    = fgallag_final_00076_00002;

            I4a02ffa2a79df824f406909aa189a404= I039c6cac5830759529595a958b7f65c9 + I3dbfbd34d1fdfd4f422d900154123b6b;
            tout_00076_00003    = fgallag_final_00076_00003;

            I3117e5029119e70846dff61d746699e7= I0584de7d919236ab138e288a27d08ff1 + Ie763738b7faf253837e1c45de255cb5e;
            tout_00077_00000    = fgallag_final_00077_00000;

            I1e4e705b3bda1451fc384cd934c0bb52= I0584de7d919236ab138e288a27d08ff1 + Iea32ebc385c6cfc9212ff37973a0a05d;
            tout_00077_00001    = fgallag_final_00077_00001;

            Ib5bea8e0072de3de2c8431ea6a35dd51= I0584de7d919236ab138e288a27d08ff1 + I449c77140475475b138d839a74078337;
            tout_00077_00002    = fgallag_final_00077_00002;

            I7d9d94022ea95ea01cddc237f3df8cb8= I0584de7d919236ab138e288a27d08ff1 + I529b763dace1924613d184c6c70c2708;
            tout_00077_00003    = fgallag_final_00077_00003;

            I3f0f9aab07427fa81fc3096c6b6d3d6d= I086402c82ec67ae09a9e6360c58904b4 + I338ccc17dc6158aec0129c8b0c02c429;
            tout_00078_00000    = fgallag_final_00078_00000;

            I12a7983041f9c298d533bad58f41d24b= I086402c82ec67ae09a9e6360c58904b4 + Iea74ecbac92e1b8f2ec7ad68d10b8e7d;
            tout_00078_00001    = fgallag_final_00078_00001;

            I78503880e5c96ec0a03c75266b1226e8= I086402c82ec67ae09a9e6360c58904b4 + Ib0b46b99e61d724ae664d9d1fec1e29f;
            tout_00078_00002    = fgallag_final_00078_00002;

            I8adeae445b33f634977957bb1a2259aa= I086402c82ec67ae09a9e6360c58904b4 + I7a600aeb6cf8c3311c10afa4d82767a1;
            tout_00078_00003    = fgallag_final_00078_00003;

            I73bd13f381d15e0b0198b60cee44bb42= I1cefdc831c146187c77f861b3e2d1af0 + I1ee46fec2b82cf8e5142f8e2ac5d9d8a;
            tout_00079_00000    = fgallag_final_00079_00000;

            Ic8b651c2b043a4a6e4cd259774322230= I1cefdc831c146187c77f861b3e2d1af0 + Ibd8424c228f87f85df3da6204edff2b5;
            tout_00079_00001    = fgallag_final_00079_00001;

            I76979d7df582f9306e796a03cb540963= I1cefdc831c146187c77f861b3e2d1af0 + I59d4567d3355fdae5660a1364d1b8d00;
            tout_00079_00002    = fgallag_final_00079_00002;

            If61d4585986757a525c54589ec93d8c6= I1cefdc831c146187c77f861b3e2d1af0 + I8c7aab31f8cb705ea13a41a5bd349303;
            tout_00079_00003    = fgallag_final_00079_00003;

            I1bc5766a4a3cc2b468ab8ef62eab691c= Ida9c16ae57d17b6faee8a54838860447 + I4f72d0db9fcc358c6fbec9964fbe0bbb;
            tout_00080_00000    = fgallag_final_00080_00000;

            I21585169e5fceda643bd03fddf8153be= Ida9c16ae57d17b6faee8a54838860447 + If6d436031f68ef587750c5c1dfcfffc2;
            tout_00080_00001    = fgallag_final_00080_00001;

            Idb2990946f60939136b3bfddbc7b1671= Ida9c16ae57d17b6faee8a54838860447 + I2b54a135e59945901e9c11580a29ee3d;
            tout_00080_00002    = fgallag_final_00080_00002;

            Icfbf703890f684bfc96decc429deaa04= Ida9c16ae57d17b6faee8a54838860447 + I171149dcaab2c0f0e2a10547ad95084d;
            tout_00080_00003    = fgallag_final_00080_00003;

            Id5bb42639a1c1c1d67df1c89a14a2bfc= Ia3b9fb112f39dd0ccbf7555659369efb + I8a7fb51566bf215af214cd2fb5209974;
            tout_00081_00000    = fgallag_final_00081_00000;

            I55b8ef91d667c1c1d9e58dbc86a2288a= Ia3b9fb112f39dd0ccbf7555659369efb + I97a75b8625ae2a143cf364790ae77753;
            tout_00081_00001    = fgallag_final_00081_00001;

            I17ff683da41b469c8c8b82ee32a7378a= Ia3b9fb112f39dd0ccbf7555659369efb + Idf8ebc0d747ae143aa61866e33d458c0;
            tout_00081_00002    = fgallag_final_00081_00002;

            I51f10296c38872338ec7df35ccd520d8= Ia3b9fb112f39dd0ccbf7555659369efb + I23b60ca4da2df0ec40c1df62d058deef;
            tout_00081_00003    = fgallag_final_00081_00003;

            Ia59ff33765ddf4aeb17f90a70c01d76c= Ib1bfcdc0c972aafc99116ed8c0511445 + I5f73e5faf1aca83ee0a415c9ac4a1b9a;
            tout_00082_00000    = fgallag_final_00082_00000;

            Ibf97abffb1ec40f2f0e099a814e04ab2= Ib1bfcdc0c972aafc99116ed8c0511445 + Ice6db5ba70d3c7499df6723a2df56bfe;
            tout_00082_00001    = fgallag_final_00082_00001;

            I3efc3271e18a1e350473dcf3375088aa= Ib1bfcdc0c972aafc99116ed8c0511445 + Ic0954671eb1dc893c3932e456800fadf;
            tout_00082_00002    = fgallag_final_00082_00002;

            I1efd1220ea9100f2fb4f169ceaf462a5= Ib1bfcdc0c972aafc99116ed8c0511445 + I7978d2d800b4438d0644ae3df6bcac9c;
            tout_00082_00003    = fgallag_final_00082_00003;

            I9af399f27c8e2b62b7f3fc6481ef9318= I7adff505c50450a04f1717cac1adebe7 + If845af0d620024f04525244753ba5d18;
            tout_00083_00000    = fgallag_final_00083_00000;

            I171bb4ee9be2f92e4d82997108572426= I7adff505c50450a04f1717cac1adebe7 + Ie7820d1a242bc28c19ec32d2c91e47b7;
            tout_00083_00001    = fgallag_final_00083_00001;

            Ib13cd76c20fcaf95f26f4914380c4fcf= I7adff505c50450a04f1717cac1adebe7 + Id50f18f642f3b00ffa34986f78a0eae6;
            tout_00083_00002    = fgallag_final_00083_00002;

            Iafb219f1c8c6883e01fbfb4c887c8d6a= I7adff505c50450a04f1717cac1adebe7 + Ibc4eddc0f1768e9ec7e38e951a28ec42;
            tout_00083_00003    = fgallag_final_00083_00003;

            I94fc9b0bdd2b0a89a9f6351f1fdd4ff5= I699feb4382974a02b21cb387c13f7f3f + Icfef12499b53cd84f0aae067f30c17d0;
            tout_00084_00000    = fgallag_final_00084_00000;

            Ia9ceb45f33402293c162cef4037ba007= I699feb4382974a02b21cb387c13f7f3f + I1039bc43e88eee527d2ed6adb8c7d1ba;
            tout_00084_00001    = fgallag_final_00084_00001;

            I0fa4e12e62e8a30b3b8045143b344b4f= I699feb4382974a02b21cb387c13f7f3f + I5b64997d083769666741c794dd92fb7f;
            tout_00084_00002    = fgallag_final_00084_00002;

            Icec1c637d24ca277bb2e488257e92a40= I699feb4382974a02b21cb387c13f7f3f + I1c97fd1d21a31af8b5498a79b1a3e7b6;
            tout_00084_00003    = fgallag_final_00084_00003;

            Ie9aca08b988fad20904545fe070defd5= Idc99c3b23e49aca3c98f0685ea34441c + I83d71a89f35eb73265ee3e54184e1277;
            tout_00085_00000    = fgallag_final_00085_00000;

            Ie82304b2c8583f967649475e309e68fa= Idc99c3b23e49aca3c98f0685ea34441c + I3caf1211dcbcdc746a3e4c7fbbdae4a8;
            tout_00085_00001    = fgallag_final_00085_00001;

            I60da0fb8a2c0669d5f9037ae99b23565= Idc99c3b23e49aca3c98f0685ea34441c + I49f5f87662fbb540d72c94bfd1acd060;
            tout_00085_00002    = fgallag_final_00085_00002;

            Id8c19a3547c17ed513d2d857adc66885= Idc99c3b23e49aca3c98f0685ea34441c + Ie4f063eeaf7ee3f033e2a01ffaca623e;
            tout_00085_00003    = fgallag_final_00085_00003;

            Id74984743844e9495ea0f528a391f4b8= Ib67318fa6954ec8f3247927d34e74f8c + Ie45aaf966aa0a94803050b5f43d69e6c;
            tout_00086_00000    = fgallag_final_00086_00000;

            I9edcdd5b927b3f6b3a4c7cacebeb4a82= Ib67318fa6954ec8f3247927d34e74f8c + I9275bb36e58e0f17964e13ee7f027ab7;
            tout_00086_00001    = fgallag_final_00086_00001;

            Ic89597a95f50382cd3a2730896735d55= Ib67318fa6954ec8f3247927d34e74f8c + I1b6d20c64b9f23fb6c30f723546aa285;
            tout_00086_00002    = fgallag_final_00086_00002;

            Ibb7d203dfc75bf6211b09ab94877f93d= Ib67318fa6954ec8f3247927d34e74f8c + Ibb3d57d510cad00064a331f61f6400a2;
            tout_00086_00003    = fgallag_final_00086_00003;

            Id2f2e6837c83973cb2173454433acb88= I8774ce3f11362915c4331d1026e452dd + I80f2e8f6743e28e86e4d85b295e2f768;
            tout_00087_00000    = fgallag_final_00087_00000;

            I1259d5918f8d65b4b22ccfef22fe3afa= I8774ce3f11362915c4331d1026e452dd + I9bc2d5692474b8368c570d92835191b3;
            tout_00087_00001    = fgallag_final_00087_00001;

            Ib84e8c6e7fd9d7762e6e7e508d5ee40a= I8774ce3f11362915c4331d1026e452dd + I30080cc6c03bbe933165d266558a822c;
            tout_00087_00002    = fgallag_final_00087_00002;

            Ia032017912715abde99ffdf5ba732c5f= I8774ce3f11362915c4331d1026e452dd + I9485ae915474a31562ce358666d66245;
            tout_00087_00003    = fgallag_final_00087_00003;

            I55c310bfefb635448ef9c25c5d15987e= I2392b2d17ffed6073875fbe8e92534cf + Ifd958901d2ea2284f506e04a058012fa;
            tout_00088_00000    = fgallag_final_00088_00000;

            I92c0f229cf7fdb2cc0fe4d84f4d9b11d= I2392b2d17ffed6073875fbe8e92534cf + I1070940dc2ef6e8ee3d1227ec9ff3162;
            tout_00088_00001    = fgallag_final_00088_00001;

            I5570eb486d238fd96f9a59b174f5a22a= I2392b2d17ffed6073875fbe8e92534cf + Ia54b6f7044a831020e49f1bf48bc063a;
            tout_00088_00002    = fgallag_final_00088_00002;

            If6f01d24acf4a8b38bdbb1b366cd9a47= I3a4f0d3e32596ef05477f494768d4266 + I7c0f872988488ac69815d288885dfd2f;
            tout_00089_00000    = fgallag_final_00089_00000;

            Iff29fff36064aa4f9d339d4c62956e61= I3a4f0d3e32596ef05477f494768d4266 + Id2808e0f40992c79ead4da7c734e5b79;
            tout_00089_00001    = fgallag_final_00089_00001;

            I818d7cae6f1b80ac452dbfc073ccfe7a= I3a4f0d3e32596ef05477f494768d4266 + Ie71c7babb5d17378d40444b6bbd4e7a6;
            tout_00089_00002    = fgallag_final_00089_00002;

            I77ecfe991c6ec778495d7d5e5e442eca= Icd08ff59cf6be3ba97698dd55703339e + I75f9d3a41019dca3044a1c2cf7069662;
            tout_00090_00000    = fgallag_final_00090_00000;

            Ie7c6a56e8b6f7756bb5a24bdfd6a855e= Icd08ff59cf6be3ba97698dd55703339e + I6e7e27bb176196e4493bf9c45ca19719;
            tout_00090_00001    = fgallag_final_00090_00001;

            I9f9bc8eb8b2978a3dc529c34516fdf75= Icd08ff59cf6be3ba97698dd55703339e + Ia0977b79857bdbf058535c30e338c38a;
            tout_00090_00002    = fgallag_final_00090_00002;

            Ie3c0e5a4b00a92357a5d37e527d59b61= I985fb7ed22a8476ea322c9e3c2b3851c + I08e907b0619bec3ef2cf4cb3779e0794;
            tout_00091_00000    = fgallag_final_00091_00000;

            I9b9a9486420e7d4aa105c48dd50aa74d= I985fb7ed22a8476ea322c9e3c2b3851c + I64c4bb0d40d80ec52aab61ce46954f43;
            tout_00091_00001    = fgallag_final_00091_00001;

            Id12199a504f7aa298fffaaedd1aacc99= I985fb7ed22a8476ea322c9e3c2b3851c + I600ea1371a2be66430ac9534583b512b;
            tout_00091_00002    = fgallag_final_00091_00002;

            I813691fd8ea36626d32c8d2562163f32= Ib985709316b1b0a9d3fa3c1eaf6c641f + I1391018fb93372ccc2fcc08700e38b65;
            tout_00092_00000    = fgallag_final_00092_00000;

            I5fd3aaddc3eb8afeb82768b45e2d53d7= Ib985709316b1b0a9d3fa3c1eaf6c641f + I749b9c345f23aae03c595a2c76126ecb;
            tout_00092_00001    = fgallag_final_00092_00001;

            I1ac281eab6c7459e835fe992142b7857= Ib985709316b1b0a9d3fa3c1eaf6c641f + Ie230ba3c73808e102eee9e5868595e7c;
            tout_00092_00002    = fgallag_final_00092_00002;

            I49e5078c9161e8bee00fb76bc00b5288= Ib985709316b1b0a9d3fa3c1eaf6c641f + Ife5b9afdbb30c122b84d5378f9cb366d;
            tout_00092_00003    = fgallag_final_00092_00003;

            Ia697adf14616bf50d6e8178596b9fa7e= I4be898887dff6e2cebe53f135ece131b + I0982b8d7f99aceb8871c9c10448f54c5;
            tout_00093_00000    = fgallag_final_00093_00000;

            Iff3128a26dabe63b015dc6afc98a85a9= I4be898887dff6e2cebe53f135ece131b + I97e89a2ee18d2688d7c1a640318a1e0d;
            tout_00093_00001    = fgallag_final_00093_00001;

            Ifc04708ee5a7cc2b3f1850db778fa42e= I4be898887dff6e2cebe53f135ece131b + I94af4b6b9dc11935db54ba872889392d;
            tout_00093_00002    = fgallag_final_00093_00002;

            Ia405859c9dff67905b2e91bcbc06259e= I4be898887dff6e2cebe53f135ece131b + I27556d599dd1a27ee8f49e819ccbf29a;
            tout_00093_00003    = fgallag_final_00093_00003;

            I2fec8f62b28575e8f3af756db66fa232= I004db04f61fb57aba81e15cc015442b3 + I7362f08ed4e4ae309dfbfda112c56ad6;
            tout_00094_00000    = fgallag_final_00094_00000;

            I98e97c02477032ead66dc50f3f274e5a= I004db04f61fb57aba81e15cc015442b3 + I793ddbf6a5d026a57ab72984ca19deac;
            tout_00094_00001    = fgallag_final_00094_00001;

            I9f2dc5add3a4d1e6eb3116c741cd2f82= I004db04f61fb57aba81e15cc015442b3 + I3bdc5ba374f85dc61346e4868c41a6bf;
            tout_00094_00002    = fgallag_final_00094_00002;

            Ie122f7d8a48d7ad29d998b6a14b8e70f= I004db04f61fb57aba81e15cc015442b3 + Icce595233ce089eafcca3eae5e71e5f8;
            tout_00094_00003    = fgallag_final_00094_00003;

            Ib5576c996062391f44066d893dd5cb91= I8f7e3dfb2f728d4cd1e79b82b62b0406 + I88aedd7f52399f5fd435c3415f2218ca;
            tout_00095_00000    = fgallag_final_00095_00000;

            If931597aab866a74c3a3ffb1cd429583= I8f7e3dfb2f728d4cd1e79b82b62b0406 + Ibfe325e48511372569e0d98d9c4e70e3;
            tout_00095_00001    = fgallag_final_00095_00001;

            I79878bd69ed53785b8a5f025a2a00a4f= I8f7e3dfb2f728d4cd1e79b82b62b0406 + I28c3818247c7c6de11790f6692882b5a;
            tout_00095_00002    = fgallag_final_00095_00002;

            Iefb0a20652954fc2002154ea874c120a= I8f7e3dfb2f728d4cd1e79b82b62b0406 + Icc3cadf40c09be1a8c2847caf0e3e63c;
            tout_00095_00003    = fgallag_final_00095_00003;

            I646ca66e4e9f24b4fb75b38bf293b4cc= I991054370345e61638ddaf81785505bd + Ie317bbd70b9092b840c0f2713204fb9d;
            tout_00096_00000    = fgallag_final_00096_00000;

            I051f0d4c44123e3637b84a32c9a00a75= I991054370345e61638ddaf81785505bd + I8922cc37cde6ba132f632743113e42af;
            tout_00096_00001    = fgallag_final_00096_00001;

            I1876f9ec3f6f637ee40cdad7cc347f6f= I991054370345e61638ddaf81785505bd + Ia3d129fd297905bee180293c0c39d9ef;
            tout_00096_00002    = fgallag_final_00096_00002;

            Ic3d6b8dbec6cf92a9b6a17fb2f75dcd4= I991054370345e61638ddaf81785505bd + Ib43886d923b8c683004713ff25b2f90d;
            tout_00096_00003    = fgallag_final_00096_00003;

            I7d89f1db7b1015d34363ad781374de58= Ifa1f503965270d10e7a5c9a15576069b + I3521b10b97b0e74888ce385cfc772945;
            tout_00097_00000    = fgallag_final_00097_00000;

            Ife217ec4da1f1477bce034cb3545160f= Ifa1f503965270d10e7a5c9a15576069b + Icb2b390266bff241a688961136db0f51;
            tout_00097_00001    = fgallag_final_00097_00001;

            Idc5e5e98508c94b87a760f8eb36fad41= Ifa1f503965270d10e7a5c9a15576069b + I8bf8b0cf27a2654a0e7fdf3255945b67;
            tout_00097_00002    = fgallag_final_00097_00002;

            I9e72b0c823f297535f13a1b3072c2776= Ifa1f503965270d10e7a5c9a15576069b + I132d9671c582876568c0f7f5335f5227;
            tout_00097_00003    = fgallag_final_00097_00003;

            Ia81da7c58d6636ab70e0cf3e263a12c0= I24f773842a4742fb58d09cae45717b2f + I820fa56328e3919970dd64adb1d4d8e7;
            tout_00098_00000    = fgallag_final_00098_00000;

            Ibfc69ef08382c79e30cfafd89bfeff69= I24f773842a4742fb58d09cae45717b2f + I4cff1804df738cbf4f940c775236df9c;
            tout_00098_00001    = fgallag_final_00098_00001;

            I2d2afa9165b7121dc8289e9e6cdab5de= I24f773842a4742fb58d09cae45717b2f + I450c0d6ad5d3b1f18bb28e3a432b5442;
            tout_00098_00002    = fgallag_final_00098_00002;

            I065052693fd8ca87614feb60f7ef37c3= I24f773842a4742fb58d09cae45717b2f + I0859c80b42a8c60dade8f05d58ee3701;
            tout_00098_00003    = fgallag_final_00098_00003;

            I13344a81551374f665cbc17c7e94296a= I5bac7e0d778a547a0ae764fe259b6f7a + I68e5b12792a86dda0576742831d3b728;
            tout_00099_00000    = fgallag_final_00099_00000;

            If5a1d2de0715fa87d191ee5f48171676= I5bac7e0d778a547a0ae764fe259b6f7a + I512f57a40c7c8cb2f040bdde73e44ca3;
            tout_00099_00001    = fgallag_final_00099_00001;

            I02b256f74ee86b42ff1eba5e3d242737= I5bac7e0d778a547a0ae764fe259b6f7a + I58447d6ae49a6be2d043477a06f83df0;
            tout_00099_00002    = fgallag_final_00099_00002;

            Ic113fc051eefaef846f440e98f2f8913= I5bac7e0d778a547a0ae764fe259b6f7a + Ib3690ec149adde94343d3e617931a287;
            tout_00099_00003    = fgallag_final_00099_00003;

            Iabeab9bdd0bd82dd145218b563b5dac1= I255577ebee6768871df0224fc1db2db3 + I6c661048307c23c699d4b3636564de0f;
            tout_00100_00000    = fgallag_final_00100_00000;

            If9ce0a09e3a4e816dda002a24319ac0b= I255577ebee6768871df0224fc1db2db3 + I557ef77ce931535467a07a8d70145f55;
            tout_00100_00001    = fgallag_final_00100_00001;

            Ib5a7d72c36e41754033a64fbe0718784= I255577ebee6768871df0224fc1db2db3 + I41f2bf9ff00f983ad1298c8c83b041cb;
            tout_00100_00002    = fgallag_final_00100_00002;

            I41df12c7dee8526abf92b8e98965fa06= Ia7fb4af3d3529a32f902a52cf5598474 + I8be4be8471625db0749e6385f87d2dcc;
            tout_00101_00000    = fgallag_final_00101_00000;

            I83dfbd224e7465a6fd769e407182829a= Ia7fb4af3d3529a32f902a52cf5598474 + Ib451127b69a0a800332a712af77c6d29;
            tout_00101_00001    = fgallag_final_00101_00001;

            Ie57bba5092ec318456365b81b36aaa65= Ia7fb4af3d3529a32f902a52cf5598474 + Ib5414585cd6976cfce42e42190cc08d7;
            tout_00101_00002    = fgallag_final_00101_00002;

            Ibcf043d24474ab8c1002d15fde2d7da2= I2c98806141f064c9e92935b23a84ede1 + I7651176b0a74846108fbaabc5cc4900a;
            tout_00102_00000    = fgallag_final_00102_00000;

            I2e3385871c6ed8cf9519f273c8a19fda= I2c98806141f064c9e92935b23a84ede1 + Ie1e9326e4eee006ec07abb6bb7d269a5;
            tout_00102_00001    = fgallag_final_00102_00001;

            I664917b9f44515bf556d69ade4ca408c= I2c98806141f064c9e92935b23a84ede1 + I1ca59325ff30db83df5bf0a2cd9706b6;
            tout_00102_00002    = fgallag_final_00102_00002;

            I28deacdec0fbd0bce49b654c2620ac38= I5680847bc8d224fa4ed93b2fc0d841e1 + I8fd26d47ecd4cdd08294cf6133468d17;
            tout_00103_00000    = fgallag_final_00103_00000;

            Ibdfc4852c620f573f929584e6b816f35= I5680847bc8d224fa4ed93b2fc0d841e1 + I38e2dbba093928b874d447362d89b291;
            tout_00103_00001    = fgallag_final_00103_00001;

            I5a69b2bbb63ab919ea2270503cd326f1= I5680847bc8d224fa4ed93b2fc0d841e1 + Ie2f5b03f3b136e651b8aba92a30d298a;
            tout_00103_00002    = fgallag_final_00103_00002;

            I2eccd8d60a19481fa595566f51c7aa4e= I365254279ebb10dd7ba0b3482d5e34cd + I0c1e22375d5e023c24519901b92eceb5;
            tout_00104_00000    = fgallag_final_00104_00000;

            I49eb4bba42440657fe04b711eedfa67f= I365254279ebb10dd7ba0b3482d5e34cd + Idd1b6014de2f053554ed09c29bf3e640;
            tout_00104_00001    = fgallag_final_00104_00001;

            I9ed8323951af0de78ae89153cbf9e9eb= I365254279ebb10dd7ba0b3482d5e34cd + I97f2813ec39bbf1513faf66b3e38838a;
            tout_00104_00002    = fgallag_final_00104_00002;

            I1d00816529836546b514f54b1275d39e= I365254279ebb10dd7ba0b3482d5e34cd + I0a3323aac825506435068f6746aee974;
            tout_00104_00003    = fgallag_final_00104_00003;

            Icc58b9a24fb9ef7e8fa5f13a2cc0a0cb= I365254279ebb10dd7ba0b3482d5e34cd + I312ce79a8dd2ce3d37c930d42640509b;
            tout_00104_00004    = fgallag_final_00104_00004;

            I9339aef608b029175b488e82f5b3f1bb= I57bf4ad773cc058ae1bb7b1911dc3174 + Id60cbf534604e5dba988050ef5abe625;
            tout_00105_00000    = fgallag_final_00105_00000;

            Ibd2f24860b701ab46e0c436d774e43f9= I57bf4ad773cc058ae1bb7b1911dc3174 + I40e99289d5762e77a3766eb8251eef00;
            tout_00105_00001    = fgallag_final_00105_00001;

            I37fe66ec8927f27f646b304500400ccf= I57bf4ad773cc058ae1bb7b1911dc3174 + I9e09c25be9f877c1e1aaf79bf12c7943;
            tout_00105_00002    = fgallag_final_00105_00002;

            I4bd6a48f494cf633a857b8ccbd67af68= I57bf4ad773cc058ae1bb7b1911dc3174 + I30253dc91301ca27b5732312c01145e0;
            tout_00105_00003    = fgallag_final_00105_00003;

            Icd7a7566438dc67e77f138ac814844f0= I57bf4ad773cc058ae1bb7b1911dc3174 + I467d5e2554ef25873e0b44e947ee0011;
            tout_00105_00004    = fgallag_final_00105_00004;

            Ic3d4239413333883dd926c7a42c0a87f= I57072dfb29c4a3d2e2b40e46e62f0d95 + Ia66c399023e500ed67197dcf236f5d42;
            tout_00106_00000    = fgallag_final_00106_00000;

            Ib8298d1ead61bc00eb31599b3087d769= I57072dfb29c4a3d2e2b40e46e62f0d95 + Ic66af6c3c0268cfb0e9f0776c4f4e961;
            tout_00106_00001    = fgallag_final_00106_00001;

            I23dbe33ce46f94d3dff1e6d391305609= I57072dfb29c4a3d2e2b40e46e62f0d95 + Icaae0fb0f460f68d690ab00697355a49;
            tout_00106_00002    = fgallag_final_00106_00002;

            I138286817f424c76e8a4f30540b0530b= I57072dfb29c4a3d2e2b40e46e62f0d95 + I0d66aa55747362354aa81d96057bc4c2;
            tout_00106_00003    = fgallag_final_00106_00003;

            I30c645a78b900306864a1ab23e923bde= I57072dfb29c4a3d2e2b40e46e62f0d95 + Ice73b514709469fd21cd254bf4ceadd9;
            tout_00106_00004    = fgallag_final_00106_00004;

            Id88681d0fe3ea62530166938503db05a= Id8cafb6f76321bdaba9711133be7be99 + I54cfd68212d97a2cc8241ef429429453;
            tout_00107_00000    = fgallag_final_00107_00000;

            I808008402174fa4edf42783135c0c3a9= Id8cafb6f76321bdaba9711133be7be99 + If8aa3ec1b5a4a3c122da82467be917da;
            tout_00107_00001    = fgallag_final_00107_00001;

            I3ad4d02ea2e52a49b6fa4f1da9b58149= Id8cafb6f76321bdaba9711133be7be99 + I53309409a6059c3bd39f037c23ec3458;
            tout_00107_00002    = fgallag_final_00107_00002;

            I39486eecb7bbfecf26573a7a5876feb9= Id8cafb6f76321bdaba9711133be7be99 + I7e28234bdf66ab5489d36d15678db797;
            tout_00107_00003    = fgallag_final_00107_00003;

            I21e8ea20029fb2cb62103405b81b21b0= Id8cafb6f76321bdaba9711133be7be99 + I45ba06a6d6f00c174b1439a6f226a085;
            tout_00107_00004    = fgallag_final_00107_00004;

            Id0b67fa451e276889e02779ddb667904= I6344e71ca2b0fd39d36caedd889c3085 + I786dfcaa131b99c254aaff15bd2c2b6d;
            tout_00108_00000    = fgallag_final_00108_00000;

            Ic328d25a58ec4559b753da3bcff938de= I6344e71ca2b0fd39d36caedd889c3085 + Idad14b6383b9af54eb35e72ff3d10035;
            tout_00108_00001    = fgallag_final_00108_00001;

            I49c44c2f2522e086c2db8a00647ba35c= I6344e71ca2b0fd39d36caedd889c3085 + Ic8a272f82736fd599fb3250e970edf9b;
            tout_00108_00002    = fgallag_final_00108_00002;

            Id4152a04385391294f4b8a18df2cb9ee= I0c99a68e0bed90afce18807acf7d55bb + I3d6a685a1913bd8be01fddbce1edec2e;
            tout_00109_00000    = fgallag_final_00109_00000;

            I5b0213a3df61e94fd0b744a8141f7502= I0c99a68e0bed90afce18807acf7d55bb + I8c0069e8756bcff203ce21ae3170aa42;
            tout_00109_00001    = fgallag_final_00109_00001;

            If0ad11ed403cbbed68614b01e2a3793e= I0c99a68e0bed90afce18807acf7d55bb + I5b9710b16effc8bf0695517c6e651836;
            tout_00109_00002    = fgallag_final_00109_00002;

            Icfa1170bc73534bee13778bc3b88a2f7= I1c95650979c86310ae2a949961c9db11 + I57ac487adc18165136e9b3c7c50f95ad;
            tout_00110_00000    = fgallag_final_00110_00000;

            Ife1bd938a0dd06d8d3cf30ff41a303b2= I1c95650979c86310ae2a949961c9db11 + Ib484aa64b795f7e36198b800f302164f;
            tout_00110_00001    = fgallag_final_00110_00001;

            I4a09cb1b99b476fa6fae0bc44c41a041= I1c95650979c86310ae2a949961c9db11 + I038b42a83025f5eaebf45799d1ebe7b0;
            tout_00110_00002    = fgallag_final_00110_00002;

            Ie08cf323944813e4b9e2d59a680ffe8d= I04eaefa5d133e53494fc270b07be7043 + I7097c9518bb3351818b96f31ed49c6d3;
            tout_00111_00000    = fgallag_final_00111_00000;

            I85fc307fb52d58550eeecd33bc4207a4= I04eaefa5d133e53494fc270b07be7043 + I41af7e4c97fc04154fe6de66b82499f5;
            tout_00111_00001    = fgallag_final_00111_00001;

            Id00dd13741fe621d0a240bdc92318f55= I04eaefa5d133e53494fc270b07be7043 + I73ddd7cf9272ceab5a663e2244e72d7e;
            tout_00111_00002    = fgallag_final_00111_00002;

            Idc8e891fd432df75a4eb133ce35ecec4= I4a64fa2412eb8058c2dfd9351d7b297d + I2f9e56d570e72714a06c59aa9e4334c0;
            tout_00112_00000    = fgallag_final_00112_00000;

            I2a51cada20cbd14f7d5a289599e68b53= I4a64fa2412eb8058c2dfd9351d7b297d + Ida5b16851dc06534844a0b037d74feb3;
            tout_00112_00001    = fgallag_final_00112_00001;

            I65a701d1e083e501544bb0fce24f0c4e= I4a64fa2412eb8058c2dfd9351d7b297d + Ia48f0029e9e76386f3dd70aacd9adbfa;
            tout_00112_00002    = fgallag_final_00112_00002;

            If3020a9109ac83274b5bafac18d176de= I4a64fa2412eb8058c2dfd9351d7b297d + I16507fab8f9076bfeb419896fa7cdc1d;
            tout_00112_00003    = fgallag_final_00112_00003;

            Iaa6bd55038c2ae911e4df08f707c55f5= Ie8bb2fcb752c6a33254963d1ebb4130d + I58f0b81a46549cab8e74ecbc285df23a;
            tout_00113_00000    = fgallag_final_00113_00000;

            Id49065cedf20e13abac8971534bb8b0e= Ie8bb2fcb752c6a33254963d1ebb4130d + I37998a91d20db2248ebdd8e661d42f70;
            tout_00113_00001    = fgallag_final_00113_00001;

            I0bb64952d77b59803a561e14b950b9b1= Ie8bb2fcb752c6a33254963d1ebb4130d + Ib4695d4389db72c5ac7e31809072c290;
            tout_00113_00002    = fgallag_final_00113_00002;

            I01e295a6ab88c6f34b44efcc32a23233= Ie8bb2fcb752c6a33254963d1ebb4130d + I3dd1f28cf199299aba54e47a429c9b11;
            tout_00113_00003    = fgallag_final_00113_00003;

            I2acf864d587b7681ca0fb6e2e2bea617= Iac05b7e3ae18f948b72c356ccfb8000f + I05eadf11cdc6c2f2b021e33f2438fa49;
            tout_00114_00000    = fgallag_final_00114_00000;

            Idfd0410b37713e8808f8bea81e2af881= Iac05b7e3ae18f948b72c356ccfb8000f + I1171dc208d5db1024dc3f09a90c78ca0;
            tout_00114_00001    = fgallag_final_00114_00001;

            I02861f333b5adfd4962356cdf5a11f23= Iac05b7e3ae18f948b72c356ccfb8000f + I3d601db540da359ae4d22f960d3d5af8;
            tout_00114_00002    = fgallag_final_00114_00002;

            I4ddbc3daa65b111cb0d45e13d62cc292= Iac05b7e3ae18f948b72c356ccfb8000f + I49d9203dc6f8c17f17383e8f7e01f005;
            tout_00114_00003    = fgallag_final_00114_00003;

            Id363d158feb8fec19b5f3d73d84f0068= I27da3f75cca6c49e55db90306aa68e94 + I72db05084d30d7c59ba1cb06d3b09400;
            tout_00115_00000    = fgallag_final_00115_00000;

            I8ec9b7a6e65e727abbed336ce240a4cf= I27da3f75cca6c49e55db90306aa68e94 + I8d4e3962525c424786ae822a6981a5e6;
            tout_00115_00001    = fgallag_final_00115_00001;

            I128fa1e99b7eb9b6905c2cfd26b95ab4= I27da3f75cca6c49e55db90306aa68e94 + Ica4ec1647bdb5a3aad6db6b447bd7995;
            tout_00115_00002    = fgallag_final_00115_00002;

            I93d459b6da42a205c91c48622f0c5032= I27da3f75cca6c49e55db90306aa68e94 + Ibeec86c75d950ee00dd63a2930f08a24;
            tout_00115_00003    = fgallag_final_00115_00003;

            I1243cc8d5dddf7dd65b40c0b3b958b9e= Idc7fed723190098341225fe01ba65ced + Ic95668328a2121027436f682bac50b9c;
            tout_00116_00000    = fgallag_final_00116_00000;

            I238df7e09d42bc93a972da349a00f511= Idc7fed723190098341225fe01ba65ced + I82a14e1ee4723e7d9a13c1f2b8b13691;
            tout_00116_00001    = fgallag_final_00116_00001;

            Ic658b2afdc7331653fc84d6372d47418= Idc7fed723190098341225fe01ba65ced + I47b2438c3680b2d816168df37d7c491c;
            tout_00116_00002    = fgallag_final_00116_00002;

            If39be111eb101c9c983fe0baa9a1cb18= Ife9065805598960919ee4f14c3cc6fd4 + Id683d693cd50645c3d6d657aa1c8bdb2;
            tout_00117_00000    = fgallag_final_00117_00000;

            I9d19d5b7d8b256c1707de97a4549c458= Ife9065805598960919ee4f14c3cc6fd4 + I461398638cb8280f1779915298540b00;
            tout_00117_00001    = fgallag_final_00117_00001;

            I6c2fffe204091f7f64aea16b0ac98769= Ife9065805598960919ee4f14c3cc6fd4 + I5983bf2c6c90b872ee6cf58b5e520311;
            tout_00117_00002    = fgallag_final_00117_00002;

            Ic4ba4d2e5c12d9f1dd233d64929f1072= I717c5c2d6a2be61593492ae5f17a112f + I2b49d74cb130542f2ca99534e2c513b1;
            tout_00118_00000    = fgallag_final_00118_00000;

            Ia9dec5831998d472d11429e5a7e60ed8= I717c5c2d6a2be61593492ae5f17a112f + Idbea892c8109117f90b453efe8ae25af;
            tout_00118_00001    = fgallag_final_00118_00001;

            Ieaaf52c1e663f260292bc1529718d681= I717c5c2d6a2be61593492ae5f17a112f + I6745cacecb7ee86cf3c7ad7eeee6048f;
            tout_00118_00002    = fgallag_final_00118_00002;

            I37061896a09588a73445deed73d3746c= I4c31fa8e6eb648439cdae1de1afe0d6f + Ifd77e040c5f82790b1d5636a42fca602;
            tout_00119_00000    = fgallag_final_00119_00000;

            I02f25b80945b6f58193fb37add3da2d8= I4c31fa8e6eb648439cdae1de1afe0d6f + I28aa517220bf597cf898660f698ef19d;
            tout_00119_00001    = fgallag_final_00119_00001;

            I19045602bb77f12666ebd44f813db2c5= I4c31fa8e6eb648439cdae1de1afe0d6f + Ib9672d20643d856ff31905ab14c0ac87;
            tout_00119_00002    = fgallag_final_00119_00002;

            I4abdc8d5318d2922696a8aaee46ffa59= Iead549a9af27f1fced7d9c36e7b5c3f5 + Ic28b148967a5b3d05409976fa9001ac8;
            tout_00120_00000    = fgallag_final_00120_00000;

            Ie139f2048f346d82623c8fc6d40c9acc= Iead549a9af27f1fced7d9c36e7b5c3f5 + Ie81315a3a14a5ef879d8e3f405936365;
            tout_00120_00001    = fgallag_final_00120_00001;

            I8d99c96e203fafc81d13ce5aee925d75= Iead549a9af27f1fced7d9c36e7b5c3f5 + Ia605d14205926b3edc6d1c2f69f70ac0;
            tout_00120_00002    = fgallag_final_00120_00002;

            I37b0bdeb3cc54d6a97720c4912c67832= Iead549a9af27f1fced7d9c36e7b5c3f5 + Id555c88cf7f0904db74d45cc75c8f5d6;
            tout_00120_00003    = fgallag_final_00120_00003;

            I08257e9e6c74c60448e22fb9855f0825= Iead549a9af27f1fced7d9c36e7b5c3f5 + Ib9dfea1f34a120eda30d5bd919365a6a;
            tout_00120_00004    = fgallag_final_00120_00004;

            I32188cca2fc715698fc05b0fc6506434= I10422eb79364e7d0e21e1643d9060331 + I1a5f22b4e326d1684c0a8c7a7e754ab4;
            tout_00121_00000    = fgallag_final_00121_00000;

            I88f1cbab9b8fa3802345f745d024931c= I10422eb79364e7d0e21e1643d9060331 + I2c1f2476efe593829ade470fe8ec2526;
            tout_00121_00001    = fgallag_final_00121_00001;

            Idf548c0e78bd221bf9f612f27002fae0= I10422eb79364e7d0e21e1643d9060331 + I8daf79a0a2ee1bac7f055af441539fa4;
            tout_00121_00002    = fgallag_final_00121_00002;

            Iedfd2e04f5740d283388639dde3ecdb5= I10422eb79364e7d0e21e1643d9060331 + I63f82f075d53205b5b556c0054f1a0b8;
            tout_00121_00003    = fgallag_final_00121_00003;

            I7088c83eacff6f1dfb134f79d469c8f1= I10422eb79364e7d0e21e1643d9060331 + Ia7bf82c9e5ca4467b5e50beeaeb975e9;
            tout_00121_00004    = fgallag_final_00121_00004;

            I6f8431671331f4ca7ea19656e0677cd4= I914cb87eba8baa40cd515334e59f26b2 + Iac3cb5b4481687fcf430c8bf52cfb74d;
            tout_00122_00000    = fgallag_final_00122_00000;

            I1e31259e267e04920cbbd16bd7aa18bc= I914cb87eba8baa40cd515334e59f26b2 + Ia17295aec0a40c2b46a595dacfede2d5;
            tout_00122_00001    = fgallag_final_00122_00001;

            If54d9f8088e67e44cfa3026f5a520fd7= I914cb87eba8baa40cd515334e59f26b2 + I0d96336eb4d5071d7e1d350e86513b25;
            tout_00122_00002    = fgallag_final_00122_00002;

            I6fd2c0746407b23aec5dff1e083f5fca= I914cb87eba8baa40cd515334e59f26b2 + I2587a5800a5a9ffeabc4dca503e3d964;
            tout_00122_00003    = fgallag_final_00122_00003;

            Ib2147a19b44d361da628a628fbfaa988= I914cb87eba8baa40cd515334e59f26b2 + I327c9acb8934729b4ea5486787afa2e8;
            tout_00122_00004    = fgallag_final_00122_00004;

            Ie804d1f4b241a2de3e9d9c7c876d914a= I32ed679af4ab759901aee43c9d93eb67 + Ib65ff82aff398f6ff7ba711a36f41ee4;
            tout_00123_00000    = fgallag_final_00123_00000;

            I6cd1e6db57e06d8f5e60a31f48ae4809= I32ed679af4ab759901aee43c9d93eb67 + Ic2b20168744fafbe15037ed7fa83da72;
            tout_00123_00001    = fgallag_final_00123_00001;

            I3e0e8832d5338423284ac4b2a0c5f3f5= I32ed679af4ab759901aee43c9d93eb67 + I20beb3fdbe91936f74a200cd8ec9817b;
            tout_00123_00002    = fgallag_final_00123_00002;

            I6ac006d79e95e222cdc66754b67a08ed= I32ed679af4ab759901aee43c9d93eb67 + I83292bcda4645233d8e8a1dfe8e5f60b;
            tout_00123_00003    = fgallag_final_00123_00003;

            I29087dda1a527842aeb3d35d66c853cb= I32ed679af4ab759901aee43c9d93eb67 + Ieddef08050c38d07e5d38f5bb7b099c0;
            tout_00123_00004    = fgallag_final_00123_00004;

            Ia67e5920bbac700dfee52cd96b15963e= Id376dfa5141402f4d41a8858180ed87e + I5b53fd45210b92703cb10d583f471ab9;
            tout_00124_00000    = fgallag_final_00124_00000;

            I1f6ecd894d90547f661e7a3888d048bb= Id376dfa5141402f4d41a8858180ed87e + I74b3c9dd3a8168aacd4369b9ff68fdfd;
            tout_00124_00001    = fgallag_final_00124_00001;

            I3112e793c6e79e1f5da2776e69a34e3c= Id376dfa5141402f4d41a8858180ed87e + I39f9e8430db114991bfb27cc46ef3e39;
            tout_00124_00002    = fgallag_final_00124_00002;

            I79152f32b45ed5b4a5302f6460707b01= I98a384bc62ee03f5ad7df20ef2d9af95 + I7095040b38bf9d6b5229c11d2a0d7c57;
            tout_00125_00000    = fgallag_final_00125_00000;

            I3d16e7d6b190639b88a217f19ac63233= I98a384bc62ee03f5ad7df20ef2d9af95 + Ibec442c099da091afcf75a7c970bf8ea;
            tout_00125_00001    = fgallag_final_00125_00001;

            Ia1be780c686163cea54b62d6ede72dc6= I98a384bc62ee03f5ad7df20ef2d9af95 + I56aa548618a4a15e9a35e04f5eeb823f;
            tout_00125_00002    = fgallag_final_00125_00002;

            Ic398c31a2a6ca89d0236534589a5919b= Icfed259ca2bb2732d8e0c26ef67cd4cf + I2c487770d606451440eecf358202db32;
            tout_00126_00000    = fgallag_final_00126_00000;

            Ie91c3202bc957b350d1915000564392f= Icfed259ca2bb2732d8e0c26ef67cd4cf + I143f5e324716a94d24ada126886bf895;
            tout_00126_00001    = fgallag_final_00126_00001;

            I687957f5300b0d4f50d6893cc556bf25= Icfed259ca2bb2732d8e0c26ef67cd4cf + I1908897b529ca04df7e7da395be4a8ce;
            tout_00126_00002    = fgallag_final_00126_00002;

            I7816b368e8e8b8dd69383b2c9327120d= I20861535c450d6e6bf11c45dac120454 + Ib1f1aef6c0a9291553b62fd555feb2e7;
            tout_00127_00000    = fgallag_final_00127_00000;

            I5f021f4a664205afbe0761af4c8914f1= I20861535c450d6e6bf11c45dac120454 + I1ea33707e40a2e41513fdb3118371437;
            tout_00127_00001    = fgallag_final_00127_00001;

            I69728004b59b5206a03a8e2087834f7d= I20861535c450d6e6bf11c45dac120454 + Ib2bbd59cd6098608ed53ac556036534f;
            tout_00127_00002    = fgallag_final_00127_00002;

            Ibbe1d623f8f5f3aa7fc70197acc6df5e= I013929385ad819ddfcfcc59c22902ee3 + I118726375ca9381e45f001965fcefc5b;
            tout_00128_00000    = fgallag_final_00128_00000;

            I4cb9f74288811592fd97fdff52bd6fe7= I013929385ad819ddfcfcc59c22902ee3 + Ia7520053a7c4a94437c6a780b03a28a5;
            tout_00128_00001    = fgallag_final_00128_00001;

            Ibb471dbccd39d41e951e98348812e343= I013929385ad819ddfcfcc59c22902ee3 + I42455e7e4d0c63f97702d204d18a446e;
            tout_00128_00002    = fgallag_final_00128_00002;

            I7f37d68f8ddcf8b4d5e99fb51eada873= I013929385ad819ddfcfcc59c22902ee3 + If004552b2047ab1cf23bb50375460b01;
            tout_00128_00003    = fgallag_final_00128_00003;

            I72ded7153883418a712ef967439d2159= I34fffcb07fe82f11fe142f7c37f39155 + I88bd8012c93dd9e2ed52ea5e9b8b0004;
            tout_00129_00000    = fgallag_final_00129_00000;

            Ie071e08299bff6bbdbe1f84703aaec08= I34fffcb07fe82f11fe142f7c37f39155 + I7e685b06df8a8c2ac351fa9f9b76a81d;
            tout_00129_00001    = fgallag_final_00129_00001;

            I1b79aa38a39ccfc839260af89aa78e7a= I34fffcb07fe82f11fe142f7c37f39155 + I2603e0b8b93f6680e44c9c8883f6512c;
            tout_00129_00002    = fgallag_final_00129_00002;

            I7384296e4190d83fb9d9a92cf965125b= I34fffcb07fe82f11fe142f7c37f39155 + If97092e1e2147de199c94a23831cf6b9;
            tout_00129_00003    = fgallag_final_00129_00003;

            Ie03034ce6233ca24effe53a2c0c8f6f3= I61ca60fde05ed88cce714dcd8c13b827 + I0f6cb7a5a31d6f2f6178632c0c898bc6;
            tout_00130_00000    = fgallag_final_00130_00000;

            Ic298f77f42fc1d41cce684790036ecfe= I61ca60fde05ed88cce714dcd8c13b827 + I4c6d3d6fc2d10066a744fdd9405a7902;
            tout_00130_00001    = fgallag_final_00130_00001;

            I805269f95afbeb6b93182f68868d08eb= I61ca60fde05ed88cce714dcd8c13b827 + I716ee53e79883f69aa045380a357e913;
            tout_00130_00002    = fgallag_final_00130_00002;

            I881328804c45b06767af51e11182b27b= I61ca60fde05ed88cce714dcd8c13b827 + Ibf74a4dfaab7f7f538d2b5fac7394b63;
            tout_00130_00003    = fgallag_final_00130_00003;

            I958993626e6e44e12f7c1e8026914680= I4907dd45c158dc7e0041c64f1fb388f6 + Ifbe479e5cab3cba43444bec1e12e72a0;
            tout_00131_00000    = fgallag_final_00131_00000;

            If31528d1fc3a083ebc364e75cdd9c71f= I4907dd45c158dc7e0041c64f1fb388f6 + I62fdc8936121a2707d94cf3bd6e660ac;
            tout_00131_00001    = fgallag_final_00131_00001;

            I4703b8d5a9033027889bfa8685e09e4f= I4907dd45c158dc7e0041c64f1fb388f6 + I42c1d469ff97913cbf15e3ebee6fdfa8;
            tout_00131_00002    = fgallag_final_00131_00002;

            I22d8e84d2db4b07111b7fdc6eef34cc8= I4907dd45c158dc7e0041c64f1fb388f6 + I991a7a7d562eb0a8b4b8d8f008ef2225;
            tout_00131_00003    = fgallag_final_00131_00003;

            I8b7c6df3b5ea575caab7820c95974608= I2c8f6a9b9f655b317bb0af4d60fdbc4b + I8c2e0c83a8204d6b21e0e3e458d56f05;
            tout_00132_00000    = fgallag_final_00132_00000;

            Ia8aa76bccf7eb310a9356e8b7ea1609d= I2c8f6a9b9f655b317bb0af4d60fdbc4b + Id435b68afb53bef4afc7b70a9512e955;
            tout_00132_00001    = fgallag_final_00132_00001;

            If9de547bf469b8424f1625e990f72b04= I2c8f6a9b9f655b317bb0af4d60fdbc4b + I56d1025271f1f7704a40dd7f0df02b0b;
            tout_00132_00002    = fgallag_final_00132_00002;

            I27d51b2015ea9af9bc345adabdb07b6f= I2c8f6a9b9f655b317bb0af4d60fdbc4b + I64c3d7be41abaa17d6992f9af8e72789;
            tout_00132_00003    = fgallag_final_00132_00003;

            I93dddce2a0dc01ecb3039fac5cf04011= Ic7dff631559304ec59f0696c66436d62 + Ia1499972c4995268acd828c1289f353d;
            tout_00133_00000    = fgallag_final_00133_00000;

            I746da2c1d5a620eb7e749f72f0f04a06= Ic7dff631559304ec59f0696c66436d62 + I0071f2168787bd42ab7f2370aed9d0f5;
            tout_00133_00001    = fgallag_final_00133_00001;

            I1e15f8d6fdb4ac732768d0cf73af829e= Ic7dff631559304ec59f0696c66436d62 + I4600963866dcb9bbea2515c805f885cb;
            tout_00133_00002    = fgallag_final_00133_00002;

            Ib719e667d7ba857f4f7432a245f4a30f= Ic7dff631559304ec59f0696c66436d62 + Icb91e63ebabc7a75a54eb7c731df4fa0;
            tout_00133_00003    = fgallag_final_00133_00003;

            I4c6eec4a0c46e4f5d7c9734df48a16bb= I6a239d3e55b4a9a3be9989a85bbec545 + I3d1dd8b9c7c6d3913f7ac369ad7e625c;
            tout_00134_00000    = fgallag_final_00134_00000;

            I95623ec1fd5516040a9492aae0fc2b70= I6a239d3e55b4a9a3be9989a85bbec545 + I6261e0d339762cb2364421e6b87086cb;
            tout_00134_00001    = fgallag_final_00134_00001;

            I69017b49c11de463fe6d881e5c96a1aa= I6a239d3e55b4a9a3be9989a85bbec545 + Ib235af5b28d56f24372d3f0af816f2c2;
            tout_00134_00002    = fgallag_final_00134_00002;

            I4fb9ed32471aa614ce6923f6a2279b36= I6a239d3e55b4a9a3be9989a85bbec545 + I673d1d0d0daab99bd940c46cc14ef55a;
            tout_00134_00003    = fgallag_final_00134_00003;

            I2f0bc217c8a39d71adc1fc45c10b81c3= I630f905e55f08e7d1569a08e937ad216 + I79fe46308b93fbb24245fe1c75edf4a5;
            tout_00135_00000    = fgallag_final_00135_00000;

            I0f1c6bb577ea2b8b2ab636e64378544b= I630f905e55f08e7d1569a08e937ad216 + I31e5b2cdc3dc571eafa37510076bcc64;
            tout_00135_00001    = fgallag_final_00135_00001;

            I7a248af9d606c566e03977e985c280e0= I630f905e55f08e7d1569a08e937ad216 + Ia9e102d8679943c079f16c0228f0f0d1;
            tout_00135_00002    = fgallag_final_00135_00002;

            I0bf9d47bff47277de1e72518e8d88362= I630f905e55f08e7d1569a08e937ad216 + I62cadbd70b07a6a7a2974c7c392696b3;
            tout_00135_00003    = fgallag_final_00135_00003;

            I24b6f4f68f291dc50caf03dc902282cf= I8d13eb3669785c4279c685763d4f3fad + Ia8d3667adc34b2b50acf7edb970538d8;
            tout_00136_00000    = fgallag_final_00136_00000;

            I79335b28eea15735f760b7a8b803e93a= I8d13eb3669785c4279c685763d4f3fad + If9f2a53dbf6e9b9a335a7657b7a2b468;
            tout_00136_00001    = fgallag_final_00136_00001;

            I0b14b34b06cfa90539c2abca5639abec= I8d13eb3669785c4279c685763d4f3fad + I68c85727adecde0aa8aa66ed08c4b502;
            tout_00136_00002    = fgallag_final_00136_00002;

            I26878777354945712f834740b17dabcb= I8d13eb3669785c4279c685763d4f3fad + Icd8257d7f53d93db989eb56eaeb7e593;
            tout_00136_00003    = fgallag_final_00136_00003;

            I6cc5daed4de5950c02c0a57b993e22fc= I25a6f3de9a9a01cbbdd32ed848561aa4 + I03bea609a189246a2375b355df47cf81;
            tout_00137_00000    = fgallag_final_00137_00000;

            I52c382d5b0c4829127c011fae402ce04= I25a6f3de9a9a01cbbdd32ed848561aa4 + Iaec2f15665e83416bc140890f3cdde9a;
            tout_00137_00001    = fgallag_final_00137_00001;

            I46ea9871e867034daa2d0501038f15e0= I25a6f3de9a9a01cbbdd32ed848561aa4 + Ia7046faae1ab05978e4b32bd44049fb9;
            tout_00137_00002    = fgallag_final_00137_00002;

            Ibb8a202599550e87831647a93a14181a= I25a6f3de9a9a01cbbdd32ed848561aa4 + I05931ceae6eff26e5a66a44a54d628ae;
            tout_00137_00003    = fgallag_final_00137_00003;

            Ibb79f2ce0b6028ebb638fc6661444cf1= Iba3dd4b2c2c85c4cfe770d9b52ef4634 + Ia784f35a5a46837b69eb048dabf84052;
            tout_00138_00000    = fgallag_final_00138_00000;

            I0d0c07d65eda2eee01df9c330c0d6f4a= Iba3dd4b2c2c85c4cfe770d9b52ef4634 + Iab354cc9ac1173335c0efeef694f3567;
            tout_00138_00001    = fgallag_final_00138_00001;

            Ie6940736944bac9be609b8d58b2cb13c= Iba3dd4b2c2c85c4cfe770d9b52ef4634 + If3a79ede332c39a8d2a276de833242f6;
            tout_00138_00002    = fgallag_final_00138_00002;

            I472a71363435cb3ec054e00f9123ae64= Iba3dd4b2c2c85c4cfe770d9b52ef4634 + I306fec0aa68a0396053a6e0fa1cda38f;
            tout_00138_00003    = fgallag_final_00138_00003;

            I553223e9166dcbddd1a51d0f92d68f28= Ie1b744387b5200a504e4874e14d2f282 + Ic8d47ff5d6c31601a57df868da78c2d4;
            tout_00139_00000    = fgallag_final_00139_00000;

            I495309d795905a53b0a3d3daa4f1f9d0= Ie1b744387b5200a504e4874e14d2f282 + I25c324feaca84e80f58075597e8c448f;
            tout_00139_00001    = fgallag_final_00139_00001;

            I21d358fd7673c4392f4e4b3d3a858b2c= Ie1b744387b5200a504e4874e14d2f282 + If64aa8c220b9ab6652e081da7e404e80;
            tout_00139_00002    = fgallag_final_00139_00002;

            Ia1a60175112362f015c5531f7c48b90b= Ie1b744387b5200a504e4874e14d2f282 + Idee8c8144207d676d1f2f9064bbdff45;
            tout_00139_00003    = fgallag_final_00139_00003;

            I5644ece811bddcec04c9e3559c86109d= Icf76cb69aedf4db01cd3444f4c4ba471 + Ib504b808f724ca6032e7c746517cd4fd;
            tout_00140_00000    = fgallag_final_00140_00000;

            I37d2f9d3f05cb90e2d45bd578299885c= Icf76cb69aedf4db01cd3444f4c4ba471 + Ic308a5413f38b96d244cac3b0bc9462c;
            tout_00140_00001    = fgallag_final_00140_00001;

            Ie7d10f3c0f8b0add66d2cdd4435ccc88= Icf76cb69aedf4db01cd3444f4c4ba471 + Ia4131464996aabab8aae1db85f6a50e4;
            tout_00140_00002    = fgallag_final_00140_00002;

            I3c37396a1cef2f9e42b8ccc126db6eda= Icf76cb69aedf4db01cd3444f4c4ba471 + I5855124d566af739caa6511f8598f2c5;
            tout_00140_00003    = fgallag_final_00140_00003;

            I2f82390734079b8d289d48a6682cc624= I4857b5b50556c8e7fff4b2d3e08e4b28 + I8edbe77bacf1975e014faeee6b861980;
            tout_00141_00000    = fgallag_final_00141_00000;

            I9061728c3163ae684e8c5aec3e807868= I4857b5b50556c8e7fff4b2d3e08e4b28 + I1338d211b5d2d409bfe0df76d2ca2701;
            tout_00141_00001    = fgallag_final_00141_00001;

            I672d7ecc28a788c2602aff76187aa568= I4857b5b50556c8e7fff4b2d3e08e4b28 + I75838ca09e301b8e1301cbf603a1f8c2;
            tout_00141_00002    = fgallag_final_00141_00002;

            I660b2fe99cd0bcaac34e9540118b54bc= I4857b5b50556c8e7fff4b2d3e08e4b28 + I50729db4a8e04f18979707df14cb2419;
            tout_00141_00003    = fgallag_final_00141_00003;

            I6aa263fc2a061d2c4059b08309f860f4= I0a1e9cf99f1d4725327615f50fcc3ad0 + I675ab6c4fb93b006f3fcafc985fbc405;
            tout_00142_00000    = fgallag_final_00142_00000;

            If3aef2d755013d195fd44f734365d7dc= I0a1e9cf99f1d4725327615f50fcc3ad0 + Ia9c043c5e8873fd13e39cf6bd8136c51;
            tout_00142_00001    = fgallag_final_00142_00001;

            I3ad2e0bbff17683824f575deff82c6bc= I0a1e9cf99f1d4725327615f50fcc3ad0 + I566221060f06e724676ec9bec861d7de;
            tout_00142_00002    = fgallag_final_00142_00002;

            I5087dc4b32d29bfd7bad49026fa58a5d= I0a1e9cf99f1d4725327615f50fcc3ad0 + Ia3cb3ea64576a3e7332e1fb55953aa3e;
            tout_00142_00003    = fgallag_final_00142_00003;

            I8a7d893f3ef6d6a93ba552320d901599= Ie844f4c446983ce381b0bc4c0e8ef7d7 + I082aa8c413d7ef8f054b1c2857cbe39f;
            tout_00143_00000    = fgallag_final_00143_00000;

            Ic057537712e09fa794918e5cde87e084= Ie844f4c446983ce381b0bc4c0e8ef7d7 + Ia0932b3fd6a5ae6da2bacd2b86ba3a43;
            tout_00143_00001    = fgallag_final_00143_00001;

            I0cbab5173052c450504e3a7d15ffda52= Ie844f4c446983ce381b0bc4c0e8ef7d7 + Id682e531735437bc24abbf3d3d51e18b;
            tout_00143_00002    = fgallag_final_00143_00002;

            I81ee40feb7abd0fec3faee653f778f5f= Ie844f4c446983ce381b0bc4c0e8ef7d7 + I3cb1f233951d49f985b0deac6e052bfd;
            tout_00143_00003    = fgallag_final_00143_00003;

            Ia344347a85d4e6afafa2ee3487e65def= I6067f47cccceea96ac46ff0d457b25f2 + If56555b7cf539750706cf678030ccdb2;
            tout_00144_00000    = fgallag_final_00144_00000;

            I038fce1597157a3d95bd9579cc2dcbc6= I6067f47cccceea96ac46ff0d457b25f2 + I097722547450582dc5776bdaff914741;
            tout_00144_00001    = fgallag_final_00144_00001;

            I546585b819c289d855cd098818792e90= I6067f47cccceea96ac46ff0d457b25f2 + I0e2f746715b901feb69f6b3c94f3a828;
            tout_00144_00002    = fgallag_final_00144_00002;

            Ibc3a6609765818327e79519f3e348494= I6067f47cccceea96ac46ff0d457b25f2 + I7015def91103398e54f446ce3e43af01;
            tout_00144_00003    = fgallag_final_00144_00003;

            Id1c71a2a34f9e6239559d28fe2780907= Ifd6fd1f3cbf8884ca7f64bc42278e4fa + I8d0f440df332ea96e2d56eec490fbd51;
            tout_00145_00000    = fgallag_final_00145_00000;

            I1cd6cf5f8119d5e6b4ca40694399b1c2= Ifd6fd1f3cbf8884ca7f64bc42278e4fa + I3bfcd63e92f1949234ab1d2701dbb499;
            tout_00145_00001    = fgallag_final_00145_00001;

            I15e2a1b4356785d73e2ab5d51f1f5ec0= Ifd6fd1f3cbf8884ca7f64bc42278e4fa + Ia8849f78971a45ed0daa2489e7d27dd7;
            tout_00145_00002    = fgallag_final_00145_00002;

            I803aeb29e66384bfc62744a841bcc83e= Ifd6fd1f3cbf8884ca7f64bc42278e4fa + I04874bd1bf257f205b5189c8c20e5a12;
            tout_00145_00003    = fgallag_final_00145_00003;

            Ib6e220dd4f54410239dd0c791d84a700= Iaec9fd9e79371676bfa8ff14b4feae52 + I7cdc5ada6fc68ee31fd4062e2ff004d3;
            tout_00146_00000    = fgallag_final_00146_00000;

            I8a009007fec23f4d492b0da1b6b404fa= Iaec9fd9e79371676bfa8ff14b4feae52 + Ie0622ff815747e4a9f368c74787026ec;
            tout_00146_00001    = fgallag_final_00146_00001;

            I5f89adcb1ba235a74639eca119fb2655= Iaec9fd9e79371676bfa8ff14b4feae52 + I0cf5cb4cd472502b84dbf6fe1af0be78;
            tout_00146_00002    = fgallag_final_00146_00002;

            I8fd2b001ff154e4760ead2df355c80da= Iaec9fd9e79371676bfa8ff14b4feae52 + I937e3a8ede2305ea7c1750283224a870;
            tout_00146_00003    = fgallag_final_00146_00003;

            I581569cc2e63bc68a8466b07ca471b25= I500757c4eda5d3d899aee47b87da585b + I3f0bba472e912f11dea8e788fbc1cb63;
            tout_00147_00000    = fgallag_final_00147_00000;

            Ia9cfdea21a65b0270de42cef7ebbf822= I500757c4eda5d3d899aee47b87da585b + Ie559401a3a913400dc5e3e5641297fa6;
            tout_00147_00001    = fgallag_final_00147_00001;

            Id66a233d2e312aff939549dfa96a8cf0= I500757c4eda5d3d899aee47b87da585b + I4936f823841b0ffe32f801f5134c0211;
            tout_00147_00002    = fgallag_final_00147_00002;

            Ie479c12c25a1964c3804936d45725bdc= I500757c4eda5d3d899aee47b87da585b + Ia7206430a739a11af4d860096eedd6c3;
            tout_00147_00003    = fgallag_final_00147_00003;

            Ie30d8770ab7e6643fcb67463f6999125= I47bf091b0fa74ad511a760bad9d2506c + I72c2256ba47cf03f95143df8f741fd83;
            tout_00148_00000    = fgallag_final_00148_00000;

            I4a17ff532c9341e80f7ed0626f728054= I47bf091b0fa74ad511a760bad9d2506c + I1092325b801600fa7ec85fa640167da9;
            tout_00148_00001    = fgallag_final_00148_00001;

            I597bc1ec224007a78c25f7eea24c2c3e= I47bf091b0fa74ad511a760bad9d2506c + Ibf4c2c00f8e012e9498361bfd3c5b06e;
            tout_00148_00002    = fgallag_final_00148_00002;

            If198ec15fcf66e97e69f88f718979c2b= Ia4c3d0cd9957f678880de5775de76e0d + If26d90629e70c5a871e6f5b14471b8cf;
            tout_00149_00000    = fgallag_final_00149_00000;

            I6aa13ef29cf7e86ec83affca4fa11e42= Ia4c3d0cd9957f678880de5775de76e0d + Iebd050e29044153d5881ef80b2db8c28;
            tout_00149_00001    = fgallag_final_00149_00001;

            Ide136b08f4b6211bca8cccf494a0baa5= Ia4c3d0cd9957f678880de5775de76e0d + I899e5f03cd1d52d11f898959559aaeea;
            tout_00149_00002    = fgallag_final_00149_00002;

            Ieeab247764c23256749776b0a164314d= If5f957fa2f055b1c2c28e8d7cfe3e9ad + I4c03a6569d1b954d088053e38827e811;
            tout_00150_00000    = fgallag_final_00150_00000;

            I210e9ff7f4588185bd712915954543ce= If5f957fa2f055b1c2c28e8d7cfe3e9ad + I0c5250aaca86185fed5978438c8861b6;
            tout_00150_00001    = fgallag_final_00150_00001;

            I59186d5219833d6dd2e813a2910a61f5= If5f957fa2f055b1c2c28e8d7cfe3e9ad + I59c80c7ec26f43308b1a646c47160568;
            tout_00150_00002    = fgallag_final_00150_00002;

            I0c8b2bb61a9c3a67ac7e03e40be2b98e= I3608378a5da8c66bef58528d56192530 + Ibf1c9d86665f696d91c554db748ff42b;
            tout_00151_00000    = fgallag_final_00151_00000;

            Ide24c1f9033e7057262da1bc4762b840= I3608378a5da8c66bef58528d56192530 + I49ccb3e14fe61618806e791ecb4f4eae;
            tout_00151_00001    = fgallag_final_00151_00001;

            I4677558b9faf190e7960cfa9b8ee00fd= I3608378a5da8c66bef58528d56192530 + I8a954a331d36266465a0813d2e8b319b;
            tout_00151_00002    = fgallag_final_00151_00002;

            Ie38ab94215851e531d2100b6602d5fa5= Ie6dead855e00ea0a8e6a9b7503aaebb8 + I239a992ebb62899120a74b1c9e6cc4b4;
            tout_00152_00000    = fgallag_final_00152_00000;

            I3f5119e8fac99376aa38e4765b8b0f99= Ie6dead855e00ea0a8e6a9b7503aaebb8 + I2e802c75c6ce34b05943b678ecbfacb1;
            tout_00152_00001    = fgallag_final_00152_00001;

            Ie8040301d224f78c1fd18bfe9e29e5ba= Ie6dead855e00ea0a8e6a9b7503aaebb8 + I05ecce409cca00ea5b0df25de5a50cf2;
            tout_00152_00002    = fgallag_final_00152_00002;

            Ied989966cebf0d730633606c5182a249= Ie6dead855e00ea0a8e6a9b7503aaebb8 + Ib49e53ca8efd9564ee9572eb3089bb51;
            tout_00152_00003    = fgallag_final_00152_00003;

            Ib8818bc4ca106ae38cacd5c20083aa08= I3bae5e6862e003a8b9a476f72cc6858b + I420e2c5a8745133f6263a71b458f1e2f;
            tout_00153_00000    = fgallag_final_00153_00000;

            Ibf08556fc39044222321912e84a4436b= I3bae5e6862e003a8b9a476f72cc6858b + I9fce6091885f1bb97d29fb1f543b1a38;
            tout_00153_00001    = fgallag_final_00153_00001;

            I985e2740ac0f656da8f9dd973bca99e6= I3bae5e6862e003a8b9a476f72cc6858b + I2de1ca2c390bdd3011fff4a359bb5332;
            tout_00153_00002    = fgallag_final_00153_00002;

            I73012d2d9f6f237bc50bbffc199e012b= I3bae5e6862e003a8b9a476f72cc6858b + Icbde2c6230e9cc67ef12031e38bb344f;
            tout_00153_00003    = fgallag_final_00153_00003;

            Iefd0d59e58623b14437b17297fdbf4ff= I4431adecba8be9e5f21bc6b3e1f8cb10 + Ia47f7fb27f2d965cfd2989569c257356;
            tout_00154_00000    = fgallag_final_00154_00000;

            I68d2443e98f2fd3fa3baf96f98e1f4bc= I4431adecba8be9e5f21bc6b3e1f8cb10 + I034fb3850485fae2d1358041a1c41888;
            tout_00154_00001    = fgallag_final_00154_00001;

            Ia2d1b6833cd8ed02f05281e508e4d716= I4431adecba8be9e5f21bc6b3e1f8cb10 + Id968b34075e351ab01d65abcb4ed8cca;
            tout_00154_00002    = fgallag_final_00154_00002;

            I512e2251bef73108eb0f3e01e79ca3fb= I4431adecba8be9e5f21bc6b3e1f8cb10 + I2e22e867f6f84a7807b82f64a147022e;
            tout_00154_00003    = fgallag_final_00154_00003;

            I9bf64811d14ca8b4c633342ad22669a3= I21c7a2885126d532d00484376588a469 + I174fcbc2ee01fc55edbc8238e5da7f0c;
            tout_00155_00000    = fgallag_final_00155_00000;

            I45a910acd40d5b9417bdfdc50cddf241= I21c7a2885126d532d00484376588a469 + Ia40dad546d9c852e2fa8942c62a1c1f8;
            tout_00155_00001    = fgallag_final_00155_00001;

            Ibbcf5c5f4528b03508b506c43e4511c4= I21c7a2885126d532d00484376588a469 + Icd9a876a0feb16ea62bcad5be2004dac;
            tout_00155_00002    = fgallag_final_00155_00002;

            I2b8b54048e164ef2f1c072517fdfe400= I21c7a2885126d532d00484376588a469 + Id9704e1d8096cd28577c5c357d30b7a4;
            tout_00155_00003    = fgallag_final_00155_00003;

            Ia48d8883fe4f685477da6b4b05ecd387= I2c4d7339ff2fe68d060dd8d961dcab8c + I6dc671e73b4e9c70cabfdeaac2e5c40b;
            tout_00156_00000    = fgallag_final_00156_00000;

            I276395da1f3f1ae246b082408be2cb80= I2c4d7339ff2fe68d060dd8d961dcab8c + Iacf6340a29a5592b61ea875304a2de48;
            tout_00156_00001    = fgallag_final_00156_00001;

            I4d0e2e01d9abf9ce839fe650abfaaddd= I2c4d7339ff2fe68d060dd8d961dcab8c + I487391402b6aa27bf212724a37ea9c33;
            tout_00156_00002    = fgallag_final_00156_00002;

            I7e4e7909094f762c54137cbee99255e5= I2c4d7339ff2fe68d060dd8d961dcab8c + I4b8554cab486a4fc1e14884a6495016e;
            tout_00156_00003    = fgallag_final_00156_00003;

            I761255e100d161b25645ca3a5187e82a= Iee518b15b067eec58cccfa37f7432ea5 + I94e89b3a841f9760e3967c97e86d7160;
            tout_00157_00000    = fgallag_final_00157_00000;

            Icc2ce1fa3cde69256378ec3f4a07b0fc= Iee518b15b067eec58cccfa37f7432ea5 + I5975ef8f6cf53cf2132cdd9d707e7912;
            tout_00157_00001    = fgallag_final_00157_00001;

            Idd99afa80ca23644675d3edd60e74fe4= Iee518b15b067eec58cccfa37f7432ea5 + I6c19936ca2edeb0e261e880a1055e964;
            tout_00157_00002    = fgallag_final_00157_00002;

            I486bcb4fb0af80c98c2ea21ac64f7a90= Iee518b15b067eec58cccfa37f7432ea5 + Iaa235d085a5916a3b0814c3ed2a9026f;
            tout_00157_00003    = fgallag_final_00157_00003;

            I759cca2c0003fc2c2af7709c5ebc59f7= I42145be9c2a80288ba4a2edd91f661a3 + I8d431a0524241fa54cf6dd1e79de4c74;
            tout_00158_00000    = fgallag_final_00158_00000;

            I1d5ce9f132cd1f46e96b511c77234e21= I42145be9c2a80288ba4a2edd91f661a3 + I7b8da162c08f8aa2ae90522ee1526cf6;
            tout_00158_00001    = fgallag_final_00158_00001;

            I032e26ea05e88c6d325a810b67e82306= I42145be9c2a80288ba4a2edd91f661a3 + I7fc190647082a3d71614f46f670167bc;
            tout_00158_00002    = fgallag_final_00158_00002;

            I0f72df5225a1fec2f276fd3c9138e8c3= I42145be9c2a80288ba4a2edd91f661a3 + I5d86ce0b58c0b281d747116a9069ef33;
            tout_00158_00003    = fgallag_final_00158_00003;

            I0d18cf087b2335f1b9e1a621acd5379f= I9dc297ad41fafcda77f5347f331cfc25 + I59547aacdcfde31dc016ec2acbb2f4b4;
            tout_00159_00000    = fgallag_final_00159_00000;

            I7684fc23c57105e856050a45640f2bfd= I9dc297ad41fafcda77f5347f331cfc25 + Ie4749f8e9ad2b370f9f9814b5a463c43;
            tout_00159_00001    = fgallag_final_00159_00001;

            If778767ab80e59e940deeaa8a0dac99a= I9dc297ad41fafcda77f5347f331cfc25 + I495f8be463b15db906474c518e0741e2;
            tout_00159_00002    = fgallag_final_00159_00002;

            Idaf86833beb8c334f99291db9302ed29= I9dc297ad41fafcda77f5347f331cfc25 + Id20394136fb036435bb4680aac64581f;
            tout_00159_00003    = fgallag_final_00159_00003;

            I6610e8d41cea10498d95850440ce388b= I846700c79f30ca954cc2933fc94d355b + I5ffed139764d90825b9f2eddacd0eddc;
            tout_00160_00000    = fgallag_final_00160_00000;

            Ibc653e701eb995e828c8180efaa122c9= I846700c79f30ca954cc2933fc94d355b + I733c3fa4d84e5680792b16a70bb1a51d;
            tout_00160_00001    = fgallag_final_00160_00001;

            I21d36c49c9c766139b4b01df7c00a8f3= I846700c79f30ca954cc2933fc94d355b + I3c057d64cf4fca0238a874f0ced99c76;
            tout_00160_00002    = fgallag_final_00160_00002;

            I0e4ffded936d7ccfc32b410aec617df8= I846700c79f30ca954cc2933fc94d355b + I8a16afac6e470ca69634d7fe9656387a;
            tout_00160_00003    = fgallag_final_00160_00003;

            I1a5745021323efb5327d0b893962e852= I8af96a91457316e49e3f7dd5e57c82da + Ie0667fbe76244eaec0b155d69dcc9447;
            tout_00161_00000    = fgallag_final_00161_00000;

            I65547afdcd7fedb7b44bd51358eec4d2= I8af96a91457316e49e3f7dd5e57c82da + Iedb9bb14951bf67bc8865b0983490c14;
            tout_00161_00001    = fgallag_final_00161_00001;

            Iada3eb71e94ff6a6f4e5c702e83036ed= I8af96a91457316e49e3f7dd5e57c82da + Ic78949e07e643f571f23df7e8f15d9fb;
            tout_00161_00002    = fgallag_final_00161_00002;

            I077404a911da16d707a326f18717dc7a= I8af96a91457316e49e3f7dd5e57c82da + Ic4e7f690bc050f1d1f84eae7ca193e1c;
            tout_00161_00003    = fgallag_final_00161_00003;

            I6da1e92759c96aab8b9207a9acb244ab= I7d1c247500d7d32e406b2a5f7e2b745b + Id4a213e494f9c9be0fd1a307e87c756a;
            tout_00162_00000    = fgallag_final_00162_00000;

            If7110182720ffa279b1cec1305cf9889= I7d1c247500d7d32e406b2a5f7e2b745b + Idda26504e422367082caeafbb29871f9;
            tout_00162_00001    = fgallag_final_00162_00001;

            If0e20ea1696ff84329b9928d7f9e3381= I7d1c247500d7d32e406b2a5f7e2b745b + I461ebbf3a02ae63e2eb27531b1370f24;
            tout_00162_00002    = fgallag_final_00162_00002;

            I4e69ae6e73a856d4e26203fb9acf3565= I7d1c247500d7d32e406b2a5f7e2b745b + Ia60421aa427236540b4d0d08d52ff507;
            tout_00162_00003    = fgallag_final_00162_00003;

            I64c939aa568669b4567c21be09ad0e94= I66d85c030a8864505298919046056305 + I5e2331edf6e881e9f3a8c47eebda0ac4;
            tout_00163_00000    = fgallag_final_00163_00000;

            Ia88eb16f68265e322509d541eb457993= I66d85c030a8864505298919046056305 + Ieb0336a1974a2aec0966f4f59f460802;
            tout_00163_00001    = fgallag_final_00163_00001;

            I916f75e5a3858a420ab5cd4c43b13921= I66d85c030a8864505298919046056305 + Ib028686da9c849e827cf249a744b7db3;
            tout_00163_00002    = fgallag_final_00163_00002;

            Id076f99460a8f73a9fd43467216e8f8e= I66d85c030a8864505298919046056305 + Icace650ee3865bd7bbddd2d9435c5561;
            tout_00163_00003    = fgallag_final_00163_00003;

            Ib4d7aeb8544fbdc36575a55b9f67f2dc= I4841257ae596d9d3e4eb1e6f886956b0 + If2b17f9e9186542117f43d0dd342326e;
            tout_00164_00000    = fgallag_final_00164_00000;

            If65d2514892fb7ee64fa4dc37fc0fed3= I4841257ae596d9d3e4eb1e6f886956b0 + I0b0dd019d8bd24684403a29aed668b6d;
            tout_00164_00001    = fgallag_final_00164_00001;

            Ibef07e48768252e9b41baf067bb1ff5d= I4841257ae596d9d3e4eb1e6f886956b0 + I831d214dcb4f8d534b5ddaaeaeeb81ce;
            tout_00164_00002    = fgallag_final_00164_00002;

            Ib8fb61fa9cb8e92bc57c53a567891895= I4841257ae596d9d3e4eb1e6f886956b0 + I7d27d070b96b7810f667e1d1845342d3;
            tout_00164_00003    = fgallag_final_00164_00003;

            Id8f5f32cd0757b4d6861d17fcbd6e8d0= Icd6f7ec117f9ab4eda8c5eba41386ffa + Id4dc304aef5f35f6ceb91796c278e716;
            tout_00165_00000    = fgallag_final_00165_00000;

            I8be241f29e7eb258e9b3501430820b0d= Icd6f7ec117f9ab4eda8c5eba41386ffa + Ieb3f28762410fb40a0c8a8556b4b3ca0;
            tout_00165_00001    = fgallag_final_00165_00001;

            Ica8a188ea43e2f28e70b8ea4e2431dc3= Icd6f7ec117f9ab4eda8c5eba41386ffa + I6fb55222b69475b7168874423226ec9c;
            tout_00165_00002    = fgallag_final_00165_00002;

            I83ceb726e57d52698b57dc39ce585897= Icd6f7ec117f9ab4eda8c5eba41386ffa + Ida7ec09c913caa0e78a2c4cbaae517c8;
            tout_00165_00003    = fgallag_final_00165_00003;

            Ic88e7e05d83ff800b4a941ae4b424557= Ibc0498839d1d9b6dc853b8e5d7a88fa3 + I927c870d09285dcb47e6d399f319471e;
            tout_00166_00000    = fgallag_final_00166_00000;

            I7de81aaac1e5776dfb60eed2d12d4f6d= Ibc0498839d1d9b6dc853b8e5d7a88fa3 + Ib402cdbfaa9900820b85bd625415c547;
            tout_00166_00001    = fgallag_final_00166_00001;

            I37058036bd9f4331387ee4a9348541e2= Ibc0498839d1d9b6dc853b8e5d7a88fa3 + I84da4ce7441e132e775167c1cd81dbe5;
            tout_00166_00002    = fgallag_final_00166_00002;

            I570f85838c418d8501c8ccdc38a53f00= Ibc0498839d1d9b6dc853b8e5d7a88fa3 + Ic5eba898858be1f768841ead792d6d86;
            tout_00166_00003    = fgallag_final_00166_00003;

            I4aa6f0c0f5163b944f11328888af73e0= I142ebca7f155e287e38ddf45423ab0fd + I4b8d520ee88fd39d83a16432e962f731;
            tout_00167_00000    = fgallag_final_00167_00000;

            Ic7fc1f38ad4e9b2cb472ae75bc3c100c= I142ebca7f155e287e38ddf45423ab0fd + I0e7079db66c15210046b997f319ece89;
            tout_00167_00001    = fgallag_final_00167_00001;

            Ibace8d2fba25834c83b1e57195c81086= I142ebca7f155e287e38ddf45423ab0fd + I8f8273c4cb2a9ace8a09847efd4bdec7;
            tout_00167_00002    = fgallag_final_00167_00002;

            Iefc1488e3eb60b99ae08d904a15c5242= I142ebca7f155e287e38ddf45423ab0fd + I72197797a307c611fa8952533e63d7bf;
            tout_00167_00003    = fgallag_final_00167_00003;
end

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
              Ifc045af19c3f10d92d2b0dfb4fbbde38 <= {(HAM_LEN){1'b0}};
       end else begin
           if (start_d8) begin
              if (Ib325dab091dfc3a1a269adb3ea9c75cd <= HamDist_sum_mm) begin
                  Ifc045af19c3f10d92d2b0dfb4fbbde38 <= Ifc045af19c3f10d92d2b0dfb4fbbde38 + 1;
              end
           end
           else if (start_dec) begin
                  Ifc045af19c3f10d92d2b0dfb4fbbde38 <= {(HAM_LEN){1'b0}};
           end
       end
   end

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
                 HamDist_iir <= 'h0;
       end else begin
          if (start_d8) begin
             if (HamDist_loop == 0)
                 HamDist_iir <= HamDist_sum_mm;
             else
                 HamDist_iir <= HamDist_iir_prod;
          end
       end
   end

   always_comb HamDist_iir_prod = ((HamDist_iir * HamDist_iir1 + HamDist_sum_mm *HamDist_iir2 + HamDist_iir3));



   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
                 Ib325dab091dfc3a1a269adb3ea9c75cd <= {(HAM_LEN){1'b0}};
       end else begin
          if (start_d8) begin
             if (HamDist_loop == 0)
                 Ib325dab091dfc3a1a269adb3ea9c75cd <= {(HAM_LEN){1'b0}};
             else
                 Ib325dab091dfc3a1a269adb3ea9c75cd <= HamDist_sum_mm;
          end
       end
   end





   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
          converged_loops_ended <= 1'b0;
          converged_pass_fail <= 1'b0;
       end else begin
          if (start_dec) begin
               converged_loops_ended <= 1'b0;
               converged_pass_fail <= 1'b0;
          end else begin
               if (start_d9) begin
                       if (
                         (HamDist_sum_mm*100 > HamDist_iir * HamDist_loop_percentage) ||
                         (Ifc045af19c3f10d92d2b0dfb4fbbde38 > HamDist_loop_max)
                         ) begin
                         converged_loops_ended <= 1'b1;
                         converged_pass_fail <= 1'b0;
                       end else if (HamDist_sum_mm == 0) begin
                         converged_loops_ended <= 1'b1;
                         converged_pass_fail <= 1'b1;
                       end

               end  //start_d8
               else begin // else I8bf8854bebe108183caeb845c7676ae4 start_d8
                    //wait for the start_dec to clear I0d149b90e7394297301c90191ae775f0 I3262d48df5d75e3452f0f16b313b7808
                    //converged_loops_ended <= 1'b0;
                    //converged_pass_fail <= 1'b0;
               end


          end  //start_dec
       end  //rstn
   end

//tmp_bit valid Ied2b5c0139cec8ad2873829dc1117d50 start_d7
// I7fa3b767c460b54a2be4d49030b349c7 cycle I7243f8be75253afbadf7477867021f8b I13b5bfe96f3e2fe411c9f66f4a582adf I724a00e315992b82d662231ea0dcbe50 or I190ebdd6b6c2b422296a6ee2cce59699 I0aa6f4210bf373c95eda00232e93cd98
always_comb HamDist_cntr_inc_converged_valid = start_d6;

assign tmp_bit_0 = sum0_00000[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[0] = tmp_bit_0;
assign tmp_bit_1 = sum0_00001[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[1] = tmp_bit_1;
assign tmp_bit_2 = sum0_00002[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[2] = tmp_bit_2;
assign tmp_bit_3 = sum0_00003[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[3] = tmp_bit_3;
assign tmp_bit_4 = sum0_00004[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[4] = tmp_bit_4;
assign tmp_bit_5 = sum0_00005[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[5] = tmp_bit_5;
assign tmp_bit_6 = sum0_00006[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[6] = tmp_bit_6;
assign tmp_bit_7 = sum0_00007[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[7] = tmp_bit_7;
assign tmp_bit_8 = sum0_00008[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[8] = tmp_bit_8;
assign tmp_bit_9 = sum0_00009[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[9] = tmp_bit_9;
assign tmp_bit_10 = sum0_00010[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[10] = tmp_bit_10;
assign tmp_bit_11 = sum0_00011[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[11] = tmp_bit_11;
assign tmp_bit_12 = sum0_00012[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[12] = tmp_bit_12;
assign tmp_bit_13 = sum0_00013[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[13] = tmp_bit_13;
assign tmp_bit_14 = sum0_00014[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[14] = tmp_bit_14;
assign tmp_bit_15 = sum0_00015[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[15] = tmp_bit_15;
assign tmp_bit_16 = sum0_00016[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[16] = tmp_bit_16;
assign tmp_bit_17 = sum0_00017[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[17] = tmp_bit_17;
assign tmp_bit_18 = sum0_00018[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[18] = tmp_bit_18;
assign tmp_bit_19 = sum0_00019[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[19] = tmp_bit_19;
assign tmp_bit_20 = sum0_00020[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[20] = tmp_bit_20;
assign tmp_bit_21 = sum0_00021[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[21] = tmp_bit_21;
assign tmp_bit_22 = sum0_00022[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[22] = tmp_bit_22;
assign tmp_bit_23 = sum0_00023[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[23] = tmp_bit_23;
assign tmp_bit_24 = sum0_00024[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[24] = tmp_bit_24;
assign tmp_bit_25 = sum0_00025[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[25] = tmp_bit_25;
assign tmp_bit_26 = sum0_00026[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[26] = tmp_bit_26;
assign tmp_bit_27 = sum0_00027[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[27] = tmp_bit_27;
assign tmp_bit_28 = sum0_00028[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[28] = tmp_bit_28;
assign tmp_bit_29 = sum0_00029[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[29] = tmp_bit_29;
assign tmp_bit_30 = sum0_00030[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[30] = tmp_bit_30;
assign tmp_bit_31 = sum0_00031[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[31] = tmp_bit_31;
assign tmp_bit_32 = sum0_00032[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[32] = tmp_bit_32;
assign tmp_bit_33 = sum0_00033[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[33] = tmp_bit_33;
assign tmp_bit_34 = sum0_00034[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[34] = tmp_bit_34;
assign tmp_bit_35 = sum0_00035[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[35] = tmp_bit_35;
assign tmp_bit_36 = sum0_00036[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[36] = tmp_bit_36;
assign tmp_bit_37 = sum0_00037[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[37] = tmp_bit_37;
assign tmp_bit_38 = sum0_00038[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[38] = tmp_bit_38;
assign tmp_bit_39 = sum0_00039[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[39] = tmp_bit_39;
assign tmp_bit_40 = sum0_00040[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[40] = tmp_bit_40;
assign tmp_bit_41 = sum0_00041[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[41] = tmp_bit_41;
assign tmp_bit_42 = sum0_00042[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[42] = tmp_bit_42;
assign tmp_bit_43 = sum0_00043[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[43] = tmp_bit_43;
assign tmp_bit_44 = sum0_00044[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[44] = tmp_bit_44;
assign tmp_bit_45 = sum0_00045[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[45] = tmp_bit_45;
assign tmp_bit_46 = sum0_00046[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[46] = tmp_bit_46;
assign tmp_bit_47 = sum0_00047[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[47] = tmp_bit_47;
assign tmp_bit_48 = sum0_00048[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[48] = tmp_bit_48;
assign tmp_bit_49 = sum0_00049[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[49] = tmp_bit_49;
assign tmp_bit_50 = sum0_00050[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[50] = tmp_bit_50;
assign tmp_bit_51 = sum0_00051[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[51] = tmp_bit_51;
assign tmp_bit_52 = sum0_00052[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[52] = tmp_bit_52;
assign tmp_bit_53 = sum0_00053[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[53] = tmp_bit_53;
assign tmp_bit_54 = sum0_00054[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[54] = tmp_bit_54;
assign tmp_bit_55 = sum0_00055[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[55] = tmp_bit_55;
assign tmp_bit_56 = sum0_00056[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[56] = tmp_bit_56;
assign tmp_bit_57 = sum0_00057[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[57] = tmp_bit_57;
assign tmp_bit_58 = sum0_00058[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[58] = tmp_bit_58;
assign tmp_bit_59 = sum0_00059[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[59] = tmp_bit_59;
assign tmp_bit_60 = sum0_00060[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[60] = tmp_bit_60;
assign tmp_bit_61 = sum0_00061[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[61] = tmp_bit_61;
assign tmp_bit_62 = sum0_00062[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[62] = tmp_bit_62;
assign tmp_bit_63 = sum0_00063[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[63] = tmp_bit_63;
assign tmp_bit_64 = sum0_00064[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[64] = tmp_bit_64;
assign tmp_bit_65 = sum0_00065[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[65] = tmp_bit_65;
assign tmp_bit_66 = sum0_00066[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[66] = tmp_bit_66;
assign tmp_bit_67 = sum0_00067[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[67] = tmp_bit_67;
assign tmp_bit_68 = sum0_00068[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[68] = tmp_bit_68;
assign tmp_bit_69 = sum0_00069[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[69] = tmp_bit_69;
assign tmp_bit_70 = sum0_00070[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[70] = tmp_bit_70;
assign tmp_bit_71 = sum0_00071[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[71] = tmp_bit_71;
assign tmp_bit_72 = sum0_00072[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[72] = tmp_bit_72;
assign tmp_bit_73 = sum0_00073[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[73] = tmp_bit_73;
assign tmp_bit_74 = sum0_00074[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[74] = tmp_bit_74;
assign tmp_bit_75 = sum0_00075[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[75] = tmp_bit_75;
assign tmp_bit_76 = sum0_00076[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[76] = tmp_bit_76;
assign tmp_bit_77 = sum0_00077[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[77] = tmp_bit_77;
assign tmp_bit_78 = sum0_00078[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[78] = tmp_bit_78;
assign tmp_bit_79 = sum0_00079[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[79] = tmp_bit_79;
assign tmp_bit_80 = sum0_00080[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[80] = tmp_bit_80;
assign tmp_bit_81 = sum0_00081[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[81] = tmp_bit_81;
assign tmp_bit_82 = sum0_00082[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[82] = tmp_bit_82;
assign tmp_bit_83 = sum0_00083[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[83] = tmp_bit_83;
assign tmp_bit_84 = sum0_00084[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[84] = tmp_bit_84;
assign tmp_bit_85 = sum0_00085[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[85] = tmp_bit_85;
assign tmp_bit_86 = sum0_00086[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[86] = tmp_bit_86;
assign tmp_bit_87 = sum0_00087[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[87] = tmp_bit_87;
assign tmp_bit_88 = sum0_00088[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[88] = tmp_bit_88;
assign tmp_bit_89 = sum0_00089[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[89] = tmp_bit_89;
assign tmp_bit_90 = sum0_00090[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[90] = tmp_bit_90;
assign tmp_bit_91 = sum0_00091[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[91] = tmp_bit_91;
assign tmp_bit_92 = sum0_00092[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[92] = tmp_bit_92;
assign tmp_bit_93 = sum0_00093[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[93] = tmp_bit_93;
assign tmp_bit_94 = sum0_00094[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[94] = tmp_bit_94;
assign tmp_bit_95 = sum0_00095[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[95] = tmp_bit_95;
assign tmp_bit_96 = sum0_00096[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[96] = tmp_bit_96;
assign tmp_bit_97 = sum0_00097[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[97] = tmp_bit_97;
assign tmp_bit_98 = sum0_00098[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[98] = tmp_bit_98;
assign tmp_bit_99 = sum0_00099[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[99] = tmp_bit_99;
assign tmp_bit_100 = sum0_00100[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[100] = tmp_bit_100;
assign tmp_bit_101 = sum0_00101[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[101] = tmp_bit_101;
assign tmp_bit_102 = sum0_00102[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[102] = tmp_bit_102;
assign tmp_bit_103 = sum0_00103[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[103] = tmp_bit_103;
assign tmp_bit_104 = sum0_00104[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[104] = tmp_bit_104;
assign tmp_bit_105 = sum0_00105[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[105] = tmp_bit_105;
assign tmp_bit_106 = sum0_00106[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[106] = tmp_bit_106;
assign tmp_bit_107 = sum0_00107[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[107] = tmp_bit_107;
assign tmp_bit_108 = sum0_00108[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[108] = tmp_bit_108;
assign tmp_bit_109 = sum0_00109[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[109] = tmp_bit_109;
assign tmp_bit_110 = sum0_00110[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[110] = tmp_bit_110;
assign tmp_bit_111 = sum0_00111[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[111] = tmp_bit_111;
assign tmp_bit_112 = sum0_00112[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[112] = tmp_bit_112;
assign tmp_bit_113 = sum0_00113[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[113] = tmp_bit_113;
assign tmp_bit_114 = sum0_00114[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[114] = tmp_bit_114;
assign tmp_bit_115 = sum0_00115[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[115] = tmp_bit_115;
assign tmp_bit_116 = sum0_00116[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[116] = tmp_bit_116;
assign tmp_bit_117 = sum0_00117[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[117] = tmp_bit_117;
assign tmp_bit_118 = sum0_00118[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[118] = tmp_bit_118;
assign tmp_bit_119 = sum0_00119[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[119] = tmp_bit_119;
assign tmp_bit_120 = sum0_00120[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[120] = tmp_bit_120;
assign tmp_bit_121 = sum0_00121[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[121] = tmp_bit_121;
assign tmp_bit_122 = sum0_00122[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[122] = tmp_bit_122;
assign tmp_bit_123 = sum0_00123[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[123] = tmp_bit_123;
assign tmp_bit_124 = sum0_00124[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[124] = tmp_bit_124;
assign tmp_bit_125 = sum0_00125[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[125] = tmp_bit_125;
assign tmp_bit_126 = sum0_00126[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[126] = tmp_bit_126;
assign tmp_bit_127 = sum0_00127[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[127] = tmp_bit_127;
assign tmp_bit_128 = sum0_00128[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[128] = tmp_bit_128;
assign tmp_bit_129 = sum0_00129[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[129] = tmp_bit_129;
assign tmp_bit_130 = sum0_00130[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[130] = tmp_bit_130;
assign tmp_bit_131 = sum0_00131[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[131] = tmp_bit_131;
assign tmp_bit_132 = sum0_00132[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[132] = tmp_bit_132;
assign tmp_bit_133 = sum0_00133[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[133] = tmp_bit_133;
assign tmp_bit_134 = sum0_00134[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[134] = tmp_bit_134;
assign tmp_bit_135 = sum0_00135[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[135] = tmp_bit_135;
assign tmp_bit_136 = sum0_00136[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[136] = tmp_bit_136;
assign tmp_bit_137 = sum0_00137[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[137] = tmp_bit_137;
assign tmp_bit_138 = sum0_00138[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[138] = tmp_bit_138;
assign tmp_bit_139 = sum0_00139[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[139] = tmp_bit_139;
assign tmp_bit_140 = sum0_00140[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[140] = tmp_bit_140;
assign tmp_bit_141 = sum0_00141[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[141] = tmp_bit_141;
assign tmp_bit_142 = sum0_00142[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[142] = tmp_bit_142;
assign tmp_bit_143 = sum0_00143[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[143] = tmp_bit_143;
assign tmp_bit_144 = sum0_00144[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[144] = tmp_bit_144;
assign tmp_bit_145 = sum0_00145[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[145] = tmp_bit_145;
assign tmp_bit_146 = sum0_00146[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[146] = tmp_bit_146;
assign tmp_bit_147 = sum0_00147[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[147] = tmp_bit_147;
assign tmp_bit_148 = sum0_00148[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[148] = tmp_bit_148;
assign tmp_bit_149 = sum0_00149[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[149] = tmp_bit_149;
assign tmp_bit_150 = sum0_00150[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[150] = tmp_bit_150;
assign tmp_bit_151 = sum0_00151[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[151] = tmp_bit_151;
assign tmp_bit_152 = sum0_00152[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[152] = tmp_bit_152;
assign tmp_bit_153 = sum0_00153[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[153] = tmp_bit_153;
assign tmp_bit_154 = sum0_00154[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[154] = tmp_bit_154;
assign tmp_bit_155 = sum0_00155[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[155] = tmp_bit_155;
assign tmp_bit_156 = sum0_00156[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[156] = tmp_bit_156;
assign tmp_bit_157 = sum0_00157[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[157] = tmp_bit_157;
assign tmp_bit_158 = sum0_00158[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[158] = tmp_bit_158;
assign tmp_bit_159 = sum0_00159[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[159] = tmp_bit_159;
assign tmp_bit_160 = sum0_00160[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[160] = tmp_bit_160;
assign tmp_bit_161 = sum0_00161[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[161] = tmp_bit_161;
assign tmp_bit_162 = sum0_00162[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[162] = tmp_bit_162;
assign tmp_bit_163 = sum0_00163[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[163] = tmp_bit_163;
assign tmp_bit_164 = sum0_00164[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[164] = tmp_bit_164;
assign tmp_bit_165 = sum0_00165[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[165] = tmp_bit_165;
assign tmp_bit_166 = sum0_00166[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[166] = tmp_bit_166;
assign tmp_bit_167 = sum0_00167[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[167] = tmp_bit_167;
assign tmp_bit_168 = sum0_00168[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[168] = tmp_bit_168;
assign tmp_bit_169 = sum0_00169[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[169] = tmp_bit_169;
assign tmp_bit_170 = sum0_00170[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[170] = tmp_bit_170;
assign tmp_bit_171 = sum0_00171[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[171] = tmp_bit_171;
assign tmp_bit_172 = sum0_00172[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[172] = tmp_bit_172;
assign tmp_bit_173 = sum0_00173[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[173] = tmp_bit_173;
assign tmp_bit_174 = sum0_00174[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[174] = tmp_bit_174;
assign tmp_bit_175 = sum0_00175[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[175] = tmp_bit_175;
assign tmp_bit_176 = sum0_00176[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[176] = tmp_bit_176;
assign tmp_bit_177 = sum0_00177[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[177] = tmp_bit_177;
assign tmp_bit_178 = sum0_00178[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[178] = tmp_bit_178;
assign tmp_bit_179 = sum0_00179[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[179] = tmp_bit_179;
assign tmp_bit_180 = sum0_00180[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[180] = tmp_bit_180;
assign tmp_bit_181 = sum0_00181[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[181] = tmp_bit_181;
assign tmp_bit_182 = sum0_00182[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[182] = tmp_bit_182;
assign tmp_bit_183 = sum0_00183[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[183] = tmp_bit_183;
assign tmp_bit_184 = sum0_00184[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[184] = tmp_bit_184;
assign tmp_bit_185 = sum0_00185[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[185] = tmp_bit_185;
assign tmp_bit_186 = sum0_00186[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[186] = tmp_bit_186;
assign tmp_bit_187 = sum0_00187[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[187] = tmp_bit_187;
assign tmp_bit_188 = sum0_00188[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[188] = tmp_bit_188;
assign tmp_bit_189 = sum0_00189[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[189] = tmp_bit_189;
assign tmp_bit_190 = sum0_00190[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[190] = tmp_bit_190;
assign tmp_bit_191 = sum0_00191[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[191] = tmp_bit_191;
assign tmp_bit_192 = sum0_00192[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[192] = tmp_bit_192;
assign tmp_bit_193 = sum0_00193[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[193] = tmp_bit_193;
assign tmp_bit_194 = sum0_00194[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[194] = tmp_bit_194;
assign tmp_bit_195 = sum0_00195[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[195] = tmp_bit_195;
assign tmp_bit_196 = sum0_00196[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[196] = tmp_bit_196;
assign tmp_bit_197 = sum0_00197[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[197] = tmp_bit_197;
assign tmp_bit_198 = sum0_00198[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[198] = tmp_bit_198;
assign tmp_bit_199 = sum0_00199[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[199] = tmp_bit_199;
assign tmp_bit_200 = sum0_00200[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[200] = tmp_bit_200;
assign tmp_bit_201 = sum0_00201[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[201] = tmp_bit_201;
assign tmp_bit_202 = sum0_00202[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[202] = tmp_bit_202;
assign tmp_bit_203 = sum0_00203[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[203] = tmp_bit_203;
assign tmp_bit_204 = sum0_00204[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[204] = tmp_bit_204;
assign tmp_bit_205 = sum0_00205[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[205] = tmp_bit_205;
assign tmp_bit_206 = sum0_00206[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[206] = tmp_bit_206;
assign tmp_bit_207 = sum0_00207[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[207] = tmp_bit_207;

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin

// Ie4894ca167b08880bfc35862f18575eb Ied2b5c0139cec8ad2873829dc1117d50 clock start_d7 valid Ied2b5c0139cec8ad2873829dc1117d50 start_d7
          tmp_bit[0]  <=   0;
          tmp_bit[1]  <=   0;
          tmp_bit[2]  <=   0;
          tmp_bit[3]  <=   0;
          tmp_bit[4]  <=   0;
          tmp_bit[5]  <=   0;
          tmp_bit[6]  <=   0;
          tmp_bit[7]  <=   0;
          tmp_bit[8]  <=   0;
          tmp_bit[9]  <=   0;
          tmp_bit[10]  <=   0;
          tmp_bit[11]  <=   0;
          tmp_bit[12]  <=   0;
          tmp_bit[13]  <=   0;
          tmp_bit[14]  <=   0;
          tmp_bit[15]  <=   0;
          tmp_bit[16]  <=   0;
          tmp_bit[17]  <=   0;
          tmp_bit[18]  <=   0;
          tmp_bit[19]  <=   0;
          tmp_bit[20]  <=   0;
          tmp_bit[21]  <=   0;
          tmp_bit[22]  <=   0;
          tmp_bit[23]  <=   0;
          tmp_bit[24]  <=   0;
          tmp_bit[25]  <=   0;
          tmp_bit[26]  <=   0;
          tmp_bit[27]  <=   0;
          tmp_bit[28]  <=   0;
          tmp_bit[29]  <=   0;
          tmp_bit[30]  <=   0;
          tmp_bit[31]  <=   0;
          tmp_bit[32]  <=   0;
          tmp_bit[33]  <=   0;
          tmp_bit[34]  <=   0;
          tmp_bit[35]  <=   0;
          tmp_bit[36]  <=   0;
          tmp_bit[37]  <=   0;
          tmp_bit[38]  <=   0;
          tmp_bit[39]  <=   0;
          tmp_bit[40]  <=   0;
          tmp_bit[41]  <=   0;
          tmp_bit[42]  <=   0;
          tmp_bit[43]  <=   0;
          tmp_bit[44]  <=   0;
          tmp_bit[45]  <=   0;
          tmp_bit[46]  <=   0;
          tmp_bit[47]  <=   0;
          tmp_bit[48]  <=   0;
          tmp_bit[49]  <=   0;
          tmp_bit[50]  <=   0;
          tmp_bit[51]  <=   0;
          tmp_bit[52]  <=   0;
          tmp_bit[53]  <=   0;
          tmp_bit[54]  <=   0;
          tmp_bit[55]  <=   0;
          tmp_bit[56]  <=   0;
          tmp_bit[57]  <=   0;
          tmp_bit[58]  <=   0;
          tmp_bit[59]  <=   0;
          tmp_bit[60]  <=   0;
          tmp_bit[61]  <=   0;
          tmp_bit[62]  <=   0;
          tmp_bit[63]  <=   0;
          tmp_bit[64]  <=   0;
          tmp_bit[65]  <=   0;
          tmp_bit[66]  <=   0;
          tmp_bit[67]  <=   0;
          tmp_bit[68]  <=   0;
          tmp_bit[69]  <=   0;
          tmp_bit[70]  <=   0;
          tmp_bit[71]  <=   0;
          tmp_bit[72]  <=   0;
          tmp_bit[73]  <=   0;
          tmp_bit[74]  <=   0;
          tmp_bit[75]  <=   0;
          tmp_bit[76]  <=   0;
          tmp_bit[77]  <=   0;
          tmp_bit[78]  <=   0;
          tmp_bit[79]  <=   0;
          tmp_bit[80]  <=   0;
          tmp_bit[81]  <=   0;
          tmp_bit[82]  <=   0;
          tmp_bit[83]  <=   0;
          tmp_bit[84]  <=   0;
          tmp_bit[85]  <=   0;
          tmp_bit[86]  <=   0;
          tmp_bit[87]  <=   0;
          tmp_bit[88]  <=   0;
          tmp_bit[89]  <=   0;
          tmp_bit[90]  <=   0;
          tmp_bit[91]  <=   0;
          tmp_bit[92]  <=   0;
          tmp_bit[93]  <=   0;
          tmp_bit[94]  <=   0;
          tmp_bit[95]  <=   0;
          tmp_bit[96]  <=   0;
          tmp_bit[97]  <=   0;
          tmp_bit[98]  <=   0;
          tmp_bit[99]  <=   0;
          tmp_bit[100]  <=   0;
          tmp_bit[101]  <=   0;
          tmp_bit[102]  <=   0;
          tmp_bit[103]  <=   0;
          tmp_bit[104]  <=   0;
          tmp_bit[105]  <=   0;
          tmp_bit[106]  <=   0;
          tmp_bit[107]  <=   0;
          tmp_bit[108]  <=   0;
          tmp_bit[109]  <=   0;
          tmp_bit[110]  <=   0;
          tmp_bit[111]  <=   0;
          tmp_bit[112]  <=   0;
          tmp_bit[113]  <=   0;
          tmp_bit[114]  <=   0;
          tmp_bit[115]  <=   0;
          tmp_bit[116]  <=   0;
          tmp_bit[117]  <=   0;
          tmp_bit[118]  <=   0;
          tmp_bit[119]  <=   0;
          tmp_bit[120]  <=   0;
          tmp_bit[121]  <=   0;
          tmp_bit[122]  <=   0;
          tmp_bit[123]  <=   0;
          tmp_bit[124]  <=   0;
          tmp_bit[125]  <=   0;
          tmp_bit[126]  <=   0;
          tmp_bit[127]  <=   0;
          tmp_bit[128]  <=   0;
          tmp_bit[129]  <=   0;
          tmp_bit[130]  <=   0;
          tmp_bit[131]  <=   0;
          tmp_bit[132]  <=   0;
          tmp_bit[133]  <=   0;
          tmp_bit[134]  <=   0;
          tmp_bit[135]  <=   0;
          tmp_bit[136]  <=   0;
          tmp_bit[137]  <=   0;
          tmp_bit[138]  <=   0;
          tmp_bit[139]  <=   0;
          tmp_bit[140]  <=   0;
          tmp_bit[141]  <=   0;
          tmp_bit[142]  <=   0;
          tmp_bit[143]  <=   0;
          tmp_bit[144]  <=   0;
          tmp_bit[145]  <=   0;
          tmp_bit[146]  <=   0;
          tmp_bit[147]  <=   0;
          tmp_bit[148]  <=   0;
          tmp_bit[149]  <=   0;
          tmp_bit[150]  <=   0;
          tmp_bit[151]  <=   0;
          tmp_bit[152]  <=   0;
          tmp_bit[153]  <=   0;
          tmp_bit[154]  <=   0;
          tmp_bit[155]  <=   0;
          tmp_bit[156]  <=   0;
          tmp_bit[157]  <=   0;
          tmp_bit[158]  <=   0;
          tmp_bit[159]  <=   0;
          tmp_bit[160]  <=   0;
          tmp_bit[161]  <=   0;
          tmp_bit[162]  <=   0;
          tmp_bit[163]  <=   0;
          tmp_bit[164]  <=   0;
          tmp_bit[165]  <=   0;
          tmp_bit[166]  <=   0;
          tmp_bit[167]  <=   0;
          tmp_bit[168]  <=   0;
          tmp_bit[169]  <=   0;
          tmp_bit[170]  <=   0;
          tmp_bit[171]  <=   0;
          tmp_bit[172]  <=   0;
          tmp_bit[173]  <=   0;
          tmp_bit[174]  <=   0;
          tmp_bit[175]  <=   0;
          tmp_bit[176]  <=   0;
          tmp_bit[177]  <=   0;
          tmp_bit[178]  <=   0;
          tmp_bit[179]  <=   0;
          tmp_bit[180]  <=   0;
          tmp_bit[181]  <=   0;
          tmp_bit[182]  <=   0;
          tmp_bit[183]  <=   0;
          tmp_bit[184]  <=   0;
          tmp_bit[185]  <=   0;
          tmp_bit[186]  <=   0;
          tmp_bit[187]  <=   0;
          tmp_bit[188]  <=   0;
          tmp_bit[189]  <=   0;
          tmp_bit[190]  <=   0;
          tmp_bit[191]  <=   0;
          tmp_bit[192]  <=   0;
          tmp_bit[193]  <=   0;
          tmp_bit[194]  <=   0;
          tmp_bit[195]  <=   0;
          tmp_bit[196]  <=   0;
          tmp_bit[197]  <=   0;
          tmp_bit[198]  <=   0;
          tmp_bit[199]  <=   0;
          tmp_bit[200]  <=   0;
          tmp_bit[201]  <=   0;
          tmp_bit[202]  <=   0;
          tmp_bit[203]  <=   0;
          tmp_bit[204]  <=   0;
          tmp_bit[205]  <=   0;
          tmp_bit[206]  <=   0;
          tmp_bit[207]  <=   0;

       end else begin

// Ie4894ca167b08880bfc35862f18575eb Ied2b5c0139cec8ad2873829dc1117d50 clock start_d7 valid Ied2b5c0139cec8ad2873829dc1117d50 start_d7
           if (start_d7) begin
               tmp_bit[0]  <=   tmp_bit_0;
           end
           if (start_d7) begin
               tmp_bit[1]  <=   tmp_bit_1;
           end
           if (start_d7) begin
               tmp_bit[2]  <=   tmp_bit_2;
           end
           if (start_d7) begin
               tmp_bit[3]  <=   tmp_bit_3;
           end
           if (start_d7) begin
               tmp_bit[4]  <=   tmp_bit_4;
           end
           if (start_d7) begin
               tmp_bit[5]  <=   tmp_bit_5;
           end
           if (start_d7) begin
               tmp_bit[6]  <=   tmp_bit_6;
           end
           if (start_d7) begin
               tmp_bit[7]  <=   tmp_bit_7;
           end
           if (start_d7) begin
               tmp_bit[8]  <=   tmp_bit_8;
           end
           if (start_d7) begin
               tmp_bit[9]  <=   tmp_bit_9;
           end
           if (start_d7) begin
               tmp_bit[10]  <=   tmp_bit_10;
           end
           if (start_d7) begin
               tmp_bit[11]  <=   tmp_bit_11;
           end
           if (start_d7) begin
               tmp_bit[12]  <=   tmp_bit_12;
           end
           if (start_d7) begin
               tmp_bit[13]  <=   tmp_bit_13;
           end
           if (start_d7) begin
               tmp_bit[14]  <=   tmp_bit_14;
           end
           if (start_d7) begin
               tmp_bit[15]  <=   tmp_bit_15;
           end
           if (start_d7) begin
               tmp_bit[16]  <=   tmp_bit_16;
           end
           if (start_d7) begin
               tmp_bit[17]  <=   tmp_bit_17;
           end
           if (start_d7) begin
               tmp_bit[18]  <=   tmp_bit_18;
           end
           if (start_d7) begin
               tmp_bit[19]  <=   tmp_bit_19;
           end
           if (start_d7) begin
               tmp_bit[20]  <=   tmp_bit_20;
           end
           if (start_d7) begin
               tmp_bit[21]  <=   tmp_bit_21;
           end
           if (start_d7) begin
               tmp_bit[22]  <=   tmp_bit_22;
           end
           if (start_d7) begin
               tmp_bit[23]  <=   tmp_bit_23;
           end
           if (start_d7) begin
               tmp_bit[24]  <=   tmp_bit_24;
           end
           if (start_d7) begin
               tmp_bit[25]  <=   tmp_bit_25;
           end
           if (start_d7) begin
               tmp_bit[26]  <=   tmp_bit_26;
           end
           if (start_d7) begin
               tmp_bit[27]  <=   tmp_bit_27;
           end
           if (start_d7) begin
               tmp_bit[28]  <=   tmp_bit_28;
           end
           if (start_d7) begin
               tmp_bit[29]  <=   tmp_bit_29;
           end
           if (start_d7) begin
               tmp_bit[30]  <=   tmp_bit_30;
           end
           if (start_d7) begin
               tmp_bit[31]  <=   tmp_bit_31;
           end
           if (start_d7) begin
               tmp_bit[32]  <=   tmp_bit_32;
           end
           if (start_d7) begin
               tmp_bit[33]  <=   tmp_bit_33;
           end
           if (start_d7) begin
               tmp_bit[34]  <=   tmp_bit_34;
           end
           if (start_d7) begin
               tmp_bit[35]  <=   tmp_bit_35;
           end
           if (start_d7) begin
               tmp_bit[36]  <=   tmp_bit_36;
           end
           if (start_d7) begin
               tmp_bit[37]  <=   tmp_bit_37;
           end
           if (start_d7) begin
               tmp_bit[38]  <=   tmp_bit_38;
           end
           if (start_d7) begin
               tmp_bit[39]  <=   tmp_bit_39;
           end
           if (start_d7) begin
               tmp_bit[40]  <=   tmp_bit_40;
           end
           if (start_d7) begin
               tmp_bit[41]  <=   tmp_bit_41;
           end
           if (start_d7) begin
               tmp_bit[42]  <=   tmp_bit_42;
           end
           if (start_d7) begin
               tmp_bit[43]  <=   tmp_bit_43;
           end
           if (start_d7) begin
               tmp_bit[44]  <=   tmp_bit_44;
           end
           if (start_d7) begin
               tmp_bit[45]  <=   tmp_bit_45;
           end
           if (start_d7) begin
               tmp_bit[46]  <=   tmp_bit_46;
           end
           if (start_d7) begin
               tmp_bit[47]  <=   tmp_bit_47;
           end
           if (start_d7) begin
               tmp_bit[48]  <=   tmp_bit_48;
           end
           if (start_d7) begin
               tmp_bit[49]  <=   tmp_bit_49;
           end
           if (start_d7) begin
               tmp_bit[50]  <=   tmp_bit_50;
           end
           if (start_d7) begin
               tmp_bit[51]  <=   tmp_bit_51;
           end
           if (start_d7) begin
               tmp_bit[52]  <=   tmp_bit_52;
           end
           if (start_d7) begin
               tmp_bit[53]  <=   tmp_bit_53;
           end
           if (start_d7) begin
               tmp_bit[54]  <=   tmp_bit_54;
           end
           if (start_d7) begin
               tmp_bit[55]  <=   tmp_bit_55;
           end
           if (start_d7) begin
               tmp_bit[56]  <=   tmp_bit_56;
           end
           if (start_d7) begin
               tmp_bit[57]  <=   tmp_bit_57;
           end
           if (start_d7) begin
               tmp_bit[58]  <=   tmp_bit_58;
           end
           if (start_d7) begin
               tmp_bit[59]  <=   tmp_bit_59;
           end
           if (start_d7) begin
               tmp_bit[60]  <=   tmp_bit_60;
           end
           if (start_d7) begin
               tmp_bit[61]  <=   tmp_bit_61;
           end
           if (start_d7) begin
               tmp_bit[62]  <=   tmp_bit_62;
           end
           if (start_d7) begin
               tmp_bit[63]  <=   tmp_bit_63;
           end
           if (start_d7) begin
               tmp_bit[64]  <=   tmp_bit_64;
           end
           if (start_d7) begin
               tmp_bit[65]  <=   tmp_bit_65;
           end
           if (start_d7) begin
               tmp_bit[66]  <=   tmp_bit_66;
           end
           if (start_d7) begin
               tmp_bit[67]  <=   tmp_bit_67;
           end
           if (start_d7) begin
               tmp_bit[68]  <=   tmp_bit_68;
           end
           if (start_d7) begin
               tmp_bit[69]  <=   tmp_bit_69;
           end
           if (start_d7) begin
               tmp_bit[70]  <=   tmp_bit_70;
           end
           if (start_d7) begin
               tmp_bit[71]  <=   tmp_bit_71;
           end
           if (start_d7) begin
               tmp_bit[72]  <=   tmp_bit_72;
           end
           if (start_d7) begin
               tmp_bit[73]  <=   tmp_bit_73;
           end
           if (start_d7) begin
               tmp_bit[74]  <=   tmp_bit_74;
           end
           if (start_d7) begin
               tmp_bit[75]  <=   tmp_bit_75;
           end
           if (start_d7) begin
               tmp_bit[76]  <=   tmp_bit_76;
           end
           if (start_d7) begin
               tmp_bit[77]  <=   tmp_bit_77;
           end
           if (start_d7) begin
               tmp_bit[78]  <=   tmp_bit_78;
           end
           if (start_d7) begin
               tmp_bit[79]  <=   tmp_bit_79;
           end
           if (start_d7) begin
               tmp_bit[80]  <=   tmp_bit_80;
           end
           if (start_d7) begin
               tmp_bit[81]  <=   tmp_bit_81;
           end
           if (start_d7) begin
               tmp_bit[82]  <=   tmp_bit_82;
           end
           if (start_d7) begin
               tmp_bit[83]  <=   tmp_bit_83;
           end
           if (start_d7) begin
               tmp_bit[84]  <=   tmp_bit_84;
           end
           if (start_d7) begin
               tmp_bit[85]  <=   tmp_bit_85;
           end
           if (start_d7) begin
               tmp_bit[86]  <=   tmp_bit_86;
           end
           if (start_d7) begin
               tmp_bit[87]  <=   tmp_bit_87;
           end
           if (start_d7) begin
               tmp_bit[88]  <=   tmp_bit_88;
           end
           if (start_d7) begin
               tmp_bit[89]  <=   tmp_bit_89;
           end
           if (start_d7) begin
               tmp_bit[90]  <=   tmp_bit_90;
           end
           if (start_d7) begin
               tmp_bit[91]  <=   tmp_bit_91;
           end
           if (start_d7) begin
               tmp_bit[92]  <=   tmp_bit_92;
           end
           if (start_d7) begin
               tmp_bit[93]  <=   tmp_bit_93;
           end
           if (start_d7) begin
               tmp_bit[94]  <=   tmp_bit_94;
           end
           if (start_d7) begin
               tmp_bit[95]  <=   tmp_bit_95;
           end
           if (start_d7) begin
               tmp_bit[96]  <=   tmp_bit_96;
           end
           if (start_d7) begin
               tmp_bit[97]  <=   tmp_bit_97;
           end
           if (start_d7) begin
               tmp_bit[98]  <=   tmp_bit_98;
           end
           if (start_d7) begin
               tmp_bit[99]  <=   tmp_bit_99;
           end
           if (start_d7) begin
               tmp_bit[100]  <=   tmp_bit_100;
           end
           if (start_d7) begin
               tmp_bit[101]  <=   tmp_bit_101;
           end
           if (start_d7) begin
               tmp_bit[102]  <=   tmp_bit_102;
           end
           if (start_d7) begin
               tmp_bit[103]  <=   tmp_bit_103;
           end
           if (start_d7) begin
               tmp_bit[104]  <=   tmp_bit_104;
           end
           if (start_d7) begin
               tmp_bit[105]  <=   tmp_bit_105;
           end
           if (start_d7) begin
               tmp_bit[106]  <=   tmp_bit_106;
           end
           if (start_d7) begin
               tmp_bit[107]  <=   tmp_bit_107;
           end
           if (start_d7) begin
               tmp_bit[108]  <=   tmp_bit_108;
           end
           if (start_d7) begin
               tmp_bit[109]  <=   tmp_bit_109;
           end
           if (start_d7) begin
               tmp_bit[110]  <=   tmp_bit_110;
           end
           if (start_d7) begin
               tmp_bit[111]  <=   tmp_bit_111;
           end
           if (start_d7) begin
               tmp_bit[112]  <=   tmp_bit_112;
           end
           if (start_d7) begin
               tmp_bit[113]  <=   tmp_bit_113;
           end
           if (start_d7) begin
               tmp_bit[114]  <=   tmp_bit_114;
           end
           if (start_d7) begin
               tmp_bit[115]  <=   tmp_bit_115;
           end
           if (start_d7) begin
               tmp_bit[116]  <=   tmp_bit_116;
           end
           if (start_d7) begin
               tmp_bit[117]  <=   tmp_bit_117;
           end
           if (start_d7) begin
               tmp_bit[118]  <=   tmp_bit_118;
           end
           if (start_d7) begin
               tmp_bit[119]  <=   tmp_bit_119;
           end
           if (start_d7) begin
               tmp_bit[120]  <=   tmp_bit_120;
           end
           if (start_d7) begin
               tmp_bit[121]  <=   tmp_bit_121;
           end
           if (start_d7) begin
               tmp_bit[122]  <=   tmp_bit_122;
           end
           if (start_d7) begin
               tmp_bit[123]  <=   tmp_bit_123;
           end
           if (start_d7) begin
               tmp_bit[124]  <=   tmp_bit_124;
           end
           if (start_d7) begin
               tmp_bit[125]  <=   tmp_bit_125;
           end
           if (start_d7) begin
               tmp_bit[126]  <=   tmp_bit_126;
           end
           if (start_d7) begin
               tmp_bit[127]  <=   tmp_bit_127;
           end
           if (start_d7) begin
               tmp_bit[128]  <=   tmp_bit_128;
           end
           if (start_d7) begin
               tmp_bit[129]  <=   tmp_bit_129;
           end
           if (start_d7) begin
               tmp_bit[130]  <=   tmp_bit_130;
           end
           if (start_d7) begin
               tmp_bit[131]  <=   tmp_bit_131;
           end
           if (start_d7) begin
               tmp_bit[132]  <=   tmp_bit_132;
           end
           if (start_d7) begin
               tmp_bit[133]  <=   tmp_bit_133;
           end
           if (start_d7) begin
               tmp_bit[134]  <=   tmp_bit_134;
           end
           if (start_d7) begin
               tmp_bit[135]  <=   tmp_bit_135;
           end
           if (start_d7) begin
               tmp_bit[136]  <=   tmp_bit_136;
           end
           if (start_d7) begin
               tmp_bit[137]  <=   tmp_bit_137;
           end
           if (start_d7) begin
               tmp_bit[138]  <=   tmp_bit_138;
           end
           if (start_d7) begin
               tmp_bit[139]  <=   tmp_bit_139;
           end
           if (start_d7) begin
               tmp_bit[140]  <=   tmp_bit_140;
           end
           if (start_d7) begin
               tmp_bit[141]  <=   tmp_bit_141;
           end
           if (start_d7) begin
               tmp_bit[142]  <=   tmp_bit_142;
           end
           if (start_d7) begin
               tmp_bit[143]  <=   tmp_bit_143;
           end
           if (start_d7) begin
               tmp_bit[144]  <=   tmp_bit_144;
           end
           if (start_d7) begin
               tmp_bit[145]  <=   tmp_bit_145;
           end
           if (start_d7) begin
               tmp_bit[146]  <=   tmp_bit_146;
           end
           if (start_d7) begin
               tmp_bit[147]  <=   tmp_bit_147;
           end
           if (start_d7) begin
               tmp_bit[148]  <=   tmp_bit_148;
           end
           if (start_d7) begin
               tmp_bit[149]  <=   tmp_bit_149;
           end
           if (start_d7) begin
               tmp_bit[150]  <=   tmp_bit_150;
           end
           if (start_d7) begin
               tmp_bit[151]  <=   tmp_bit_151;
           end
           if (start_d7) begin
               tmp_bit[152]  <=   tmp_bit_152;
           end
           if (start_d7) begin
               tmp_bit[153]  <=   tmp_bit_153;
           end
           if (start_d7) begin
               tmp_bit[154]  <=   tmp_bit_154;
           end
           if (start_d7) begin
               tmp_bit[155]  <=   tmp_bit_155;
           end
           if (start_d7) begin
               tmp_bit[156]  <=   tmp_bit_156;
           end
           if (start_d7) begin
               tmp_bit[157]  <=   tmp_bit_157;
           end
           if (start_d7) begin
               tmp_bit[158]  <=   tmp_bit_158;
           end
           if (start_d7) begin
               tmp_bit[159]  <=   tmp_bit_159;
           end
           if (start_d7) begin
               tmp_bit[160]  <=   tmp_bit_160;
           end
           if (start_d7) begin
               tmp_bit[161]  <=   tmp_bit_161;
           end
           if (start_d7) begin
               tmp_bit[162]  <=   tmp_bit_162;
           end
           if (start_d7) begin
               tmp_bit[163]  <=   tmp_bit_163;
           end
           if (start_d7) begin
               tmp_bit[164]  <=   tmp_bit_164;
           end
           if (start_d7) begin
               tmp_bit[165]  <=   tmp_bit_165;
           end
           if (start_d7) begin
               tmp_bit[166]  <=   tmp_bit_166;
           end
           if (start_d7) begin
               tmp_bit[167]  <=   tmp_bit_167;
           end
           if (start_d7) begin
               tmp_bit[168]  <=   tmp_bit_168;
           end
           if (start_d7) begin
               tmp_bit[169]  <=   tmp_bit_169;
           end
           if (start_d7) begin
               tmp_bit[170]  <=   tmp_bit_170;
           end
           if (start_d7) begin
               tmp_bit[171]  <=   tmp_bit_171;
           end
           if (start_d7) begin
               tmp_bit[172]  <=   tmp_bit_172;
           end
           if (start_d7) begin
               tmp_bit[173]  <=   tmp_bit_173;
           end
           if (start_d7) begin
               tmp_bit[174]  <=   tmp_bit_174;
           end
           if (start_d7) begin
               tmp_bit[175]  <=   tmp_bit_175;
           end
           if (start_d7) begin
               tmp_bit[176]  <=   tmp_bit_176;
           end
           if (start_d7) begin
               tmp_bit[177]  <=   tmp_bit_177;
           end
           if (start_d7) begin
               tmp_bit[178]  <=   tmp_bit_178;
           end
           if (start_d7) begin
               tmp_bit[179]  <=   tmp_bit_179;
           end
           if (start_d7) begin
               tmp_bit[180]  <=   tmp_bit_180;
           end
           if (start_d7) begin
               tmp_bit[181]  <=   tmp_bit_181;
           end
           if (start_d7) begin
               tmp_bit[182]  <=   tmp_bit_182;
           end
           if (start_d7) begin
               tmp_bit[183]  <=   tmp_bit_183;
           end
           if (start_d7) begin
               tmp_bit[184]  <=   tmp_bit_184;
           end
           if (start_d7) begin
               tmp_bit[185]  <=   tmp_bit_185;
           end
           if (start_d7) begin
               tmp_bit[186]  <=   tmp_bit_186;
           end
           if (start_d7) begin
               tmp_bit[187]  <=   tmp_bit_187;
           end
           if (start_d7) begin
               tmp_bit[188]  <=   tmp_bit_188;
           end
           if (start_d7) begin
               tmp_bit[189]  <=   tmp_bit_189;
           end
           if (start_d7) begin
               tmp_bit[190]  <=   tmp_bit_190;
           end
           if (start_d7) begin
               tmp_bit[191]  <=   tmp_bit_191;
           end
           if (start_d7) begin
               tmp_bit[192]  <=   tmp_bit_192;
           end
           if (start_d7) begin
               tmp_bit[193]  <=   tmp_bit_193;
           end
           if (start_d7) begin
               tmp_bit[194]  <=   tmp_bit_194;
           end
           if (start_d7) begin
               tmp_bit[195]  <=   tmp_bit_195;
           end
           if (start_d7) begin
               tmp_bit[196]  <=   tmp_bit_196;
           end
           if (start_d7) begin
               tmp_bit[197]  <=   tmp_bit_197;
           end
           if (start_d7) begin
               tmp_bit[198]  <=   tmp_bit_198;
           end
           if (start_d7) begin
               tmp_bit[199]  <=   tmp_bit_199;
           end
           if (start_d7) begin
               tmp_bit[200]  <=   tmp_bit_200;
           end
           if (start_d7) begin
               tmp_bit[201]  <=   tmp_bit_201;
           end
           if (start_d7) begin
               tmp_bit[202]  <=   tmp_bit_202;
           end
           if (start_d7) begin
               tmp_bit[203]  <=   tmp_bit_203;
           end
           if (start_d7) begin
               tmp_bit[204]  <=   tmp_bit_204;
           end
           if (start_d7) begin
               tmp_bit[205]  <=   tmp_bit_205;
           end
           if (start_d7) begin
               tmp_bit[206]  <=   tmp_bit_206;
           end
           if (start_d7) begin
               tmp_bit[207]  <=   tmp_bit_207;
           end

       end
   end


`ifdef ENCRYPT
`endif

endmodule


module Ic9c2f173881d25f8976d723957809f51 #(
`include "NR_2_0_4/fgallag/GF2_LDPC_fgallag_param_inc.sv"

) (

input wire [fgallag_SEL - 1:0]       fgallag_sel ,
output reg [fgallag_WDTH  - 1:0]     fgallag,
input wire                           start_in,
output wire                          start_out,
input wire                           rstn,
input wire                           clk

);

`include "NR_2_0_4/fgallag/GF2_LDPC_fgallag_inc_inc_all.sv"

// fgallag::'h380
`include "NR_2_0_4/fgallag/GF2_LDPC_fgallag_inc_all.sv"

assign start_d_fgallag0x00000 = start_in;
assign start_out = start_d_fgallag0xffffffff_q;

always_comb
begin
     fgallag = fgallag0xffffffff_0_q;
end


endmodule







module Ic3da32f100a43f826b89a492544e7812 #(
`include "NR_2_0_4/flogtanh/GF2_LDPC_flogtanh_param_inc.sv"

) (

input wire [flogtanh_SEL - 1:0]      flogtanh_sel ,
output reg [flogtanh_WDTH  - 1:0]    flogtanh,
input wire                           start_in,
output wire                          start_out,
input wire                           rstn,
input wire                           clk

);

`include "NR_2_0_4/flogtanh/GF2_LDPC_flogtanh_inc_inc_all.sv"

// flogtanh::'h380
`include "NR_2_0_4/flogtanh/GF2_LDPC_flogtanh_inc_all.sv"

assign start_d_flogtanh0x00000 = start_in;
assign start_out = start_d_flogtanh0xffffffff_q;

always_comb
begin
     flogtanh = flogtanh0xffffffff_0_q;
end




endmodule




//C Ia642a85aab89544a289fb1f29eab689d: Ib6f6b4efd9391d1fa207d325ff1bbd60 I83878c91171338902e0fe0fb97a8c47a:0.100000 I7290d6b1f1458098d2f225877e609ba6:2.197225 percent_probability_int:'d141

 //Ic07b0b4d7660314f711a68fc47c4ab38 I48d8d6f5a3efbf52837d6b788a22859a valid code word
//y_int:
 //44010bdd34c9a17a9dc5c9798ef00a0604fe89b67904e634be0b
//syny_err:
 //0200400200100008100880c0000680200320002200
//C Ia642a85aab89544a289fb1f29eab689d: Ib6f6b4efd9391d1fa207d325ff1bbd60 I83878c91171338902e0fe0fb97a8c47a:0.038462 I7290d6b1f1458098d2f225877e609ba6:3.218876 percent_probability_int:'d206
