reg [flogtanh_WDTH -1:0] I85e2d7a9e28f224cac9188370cccc37b, Iba870e87f87c875ff098cafadf28d262;
reg [flogtanh_WDTH -1:0] I17540db3c63ade2b53e82ca752a6cd99, Icca31b5b8e9f944b504a02ba62118cc7;
reg [flogtanh_WDTH -1:0] I43b24a45247c83d2a986a6e352e7a38a, I43afe6aef28fcced58953c4b3a9b3eed;
reg [flogtanh_WDTH -1:0] I92680f7db736ef5df4e81244ffcff59b, Ieed89d20b342594d04aa6adca4cf2edf;
reg [flogtanh_WDTH -1:0] I39764779466097d56a3a65718704d030, Ibc5eb7267931e83838a653795dc809b1;
reg [flogtanh_WDTH -1:0] I1e7b702101a2cb5064b151835830a57d, Iedd54575ec8e5a76566ae1313faedb7c;
reg [flogtanh_WDTH -1:0] I57b599739f81aba00c5a7aa795ea08c8, I7b3ee2f269cb1f90235f1af617e5c3d9;
reg [flogtanh_WDTH -1:0] Ied56219095ff64722213c69d58e6b74f, I7935f561c946b80813603b40e7652f91;
reg [flogtanh_WDTH -1:0] I5fbce88eb0e5add5adc151439b070eff, I97c22b8b68524a584412c15361d761cc;
reg [flogtanh_WDTH -1:0] Ibaf106dee88a6d70caa3ca247be96938, I7d2a8ad5ee9f7a3e9d642735a85a9a23;
reg [flogtanh_WDTH -1:0] I47decd52e0f93d6281011a92a9a7081e, I07057436f307eac4f43cd5cb9274f963;
reg [flogtanh_WDTH -1:0] I4b74e2c1db97dcec11a65b57b1035acf, I2f4c421ebd4de08c8f660aa125eb06d3;
reg [flogtanh_WDTH -1:0] Ib8190cccfd6f5afb2b6cef33e5376d19, I760715bc18504dc4ef1f861035f6f8f7;
reg [flogtanh_WDTH -1:0] Icbc0f6167d607f74c80c23a3257cd2e1, If4e8fc4e2bbb39e7beb6db11b58d8232;
reg [flogtanh_WDTH -1:0] Ieac93250ec9be2ef318d48baf88b1ef5, I082a57b5a74e7e39bcf5d12acd15e272;
reg [flogtanh_WDTH -1:0] I5db1844e769af7943f93da66b475d99e, Ief8973860cdc98a7e4cce37573e3acb9;
reg [flogtanh_WDTH -1:0] I8f242f17610cae369dbfb2aaa0453b79, If72bc16b595b4a2f27b2639e2b033e39;
reg [flogtanh_WDTH -1:0] I5bebf7ec46791bfa6d1dad7eceeea034, Ibc2aacfd2026e5970b2ae172c703784b;
reg [flogtanh_WDTH -1:0] Ife8a533289756df000f25a54a51bcfe3, I71f0fb5ab1d8d8a20c53435e79081eef;
reg [flogtanh_WDTH -1:0] I5de464a27ad96e1c636efd974f129cfe, Ic7937c4ac4365348de1d96ece551555c;
reg [flogtanh_WDTH -1:0] I5f1b79389154a01c7d846f5f8774dfa7, I7f4db8e60704ff9f4b74094d188e0dda;
reg [flogtanh_WDTH -1:0] If3d70b7c1e8f802b887c01e068428a4e, I34ad34e3ccac9eb915309c29568da011;
reg [flogtanh_WDTH -1:0] Ic10bc44ab0b4ca1d588d768859f1bb35, Ia006bebb09394969493a92514c8713b5;
reg [flogtanh_WDTH -1:0] Ie3cd02462472a4430da14641cda50452, Ib2fbcacfe3daa5d49e950f5ebabf258f;
reg [flogtanh_WDTH -1:0] I3071dd54b8e3e01163a9d17df901a502, I98e3b2ac676d6e2555f2286631e0c43d;
reg [flogtanh_WDTH -1:0] I7fa902c92592761b9689aec509e9e68f, Iaaf05004e8c7866bb2ec1d46e76cd5a5;
reg [flogtanh_WDTH -1:0] I13ac2bb6eb27b06cc93e19bec590ac44, Idbde787e711114043d18cd262802b234;
reg [flogtanh_WDTH -1:0] Ied47c387d2e31433fbd752243e5e0aac, I061dc14bf9bc7b97d69893ab5b084f00;
reg [flogtanh_WDTH -1:0] I470d7fc38fd4e1b015a43ce4f898f2bd, Iaa784a3cc93b4939eb183ccc94bb8089;
reg [flogtanh_WDTH -1:0] If1f7c2655f45c9148824e4151ab448b6, Ifb75793136968aa2432e934f9e849695;
reg [flogtanh_WDTH -1:0] If120a179bc9b785016b64084d6e4d056, I3f333a2b43e5db6062346394119bfbaf;
reg [flogtanh_WDTH -1:0] I7fc7f688e30263828dfdaf9ec8ec2f7a, I3b0f64d1ae335c61b01f2209bcdc8333;
reg [flogtanh_WDTH -1:0] Ia8804339708717f01d9a9069c72f0fbb, Iccd3b8b6b6e2a4d60d81d4f367d971c7;
reg [flogtanh_WDTH -1:0] I5079e19864882aa577c73731fcee0a31, Iae2e1facdac5fd4726d1a6b77849b2f6;
reg [flogtanh_WDTH -1:0] Ia0dceddb9355f13a3a622f279c244f06, Iac2dd16556eed4d7f826f2063d8979ff;
reg [flogtanh_WDTH -1:0] I75a27f997d71f89b8beb0484ec0402d5, I879638f9da54bd5a8a5ff78f7b011739;
reg [flogtanh_WDTH -1:0] I6557d5a7415612889373a46ee77437c5, Ic4958fe74930007506b93064b9f87588;
reg [flogtanh_WDTH -1:0] Ieef6c1b5a0ec168747b3dedc3f88e803, If1618b6028dfd675842dc0fa24485ddf;
reg [flogtanh_WDTH -1:0] I892de6b0f85b4aea7ff9113d713552e2, If22a928365940b767923b37527ec904f;
reg [flogtanh_WDTH -1:0] Ie8c260c1c1a61ba194c563e25325b435, I8586e464f05f813699f9d466970085dd;
reg [flogtanh_WDTH -1:0] Ic34456cc9dc2004ffb6ac0974c98e0e4, I3bc0dcbecfbefea5fb1d0b617d0efa78;
reg [flogtanh_WDTH -1:0] I59e956b7f374eed213b25d05b702aa7b, I3ba79b98d30ac9111420c21e244bf338;
reg [flogtanh_WDTH -1:0] I3f03c8fa63d838b3d42c3f047e70fbf5, Id0e2a5919dcda34c1fcd9230d79d402c;
reg [flogtanh_WDTH -1:0] I3d899ecab223931d4c0e12833417e32b, I203eedac26099a1b191c73411c443e3d;
reg [flogtanh_WDTH -1:0] I1c56ccfd13ce759046362280dce3ef9c, I31bce9c2121ec3e7de33fd80027cdf38;
reg [flogtanh_WDTH -1:0] Icc0a9c979d7e154edb892315a4ca9cfd, I13702c5d75b212144cc0a3f060887b46;
reg [flogtanh_WDTH -1:0] Ieac7270ea1f936fea6df9fa9233a78a1, I4e3c3bcf1ca00767b813fec32d679779;
reg [flogtanh_WDTH -1:0] Id9a98abcca5f5bf46e2dce45066d2dd6, Iaabe6440ad8902891ba43f734d7c2935;
reg [flogtanh_WDTH -1:0] I240fa7efcb0d0196b865a47048e9f5e2, I69dc2265888e6ff99b608329353fb5b8;
reg [flogtanh_WDTH -1:0] I83a9fc44b887c9b860d07ba9d9a90083, I8c530fbe167efb1aca099e309bd8f250;
reg [flogtanh_WDTH -1:0] Ic20207f1d7c0f19dba8676141ca07549, Ic652a50c7dc405a941fe04abc2170434;
reg [flogtanh_WDTH -1:0] Ic4c14384ec86a331d36974bb41903efa, Ic9b544f863bc0820276ac101c90d38f0;
reg [flogtanh_WDTH -1:0] I87fab4038ff6c1bc1bcc170f9a202769, I3d5ba70412e03b55a77463d256016a7f;
reg [flogtanh_WDTH -1:0] I47e00ea6506dbd4a360baf94cf63dc2a, I842efe9f673c4d17759b83e4b6e86a4b;
reg [flogtanh_WDTH -1:0] Ia2683d4666dbf6b9f8befa2d6bdbbfcb, I23dfb343d3762798b72aec1aeb2f4b4d;
reg [flogtanh_WDTH -1:0] I1ed7dd07abe9aee415671c6222bdc16c, Ie31a29b6cf533af693f1a28483f6fb89;
reg [flogtanh_WDTH -1:0] I5ea7cfba8e7720077757862cf36ceaa2, I81ccdf38e45a3e285b02ef75c30b997d;
reg [flogtanh_WDTH -1:0] Ifb1ba203c0ec3fc5e1081393bf492c20, I3bd029d3007a94b52c72423af9f0ae79;
reg [flogtanh_WDTH -1:0] Id0417686b69b456644d09aaa861f26d4, I675db209cea9deaa18aaa4ace818d238;
reg [flogtanh_WDTH -1:0] I4c3cbe58c98f3e0fdf9c89b7143e50a3, I0a9c0baf5ac3e43feb41aec0c43df3de;
reg [flogtanh_WDTH -1:0] I0915e1427b7e3267e7ffe79d0cc782f3, Ifcd5afdf257eab5b1f6c7906290abdfd;
reg [flogtanh_WDTH -1:0] Id5a895fa3677c1f973675aebec6b41f2, I335e3a7dd9a8baa6412527ef292ea90c;
reg [flogtanh_WDTH -1:0] I023b610b050357cc816939b6508bedb9, Ie801d81c4251559ca6661da90df75c79;
reg [flogtanh_WDTH -1:0] Ia7f89e3fc13d2589f1a2a025830a8b9e, Ide9dd8e36e4508731c54d883e4a2e2ee;
reg [flogtanh_WDTH -1:0] I51c00546226c98d468b69a85d8613b4d, Iaedb40c3bffbe0928b2b23275b85ddd4;
reg [flogtanh_WDTH -1:0] Ie5f68f657e8123b2e971d4f3e5a675df, Id8e69f2913aa400a3d03702076af5c2b;
reg [flogtanh_WDTH -1:0] Ia9194d615d26094f0c3e0399ab2e3da3, I7acb86a7e521fad3f1123b86e310b18a;
reg [flogtanh_WDTH -1:0] I9f1ef03445a07c36defabb3abd5df4c4, If9f8f260dff9690b3346854b71290cc8;
reg [flogtanh_WDTH -1:0] I8f90fcb8534f00216e0f6c4a3dbad2f6, I86df045ba01e5daeb569d9ea1a3263d7;
reg [flogtanh_WDTH -1:0] I30166adbb988446bdb36723a2e4cd7c1, I2daa598dc2f08ceae2895b81ef43a742;
reg [flogtanh_WDTH -1:0] Ief50b2820a6d32e602d4963c13b3f630, I0583dbd1d4e65defd1ba2fbe2bd87d0a;
reg [flogtanh_WDTH -1:0] If51760e69ff89f244fdb9cdb0b93bda4, I1a7a8ed99d0d10bcefd5a51600d1ceb6;
reg [flogtanh_WDTH -1:0] Idf43504868969d00511ef6e8d809db66, Ic541d5047749fb2833bfa23bad86e2ae;
reg [flogtanh_WDTH -1:0] Icfc6c999050d945d3a381ba869dd6e76, Ie28cded64c2871f0632dc9ba10be2738;
reg [flogtanh_WDTH -1:0] Iec57a1e76f07f3c328f74bfe5b1da785, I02cfa4d934a334809afc76213ef6cdff;
reg [flogtanh_WDTH -1:0] Ice973d37ca9816e4e5b7221463d76636, Ic5c8fef9f84b9de0aac6d91be393d8d6;
reg [flogtanh_WDTH -1:0] I87c9f04f74686c1dee6305deb51b9007, I75c142058c4a21b970356e0575e2d025;
reg [flogtanh_WDTH -1:0] I9350b76d99dd94589a9997500354f19d, I9896c94b6a97b16d440b3c0926fc85aa;
reg [flogtanh_WDTH -1:0] Idd0acb6b0bc3d9e3a12715d4f6614149, I561431791c47fa1b7455126752aac55e;
reg [flogtanh_WDTH -1:0] Idab3e6bf2379a457d67cce07ca31ba57, I7ece0fbda1ad50ea064dd79f1b9b243c;
reg [flogtanh_WDTH -1:0] Ie2f28a6c2445f5178eecc13507b72323, I5004693a6347e9b31037639942d06504;
reg [flogtanh_WDTH -1:0] I5d3b6f0d046829b096807ab4a49bcc25, I367d8953c0e23856140cf4785d929d91;
reg [flogtanh_WDTH -1:0] I0b3c995b0a12a14265de007d90300cec, I73709d12931c354b73a1369cac5db3a9;
reg [flogtanh_WDTH -1:0] I31b53846b721e11cddea32c4b046a7fa, Ia0225847ade3d5db93ae32d6d7d83eee;
reg [flogtanh_WDTH -1:0] I1b40caccc7bf0db9618dd54d2959ee2a, I6e3a3dc54544c2601df65e24390247e4;
reg [flogtanh_WDTH -1:0] I832959dc65f560a892c99dc05dfb19ff, I2ddf3dd926d1966b8b82e421da6a9675;
reg [flogtanh_WDTH -1:0] I515dd393df02b089c3afa5ef912c945a, Ia7d3383c61357b1b2fa53a9f3728a3da;
reg [flogtanh_WDTH -1:0] I55b2317ed99a99a1afd11aff3c296683, I629e0f0fae704938defa7dccef6eb675;
reg [flogtanh_WDTH -1:0] I8122943006aece7452a503e8c20375b4, I1a296cef71412b570eaa40a564f146e2;
reg [flogtanh_WDTH -1:0] Ida9814058169631dca9f83ee34741a75, Ib34c55a2554033229a576daae46633f1;
reg If6d744ed5db03bac562b8bea5fd72479 ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 Iba870e87f87c875ff098cafadf28d262 <= 'h0;
 Icca31b5b8e9f944b504a02ba62118cc7 <= 'h0;
 I43afe6aef28fcced58953c4b3a9b3eed <= 'h0;
 Ieed89d20b342594d04aa6adca4cf2edf <= 'h0;
 Ibc5eb7267931e83838a653795dc809b1 <= 'h0;
 Iedd54575ec8e5a76566ae1313faedb7c <= 'h0;
 I7b3ee2f269cb1f90235f1af617e5c3d9 <= 'h0;
 I7935f561c946b80813603b40e7652f91 <= 'h0;
 I97c22b8b68524a584412c15361d761cc <= 'h0;
 I7d2a8ad5ee9f7a3e9d642735a85a9a23 <= 'h0;
 I07057436f307eac4f43cd5cb9274f963 <= 'h0;
 I2f4c421ebd4de08c8f660aa125eb06d3 <= 'h0;
 I760715bc18504dc4ef1f861035f6f8f7 <= 'h0;
 If4e8fc4e2bbb39e7beb6db11b58d8232 <= 'h0;
 I082a57b5a74e7e39bcf5d12acd15e272 <= 'h0;
 Ief8973860cdc98a7e4cce37573e3acb9 <= 'h0;
 If72bc16b595b4a2f27b2639e2b033e39 <= 'h0;
 Ibc2aacfd2026e5970b2ae172c703784b <= 'h0;
 I71f0fb5ab1d8d8a20c53435e79081eef <= 'h0;
 Ic7937c4ac4365348de1d96ece551555c <= 'h0;
 I7f4db8e60704ff9f4b74094d188e0dda <= 'h0;
 I34ad34e3ccac9eb915309c29568da011 <= 'h0;
 Ia006bebb09394969493a92514c8713b5 <= 'h0;
 Ib2fbcacfe3daa5d49e950f5ebabf258f <= 'h0;
 I98e3b2ac676d6e2555f2286631e0c43d <= 'h0;
 Iaaf05004e8c7866bb2ec1d46e76cd5a5 <= 'h0;
 Idbde787e711114043d18cd262802b234 <= 'h0;
 I061dc14bf9bc7b97d69893ab5b084f00 <= 'h0;
 Iaa784a3cc93b4939eb183ccc94bb8089 <= 'h0;
 Ifb75793136968aa2432e934f9e849695 <= 'h0;
 I3f333a2b43e5db6062346394119bfbaf <= 'h0;
 I3b0f64d1ae335c61b01f2209bcdc8333 <= 'h0;
 Iccd3b8b6b6e2a4d60d81d4f367d971c7 <= 'h0;
 Iae2e1facdac5fd4726d1a6b77849b2f6 <= 'h0;
 Iac2dd16556eed4d7f826f2063d8979ff <= 'h0;
 I879638f9da54bd5a8a5ff78f7b011739 <= 'h0;
 Ic4958fe74930007506b93064b9f87588 <= 'h0;
 If1618b6028dfd675842dc0fa24485ddf <= 'h0;
 If22a928365940b767923b37527ec904f <= 'h0;
 I8586e464f05f813699f9d466970085dd <= 'h0;
 I3bc0dcbecfbefea5fb1d0b617d0efa78 <= 'h0;
 I3ba79b98d30ac9111420c21e244bf338 <= 'h0;
 Id0e2a5919dcda34c1fcd9230d79d402c <= 'h0;
 I203eedac26099a1b191c73411c443e3d <= 'h0;
 I31bce9c2121ec3e7de33fd80027cdf38 <= 'h0;
 I13702c5d75b212144cc0a3f060887b46 <= 'h0;
 I4e3c3bcf1ca00767b813fec32d679779 <= 'h0;
 Iaabe6440ad8902891ba43f734d7c2935 <= 'h0;
 I69dc2265888e6ff99b608329353fb5b8 <= 'h0;
 I8c530fbe167efb1aca099e309bd8f250 <= 'h0;
 Ic652a50c7dc405a941fe04abc2170434 <= 'h0;
 Ic9b544f863bc0820276ac101c90d38f0 <= 'h0;
 I3d5ba70412e03b55a77463d256016a7f <= 'h0;
 I842efe9f673c4d17759b83e4b6e86a4b <= 'h0;
 I23dfb343d3762798b72aec1aeb2f4b4d <= 'h0;
 Ie31a29b6cf533af693f1a28483f6fb89 <= 'h0;
 I81ccdf38e45a3e285b02ef75c30b997d <= 'h0;
 I3bd029d3007a94b52c72423af9f0ae79 <= 'h0;
 I675db209cea9deaa18aaa4ace818d238 <= 'h0;
 I0a9c0baf5ac3e43feb41aec0c43df3de <= 'h0;
 Ifcd5afdf257eab5b1f6c7906290abdfd <= 'h0;
 I335e3a7dd9a8baa6412527ef292ea90c <= 'h0;
 Ie801d81c4251559ca6661da90df75c79 <= 'h0;
 Ide9dd8e36e4508731c54d883e4a2e2ee <= 'h0;
 Iaedb40c3bffbe0928b2b23275b85ddd4 <= 'h0;
 Id8e69f2913aa400a3d03702076af5c2b <= 'h0;
 I7acb86a7e521fad3f1123b86e310b18a <= 'h0;
 If9f8f260dff9690b3346854b71290cc8 <= 'h0;
 I86df045ba01e5daeb569d9ea1a3263d7 <= 'h0;
 I2daa598dc2f08ceae2895b81ef43a742 <= 'h0;
 I0583dbd1d4e65defd1ba2fbe2bd87d0a <= 'h0;
 I1a7a8ed99d0d10bcefd5a51600d1ceb6 <= 'h0;
 Ic541d5047749fb2833bfa23bad86e2ae <= 'h0;
 Ie28cded64c2871f0632dc9ba10be2738 <= 'h0;
 I02cfa4d934a334809afc76213ef6cdff <= 'h0;
 Ic5c8fef9f84b9de0aac6d91be393d8d6 <= 'h0;
 I75c142058c4a21b970356e0575e2d025 <= 'h0;
 I9896c94b6a97b16d440b3c0926fc85aa <= 'h0;
 I561431791c47fa1b7455126752aac55e <= 'h0;
 I7ece0fbda1ad50ea064dd79f1b9b243c <= 'h0;
 I5004693a6347e9b31037639942d06504 <= 'h0;
 I367d8953c0e23856140cf4785d929d91 <= 'h0;
 I73709d12931c354b73a1369cac5db3a9 <= 'h0;
 Ia0225847ade3d5db93ae32d6d7d83eee <= 'h0;
 I6e3a3dc54544c2601df65e24390247e4 <= 'h0;
 I2ddf3dd926d1966b8b82e421da6a9675 <= 'h0;
 Ia7d3383c61357b1b2fa53a9f3728a3da <= 'h0;
 I629e0f0fae704938defa7dccef6eb675 <= 'h0;
 I1a296cef71412b570eaa40a564f146e2 <= 'h0;
 Ib34c55a2554033229a576daae46633f1 <= 'h0;
 If6d744ed5db03bac562b8bea5fd72479 <= 'h0;
end
else
begin
 Iba870e87f87c875ff098cafadf28d262 <=  I85e2d7a9e28f224cac9188370cccc37b;
 Icca31b5b8e9f944b504a02ba62118cc7 <=  I17540db3c63ade2b53e82ca752a6cd99;
 I43afe6aef28fcced58953c4b3a9b3eed <=  I43b24a45247c83d2a986a6e352e7a38a;
 Ieed89d20b342594d04aa6adca4cf2edf <=  I92680f7db736ef5df4e81244ffcff59b;
 Ibc5eb7267931e83838a653795dc809b1 <=  I39764779466097d56a3a65718704d030;
 Iedd54575ec8e5a76566ae1313faedb7c <=  I1e7b702101a2cb5064b151835830a57d;
 I7b3ee2f269cb1f90235f1af617e5c3d9 <=  I57b599739f81aba00c5a7aa795ea08c8;
 I7935f561c946b80813603b40e7652f91 <=  Ied56219095ff64722213c69d58e6b74f;
 I97c22b8b68524a584412c15361d761cc <=  I5fbce88eb0e5add5adc151439b070eff;
 I7d2a8ad5ee9f7a3e9d642735a85a9a23 <=  Ibaf106dee88a6d70caa3ca247be96938;
 I07057436f307eac4f43cd5cb9274f963 <=  I47decd52e0f93d6281011a92a9a7081e;
 I2f4c421ebd4de08c8f660aa125eb06d3 <=  I4b74e2c1db97dcec11a65b57b1035acf;
 I760715bc18504dc4ef1f861035f6f8f7 <=  Ib8190cccfd6f5afb2b6cef33e5376d19;
 If4e8fc4e2bbb39e7beb6db11b58d8232 <=  Icbc0f6167d607f74c80c23a3257cd2e1;
 I082a57b5a74e7e39bcf5d12acd15e272 <=  Ieac93250ec9be2ef318d48baf88b1ef5;
 Ief8973860cdc98a7e4cce37573e3acb9 <=  I5db1844e769af7943f93da66b475d99e;
 If72bc16b595b4a2f27b2639e2b033e39 <=  I8f242f17610cae369dbfb2aaa0453b79;
 Ibc2aacfd2026e5970b2ae172c703784b <=  I5bebf7ec46791bfa6d1dad7eceeea034;
 I71f0fb5ab1d8d8a20c53435e79081eef <=  Ife8a533289756df000f25a54a51bcfe3;
 Ic7937c4ac4365348de1d96ece551555c <=  I5de464a27ad96e1c636efd974f129cfe;
 I7f4db8e60704ff9f4b74094d188e0dda <=  I5f1b79389154a01c7d846f5f8774dfa7;
 I34ad34e3ccac9eb915309c29568da011 <=  If3d70b7c1e8f802b887c01e068428a4e;
 Ia006bebb09394969493a92514c8713b5 <=  Ic10bc44ab0b4ca1d588d768859f1bb35;
 Ib2fbcacfe3daa5d49e950f5ebabf258f <=  Ie3cd02462472a4430da14641cda50452;
 I98e3b2ac676d6e2555f2286631e0c43d <=  I3071dd54b8e3e01163a9d17df901a502;
 Iaaf05004e8c7866bb2ec1d46e76cd5a5 <=  I7fa902c92592761b9689aec509e9e68f;
 Idbde787e711114043d18cd262802b234 <=  I13ac2bb6eb27b06cc93e19bec590ac44;
 I061dc14bf9bc7b97d69893ab5b084f00 <=  Ied47c387d2e31433fbd752243e5e0aac;
 Iaa784a3cc93b4939eb183ccc94bb8089 <=  I470d7fc38fd4e1b015a43ce4f898f2bd;
 Ifb75793136968aa2432e934f9e849695 <=  If1f7c2655f45c9148824e4151ab448b6;
 I3f333a2b43e5db6062346394119bfbaf <=  If120a179bc9b785016b64084d6e4d056;
 I3b0f64d1ae335c61b01f2209bcdc8333 <=  I7fc7f688e30263828dfdaf9ec8ec2f7a;
 Iccd3b8b6b6e2a4d60d81d4f367d971c7 <=  Ia8804339708717f01d9a9069c72f0fbb;
 Iae2e1facdac5fd4726d1a6b77849b2f6 <=  I5079e19864882aa577c73731fcee0a31;
 Iac2dd16556eed4d7f826f2063d8979ff <=  Ia0dceddb9355f13a3a622f279c244f06;
 I879638f9da54bd5a8a5ff78f7b011739 <=  I75a27f997d71f89b8beb0484ec0402d5;
 Ic4958fe74930007506b93064b9f87588 <=  I6557d5a7415612889373a46ee77437c5;
 If1618b6028dfd675842dc0fa24485ddf <=  Ieef6c1b5a0ec168747b3dedc3f88e803;
 If22a928365940b767923b37527ec904f <=  I892de6b0f85b4aea7ff9113d713552e2;
 I8586e464f05f813699f9d466970085dd <=  Ie8c260c1c1a61ba194c563e25325b435;
 I3bc0dcbecfbefea5fb1d0b617d0efa78 <=  Ic34456cc9dc2004ffb6ac0974c98e0e4;
 I3ba79b98d30ac9111420c21e244bf338 <=  I59e956b7f374eed213b25d05b702aa7b;
 Id0e2a5919dcda34c1fcd9230d79d402c <=  I3f03c8fa63d838b3d42c3f047e70fbf5;
 I203eedac26099a1b191c73411c443e3d <=  I3d899ecab223931d4c0e12833417e32b;
 I31bce9c2121ec3e7de33fd80027cdf38 <=  I1c56ccfd13ce759046362280dce3ef9c;
 I13702c5d75b212144cc0a3f060887b46 <=  Icc0a9c979d7e154edb892315a4ca9cfd;
 I4e3c3bcf1ca00767b813fec32d679779 <=  Ieac7270ea1f936fea6df9fa9233a78a1;
 Iaabe6440ad8902891ba43f734d7c2935 <=  Id9a98abcca5f5bf46e2dce45066d2dd6;
 I69dc2265888e6ff99b608329353fb5b8 <=  I240fa7efcb0d0196b865a47048e9f5e2;
 I8c530fbe167efb1aca099e309bd8f250 <=  I83a9fc44b887c9b860d07ba9d9a90083;
 Ic652a50c7dc405a941fe04abc2170434 <=  Ic20207f1d7c0f19dba8676141ca07549;
 Ic9b544f863bc0820276ac101c90d38f0 <=  Ic4c14384ec86a331d36974bb41903efa;
 I3d5ba70412e03b55a77463d256016a7f <=  I87fab4038ff6c1bc1bcc170f9a202769;
 I842efe9f673c4d17759b83e4b6e86a4b <=  I47e00ea6506dbd4a360baf94cf63dc2a;
 I23dfb343d3762798b72aec1aeb2f4b4d <=  Ia2683d4666dbf6b9f8befa2d6bdbbfcb;
 Ie31a29b6cf533af693f1a28483f6fb89 <=  I1ed7dd07abe9aee415671c6222bdc16c;
 I81ccdf38e45a3e285b02ef75c30b997d <=  I5ea7cfba8e7720077757862cf36ceaa2;
 I3bd029d3007a94b52c72423af9f0ae79 <=  Ifb1ba203c0ec3fc5e1081393bf492c20;
 I675db209cea9deaa18aaa4ace818d238 <=  Id0417686b69b456644d09aaa861f26d4;
 I0a9c0baf5ac3e43feb41aec0c43df3de <=  I4c3cbe58c98f3e0fdf9c89b7143e50a3;
 Ifcd5afdf257eab5b1f6c7906290abdfd <=  I0915e1427b7e3267e7ffe79d0cc782f3;
 I335e3a7dd9a8baa6412527ef292ea90c <=  Id5a895fa3677c1f973675aebec6b41f2;
 Ie801d81c4251559ca6661da90df75c79 <=  I023b610b050357cc816939b6508bedb9;
 Ide9dd8e36e4508731c54d883e4a2e2ee <=  Ia7f89e3fc13d2589f1a2a025830a8b9e;
 Iaedb40c3bffbe0928b2b23275b85ddd4 <=  I51c00546226c98d468b69a85d8613b4d;
 Id8e69f2913aa400a3d03702076af5c2b <=  Ie5f68f657e8123b2e971d4f3e5a675df;
 I7acb86a7e521fad3f1123b86e310b18a <=  Ia9194d615d26094f0c3e0399ab2e3da3;
 If9f8f260dff9690b3346854b71290cc8 <=  I9f1ef03445a07c36defabb3abd5df4c4;
 I86df045ba01e5daeb569d9ea1a3263d7 <=  I8f90fcb8534f00216e0f6c4a3dbad2f6;
 I2daa598dc2f08ceae2895b81ef43a742 <=  I30166adbb988446bdb36723a2e4cd7c1;
 I0583dbd1d4e65defd1ba2fbe2bd87d0a <=  Ief50b2820a6d32e602d4963c13b3f630;
 I1a7a8ed99d0d10bcefd5a51600d1ceb6 <=  If51760e69ff89f244fdb9cdb0b93bda4;
 Ic541d5047749fb2833bfa23bad86e2ae <=  Idf43504868969d00511ef6e8d809db66;
 Ie28cded64c2871f0632dc9ba10be2738 <=  Icfc6c999050d945d3a381ba869dd6e76;
 I02cfa4d934a334809afc76213ef6cdff <=  Iec57a1e76f07f3c328f74bfe5b1da785;
 Ic5c8fef9f84b9de0aac6d91be393d8d6 <=  Ice973d37ca9816e4e5b7221463d76636;
 I75c142058c4a21b970356e0575e2d025 <=  I87c9f04f74686c1dee6305deb51b9007;
 I9896c94b6a97b16d440b3c0926fc85aa <=  I9350b76d99dd94589a9997500354f19d;
 I561431791c47fa1b7455126752aac55e <=  Idd0acb6b0bc3d9e3a12715d4f6614149;
 I7ece0fbda1ad50ea064dd79f1b9b243c <=  Idab3e6bf2379a457d67cce07ca31ba57;
 I5004693a6347e9b31037639942d06504 <=  Ie2f28a6c2445f5178eecc13507b72323;
 I367d8953c0e23856140cf4785d929d91 <=  I5d3b6f0d046829b096807ab4a49bcc25;
 I73709d12931c354b73a1369cac5db3a9 <=  I0b3c995b0a12a14265de007d90300cec;
 Ia0225847ade3d5db93ae32d6d7d83eee <=  I31b53846b721e11cddea32c4b046a7fa;
 I6e3a3dc54544c2601df65e24390247e4 <=  I1b40caccc7bf0db9618dd54d2959ee2a;
 I2ddf3dd926d1966b8b82e421da6a9675 <=  I832959dc65f560a892c99dc05dfb19ff;
 Ia7d3383c61357b1b2fa53a9f3728a3da <=  I515dd393df02b089c3afa5ef912c945a;
 I629e0f0fae704938defa7dccef6eb675 <=  I55b2317ed99a99a1afd11aff3c296683;
 I1a296cef71412b570eaa40a564f146e2 <=  I8122943006aece7452a503e8c20375b4;
 Ib34c55a2554033229a576daae46633f1 <=  Ida9814058169631dca9f83ee34741a75;
 If6d744ed5db03bac562b8bea5fd72479 <=  Icf92b5275d264e1b6d832272a0d01a66;
end
