 reg  ['hffff:0] [$clog2('h7000+1)-1:0] Ia439aa2748f2eda0e2e55cce3a9fa0dee631b8aa10765b3a86df54c955466e56 ;
