reg [fgallag_WDTH -1:0] I9c9ab24ecd80ca61b89534e3e5adfca8, Ia6f93d7eab83c88b604f8a81a74c04e9;
reg [fgallag_WDTH -1:0] Ie92d645c17dda47f594bc34b0937caac, Ice05aa8a4d2a062da9785286081fd024;
reg [fgallag_WDTH -1:0] Ieb8b25a5f6d3cc4cead3f3845234d1d3, I6e41efdbe6eeb41b9c9b39e56f3d8b9c;
reg [fgallag_WDTH -1:0] Ibcbdbe8034a373448800d1b745cb5849, Ibe53a3b8a9caa8643361263d463290c8;
reg [fgallag_WDTH -1:0] Ibd0769c69670150d8263d9873cbf668f, Ifbcddebb5f791d2df0b2e7aa94a81c22;
reg [fgallag_WDTH -1:0] I2010cff1e77f9706d8c659482f51c898, I341146b894d9d94c2c803e6b6c464085;
reg [fgallag_WDTH -1:0] I4183447a1a1727e91b0fcabb9bec1963, Iccfcaba2f6129c8201cb97323a8e740a;
reg [fgallag_WDTH -1:0] I780bea956f609c6f3cd0ffd126f99316, I850f7b404a1ab022498350d9ef0cbdc2;
reg [fgallag_WDTH -1:0] I349cff38817dd1607e798b9a2ae6fb8b, Ie88f3ca2bc79208be9385225a7ad7268;
reg [fgallag_WDTH -1:0] I3ff605a8af8eceb2c055e842e6208958, If4137d66b193970e9ae89b8e1b00e8ca;
reg [fgallag_WDTH -1:0] Ib53b2b0d39dbe6d09f51e0af27e5986f, I877047b00cef1f6a938ed9915215e203;
reg [fgallag_WDTH -1:0] I343242367c13febc05ee63f57dd4f754, Ic9e529e5e428a666bf6bcf2041969d1e;
reg [fgallag_WDTH -1:0] Ibde6749f31c571c5209a8b36c1c8f4da, I2e8ce46a773bcf5f2c3129441a267af4;
reg [fgallag_WDTH -1:0] Ib735324969bc744cc0ab8c2b3a7c5561, Ie734c46bfea46055c73a2642b3f8a7da;
reg [fgallag_WDTH -1:0] If53ed28774233bca87090e799465e3a5, Id980a518f6b9c84062f5bd7d6f57472f;
reg [fgallag_WDTH -1:0] Ib5017be08e079fe946c365fc01461d11, I8901003e5fb9f89fddb0fa87dc5b2d05;
reg [fgallag_WDTH -1:0] I0f24b1ca1d272d4971cde83a2acfe5ac, Ia5402393b456807ca5fee0ecb219c7d9;
reg [fgallag_WDTH -1:0] I1d1f2f5dd46b3f89c5a614ebad298d13, I41d38680c5aca0364ef9c716cd4525e7;
reg [fgallag_WDTH -1:0] I09dbcf2140141aaa400ad52408f8ab41, I03ee8c787b49b08c0a5a503bd28fcca5;
reg [fgallag_WDTH -1:0] I8315726dd19b5074a78796ee704d7108, Id85bac587e9c200406f0aecafbaf3dd5;
reg [fgallag_WDTH -1:0] Idb03654ee570200d2fe82907af7095d7, Ibb5dbc2fc80aca18dbaa13b7ecdb6c20;
reg [fgallag_WDTH -1:0] I9a5f25915425b586c1c3979240ff1a54, I9b5df9c23c9a2aaa14a99abd110075cb;
reg [fgallag_WDTH -1:0] I259241ceeda0568e6c10162cd43ca1dc, Ic00f5a4dfdbbf58316107417ccc6bb74;
reg [fgallag_WDTH -1:0] I66d1b07d77d2fe21d535920b30e176ff, Ic208118fb71fea311016edcb1203407d;
reg [fgallag_WDTH -1:0] I135dcccb8e63f697fe4559b964322345, Ib3d96f215fc42ace8fddda8c64afbc05;
reg [fgallag_WDTH -1:0] Ic37c4058485edfc0ca4f12fd7a97bf93, Ie304d02670ae74fb93fb42328d43079e;
reg [fgallag_WDTH -1:0] I1400488e51bbe6c921439713342d39f8, I1a875fdb7e3681839eeb5fdb8c6b47c3;
reg [fgallag_WDTH -1:0] Iaa8359974e7a41f754b38d6a232c5e72, I85c6964245f5e3423ddfcae7ae864429;
reg [fgallag_WDTH -1:0] Ie99b9c10b4b5208374b9f4ba1bd3eeab, Idd3396a16fde9c928bfd71f9b05b98bf;
reg [fgallag_WDTH -1:0] I54462091230adebf4bf4ec0cea25e374, I3a124ec3bd01d433c39ecbfd0b153d74;
reg [fgallag_WDTH -1:0] Iba9e737dd791a2ee966dbf6958339d65, I7be57c1f60b38d43d0fe2c02175aeef5;
reg [fgallag_WDTH -1:0] Ib205f5f9a6005baa465f1b254e4014d0, I886a56b1cae34e1860e4cd2c28606a45;
reg [fgallag_WDTH -1:0] I5ea13e282884d2343e8fdbe17d7ee058, I4dfc6b1e7b358ad6a32f6682e487d962;
reg [fgallag_WDTH -1:0] I6d8ed091d5f44b3b49e8b0eb63f0d106, I4c60daf9c53a50f2a228ca9ad0d75115;
reg [fgallag_WDTH -1:0] I4109473d968250506e17f8227bc55d06, I5fa487af5385cb6dcd0bac274a2b2261;
reg [fgallag_WDTH -1:0] Ia7da78b0d37028fcd34d3d39c7e36596, If3024e217350078f9a06275cc31b6699;
reg [fgallag_WDTH -1:0] I034454a1608fbde69fffb6b28e685f9f, Ifb39ced2cc4424e46be38af68161181a;
reg [fgallag_WDTH -1:0] I6e487d671a19855fd1eae42664d9c57f, I17934cad1385024244ce8bd07b709db0;
reg [fgallag_WDTH -1:0] Ib49b6b6895bd7200dc9e026584bea017, Ie43b90c9bb7dcb76f116c75615df246b;
reg [fgallag_WDTH -1:0] I220ce4284bf6adf0e46cf524b04a0e1b, I7f095ecd42b65b1781e2290db664a73d;
reg [fgallag_WDTH -1:0] I64586e3b7241a57c2e887b651819c7f9, I4d7c79dc1c72745d5750cac86454beb8;
reg [fgallag_WDTH -1:0] Ifad0bf7a3d7d334b5f8ea0d1a973fd39, I00c66baa19546590a542100f8883d4ab;
reg [fgallag_WDTH -1:0] If060b99963382d16c1f779faf00a7128, I97293ec9139e6e252c554d9f26619f06;
reg [fgallag_WDTH -1:0] Ie80ad5b1c3c4046c80e6cb96ee51e5c0, I067a46089f564be32860d44b3c69af1a;
reg [fgallag_WDTH -1:0] I4fe400daeacdfbebafcdf7e753af2787, Ib11764f9c254c7ddf0782d0cccae0067;
reg [fgallag_WDTH -1:0] I5c1ec1001d1ea61ab7198336742ed99d, Ic63385ac292f30c59ab2ad6f8b7d8903;
reg [fgallag_WDTH -1:0] If50cfdca6c9b8000665da2513244ff24, I5d3f02e43c3a9ab32c9769c1cf45ec6c;
reg [fgallag_WDTH -1:0] I4367feaf57687befa18bc6a902573bb9, I968edb5f5a70a3d391db21db00dafe78;
reg [fgallag_WDTH -1:0] I8f2820928683d8d88d41b80a9d9832dd, I59ad05479adc69422b7e06e4507a8f7a;
reg [fgallag_WDTH -1:0] Id980002a738b3ab2a4c2ccb9d232d141, I3755b61b6fb958538b1b906a4ad1103d;
reg [fgallag_WDTH -1:0] Ib1db1798d076dc0a6fa322c47e0ac062, I0ba5990e179758e1080a8407412a9a59;
reg [fgallag_WDTH -1:0] Iba73f7b76a2e16d7d84cfbab4473143d, I7562a62ae85c4676605b60594722a950;
reg [fgallag_WDTH -1:0] Iad0a6e20283bbf4bd4114a0c70c0685e, I62c2ba2ded74107adfcbe43670718e65;
reg [fgallag_WDTH -1:0] Ic772211084626d2ed3ddc4f32b467c6c, Ie43871350b062263474a7e0dbca850ce;
reg [fgallag_WDTH -1:0] Ifcba38a9a6ca0931ba9d86396f257929, I12d1f6ac4ef39cb76907b09745b4f8ad;
reg [fgallag_WDTH -1:0] I3ae9dbf37dbadabaf8a56188eae40288, If9b05209071a1c16ecce1c28f886ee1d;
reg [fgallag_WDTH -1:0] Iae4d59e569911a81bb653cdb58c65137, Iebb87060282934e67cd1e7e8493fcf20;
reg [fgallag_WDTH -1:0] I9b12cb33d0f37813bd735c14d8be517e, I22b235f6e6f0938fe2a026f91bfd72cf;
reg [fgallag_WDTH -1:0] Ifab01268c2a1f0385dc4b18a9d488321, I185299c78eca06f6174996089a2df4d5;
reg [fgallag_WDTH -1:0] Ie0f0a8cf008e6a10d1698c11c380df97, I90f70f8385f7d8fc69fe21f42d96eeeb;
reg [fgallag_WDTH -1:0] I99aa62ad841c5bd5b1f2b6758d046784, I5d03a9d2e8ca426a10005cf5a1689f4f;
reg [fgallag_WDTH -1:0] I3fc64e5c431cd64d48f3cc5c9c86f342, I1f30e3cf906aa5a09d71f23c5be461ba;
reg [fgallag_WDTH -1:0] I65a139ae2fa69f57c3a8ed35e00e29ae, I13069dca0bc85e00a513e9fe7562b346;
reg [fgallag_WDTH -1:0] I628bc7c30b5e896c2b8f4af752b44637, Ib69a5ff88f694a3cf18fa11fcccdd9c2;
reg [fgallag_WDTH -1:0] I5c7ed27126a8097481ab5f966867783b, If4b3a419df7ce8b8cd5f2b7a26e1a629;
reg [fgallag_WDTH -1:0] I686481757183441e45d85fece1a7b514, I03b2bc96c0edf4f4c27ab02d8beda293;
reg [fgallag_WDTH -1:0] I10929316643f6670bedc63e77b293c97, Iddd38c69253e1ba79f6762c9e69857ad;
reg [fgallag_WDTH -1:0] Ia66d818d01365175f416a4de87a281bb, I3437ae400dbe3a2eb99a65a263889bb6;
reg [fgallag_WDTH -1:0] I7711386635a1760e7976d0947e0a5f8a, I0bb76633859552dc99f63b3c520037cc;
reg [fgallag_WDTH -1:0] I4b2cc8ae58d2fb89bd9095b2bb688cbe, Ifcb79d8780c0e5859fc885521a3a4070;
reg [fgallag_WDTH -1:0] Ied1035a697824a18281435fe2b7f1f56, Ia43aac10d65d1661b3d7f9968c829c21;
reg [fgallag_WDTH -1:0] I3e9ecaf8da044766c57685a1065ce10a, I6ecfb2be423754892a663315c2c74440;
reg [fgallag_WDTH -1:0] Ibebda2f9816088ea15cd5b4f555c5d33, Ic9b31062ba9aedcda0f4c91e39fe1814;
reg [fgallag_WDTH -1:0] I6043631f93e2c514d5ed6e86beffa7c6, Ie5ff9375515964757ffe821812ed8e73;
reg [fgallag_WDTH -1:0] Ibc084904fb63bb24102789357ce2cd76, I5152ee18b04c8d038ead4817bc68fa57;
reg [fgallag_WDTH -1:0] I9e82413dca68de150b81bd27ab180980, I606544d89b457531a204f0a9a061dc74;
reg [fgallag_WDTH -1:0] I4992c306a07d2e104a72dfcc37968e8c, If7bcb8673722495218ae395b5716c89a;
reg [fgallag_WDTH -1:0] I637c0445b26879a0fb9d7d94baef55e4, I755d5c8837cace07fc3c0393a6ba2a43;
reg [fgallag_WDTH -1:0] I3f1f9cecc45287a2c9487c04d8430b5b, I2051dc0ec4b2e1de6e3308c6e0ae74bd;
reg [fgallag_WDTH -1:0] Ife3d2f48786c2e11f7c4f8b4a7bb829e, I9ff8a14d8788f2e0deb7a0c1f4d0fa0d;
reg [fgallag_WDTH -1:0] I0a019e2861b41f395bd12b43cd978e59, Id017562a43e853ec27712b3f8d449361;
reg [fgallag_WDTH -1:0] I34fcd098fa2b426f98542121dae204fc, I7c408398d6b1e91c00962636fbf59b83;
reg [fgallag_WDTH -1:0] I8c9a0911720c403f2794fa5662a31207, I53387cf352304840ccae53d5b5b153e7;
reg [fgallag_WDTH -1:0] I11af377ea2ae07f2249042a6daeef846, I6d483d27683d84d2309d756d36f43ae9;
reg [fgallag_WDTH -1:0] Ib5d6d77cf92f29c1b498252859ec19ff, I1c44630f8f2d9bf2a5df81f22a67ed43;
reg [fgallag_WDTH -1:0] I1d6100bd00e7e46af792dd99286391a5, Ic7a0ea4cb5954db181b37e8072cf54fb;
reg [fgallag_WDTH -1:0] Ia6e85ec8c498ed70cb4a4e01bf8d1530, I591e5713ec07915309f4a588ea51a990;
reg [fgallag_WDTH -1:0] Icc6d40c383e5580bbac65b6c77da6528, Ibab6e2a97bd19438998b97780bdae17d;
reg [fgallag_WDTH -1:0] Id939e83f81205a66485908e0bba8504d, Icb868f4e4f276036478f3977e8d831a3;
reg [fgallag_WDTH -1:0] Ie709765eec241ae95c588fbfed18a87e, I8dde06b1ca763ca0cdd273e440de86ab;
reg [fgallag_WDTH -1:0] I497fb247a6572f689aea3e595e657fdb, I44049fcab453cba240bed48d89a664e5;
reg [fgallag_WDTH -1:0] I659b78a601b47941441dc1debcae4d46, I4c6d3af7a2d1adb1f60b61a523dd9bff;
reg [fgallag_WDTH -1:0] Ibed2d1ab1707ca759a8b09a5147a4268, I70d83e5081cd2c9051f9c6b8652462d7;
reg [fgallag_WDTH -1:0] I23c058e418bad060fb1404b248782705, Id841c70607e96ab5144c91a573a771c7;
reg [fgallag_WDTH -1:0] I95f73f2e7a5268d25f4fcaa53339c2fc, Ib9318ad9f3aa8b5fd8b8c59fe3bd1616;
reg [fgallag_WDTH -1:0] I90b927c01ca8d69239141958db410c54, I569eefbb2dbaf1e589f1cf1bc35721c7;
reg [fgallag_WDTH -1:0] I79c64b98cdd4f4a1b41ddd2480c5d62a, Id399e2be28090c81e93743f1bfe00347;
reg [fgallag_WDTH -1:0] I76071439d501dfac67b1355c33f04c79, I04b7604f3936be2c49deb140a0d1eae5;
reg [fgallag_WDTH -1:0] I3bed56f31105c1dd5524f2e04a6cdc0f, I23d474402240b1761c2f9d785cd2973b;
reg [fgallag_WDTH -1:0] I1ca06bac6a4d082efeed13d0448630fb, Ia5bbbcb8956d08a529457d6ca2c38ebc;
reg [fgallag_WDTH -1:0] Iefd7ba660203932e953d509b10032e4d, I116f8968c4a02e2a22a8ea4eb5dd3951;
reg [fgallag_WDTH -1:0] I76b3bd4ded426c469b208f83f7bb1781, I1ebdf4675d0986c912c52af538ac358d;
reg [fgallag_WDTH -1:0] I36261da4cc2946a22e80fb6f2a394753, I92cd919b7b5b4ca8984668bfbdb43d3b;
reg [fgallag_WDTH -1:0] Iaa84b434bf0040f25a2dd6af77d90df4, Ibdecc8406ba4102713fde4a51206403f;
reg [fgallag_WDTH -1:0] I1a314b0ac2b2897b23d2e9fd3e5e63f0, Ie79b340519a003c4388b90a3d8fac445;
reg [fgallag_WDTH -1:0] I64eff7490d835e24cf4e5f4d0c60e18e, I719e56962c59071b4783ff87e554a37e;
reg [fgallag_WDTH -1:0] I95c886a9726c33f2a8f2f9413c9486cb, Id2a6a7580c31d450f8c78217e8997f7e;
reg [fgallag_WDTH -1:0] Ie2fbf1593b8aa394377ccc4ef0f705b6, I74f0171925c0986fe140602b09a0caf2;
reg [fgallag_WDTH -1:0] I124a5e6d2c3103fbb4699cc2f7528a48, I5e9bef3789fd851fb793bea78beef829;
reg [fgallag_WDTH -1:0] I3625276282d727c6510f5123ee467e73, I0f3062a73289917dc123b87666bdad07;
reg [fgallag_WDTH -1:0] I771e25faed091d437e00dae0e66d088b, I238a8e826a1d8f069455ae0163d508f2;
reg [fgallag_WDTH -1:0] Iad7a84f48832522261c3495844b19dde, Iedd0e164003fd9532945df51a5408307;
reg [fgallag_WDTH -1:0] I8de675a8e37ed2b30a82e49ff6d510a0, Ib8a70644d197140114eacd4c9612dd77;
reg [fgallag_WDTH -1:0] I4bbc70e0a3a56eeb62af73e6c80006b4, Ib171958fe2af1d20130ca83b668af768;
reg [fgallag_WDTH -1:0] I5c97bebf3cd2472e43ae7312d3956bb5, I80d67b47c44a3b424d1ed4c8e357c265;
reg [fgallag_WDTH -1:0] I527847fbb55900e97761446b030ed540, Iaa9183f11cd736e6271b9e6259a807a7;
reg [fgallag_WDTH -1:0] Ie707c8b057532a88aff15ca43d1a4cef, I1f2ac0b753cee68f5e984de8994f2f0d;
reg [fgallag_WDTH -1:0] I41708d131f34ee41b74f571661e751c6, I495ac3abe6643625add1aeef4776b39e;
reg [fgallag_WDTH -1:0] I410af2866a81357ed84738c1800ee8e2, I4c8185fc93a069b6fa81b3936de2b4b0;
reg [fgallag_WDTH -1:0] Iae78b53a85d3b3441bb251688c85fe66, Ib05eddf67c2a5797e8e0e733fca4328b;
reg [fgallag_WDTH -1:0] I1c4646eab74db4876187e2e87d861e4d, I8f8316a85f64267a15f99a0b47db5f08;
reg [fgallag_WDTH -1:0] Idb04b139376a9fd83c6f921b02c31849, I69116a38d209590270e61cfe9d2e56d5;
reg [fgallag_WDTH -1:0] I64c0c3c0d18d18ed62b2b2910930f8a0, I713819fe0cf6d54393d9cd5a32a37807;
reg [fgallag_WDTH -1:0] I0c622446a77fe077062fd87448e11fec, I811d183d31135919e65f87250c0ba456;
reg [fgallag_WDTH -1:0] Ie69cbbb6131f04ccf84db28990b4dbdd, I8a99662ff2d2b8f153d6d9359b88eff5;
reg [fgallag_WDTH -1:0] Id0b467dbeaa2b30126ed60489530e29f, Ib246205f26dd43b9d1fa057a2179e4b2;
reg [fgallag_WDTH -1:0] Idac7b0bec594eccd74ac2d944da4484e, I972077c6595b44e3113b0d7a925aa913;
reg [fgallag_WDTH -1:0] I4ddb027f246fb2b145bba7b01687d39b, Idde043a5721004c3904eb2b55031e7c1;
reg [fgallag_WDTH -1:0] I754ff7341b379de55d5facc6fcc9f874, Iebfd00d9a2a6e39e6fc73f95c4f29539;
reg [fgallag_WDTH -1:0] Ia7a71696b5ebed6c80cafb33a031626e, I3e10f0cc7d257acf63a5ca7a0cb9c7cf;
reg [fgallag_WDTH -1:0] I542db58e949d7d1c542c075005fb065c, I62895b1265f950882fc5fb770dafd51d;
reg [fgallag_WDTH -1:0] I28aaa9370cb22a81b7c8d20fe7e1d347, I9f890d3f6b5edfbf106d59df07cb1b68;
reg [fgallag_WDTH -1:0] If4abfdcd468d4d98db5f32bb99303035, Icd6b85be80234c06eaeaf1347ebabb38;
reg [fgallag_WDTH -1:0] Idfc14e592719d57828f8e6dc2130e270, I1e9047545567e723fa101ab94dffa45f;
reg [fgallag_WDTH -1:0] Ia51b4598ba3f6c128ffcd421a3ba7309, Iea7a223f22fb02e29871f500b61fa205;
reg [fgallag_WDTH -1:0] Iee935e25f9fe5c7844bb0c0490cbb90f, Ida8637c3dd298410093697077abad3e0;
reg [fgallag_WDTH -1:0] I05d0b3631f8501ecafcbb321c15be5f1, Ic767ff5ab4bfc377cf1b7bae10b42d3e;
reg [fgallag_WDTH -1:0] I7ea9adf8dba141eef7a08d76105580ec, Ieafe43b66027e5b192cdd5fe25977f4c;
reg [fgallag_WDTH -1:0] Ifa4cd939b137dc050f675a493546ddf6, I41d92f30c38301789ac4155986c2a634;
reg [fgallag_WDTH -1:0] I7a6215a05dd8dbdcb421d7df535c5b67, I5c4bedc45aa3faab29c3547e29c6db68;
reg [fgallag_WDTH -1:0] Ibd0c06d4190a37b90c51d562c6019551, I1bf648fa37015e2997a689769881149c;
reg [fgallag_WDTH -1:0] I75b4b57cf9d7400feec38e037c948352, I4f38b0092062a40f0bd68bbe8911f248;
reg [fgallag_WDTH -1:0] I14a4e51be5aa98fa28cc4740e6446747, I74c408ce157c47049698b52949d1fd38;
reg [fgallag_WDTH -1:0] I43196769a96d15dd03318e43b48a6b4d, I3ed597f1774bf9274566cb5fc7dbbdc5;
reg [fgallag_WDTH -1:0] I8494b9c75594140fabc1158bacf4438a, I8d111345e29debfc7addbb913d4e9054;
reg [fgallag_WDTH -1:0] I931bf44a358d9fd91d31aa78d3e16312, I8d19b379f6693601f18ea748bbbadf9b;
reg [fgallag_WDTH -1:0] I5355f3939098f1ae0aa0f254b8e7e163, I68521e797f1f404e6a190855b1a322f1;
reg [fgallag_WDTH -1:0] I6228ab1c737aec5845684c0eff41dac4, I5ecffa51c73d64359ba32c2cf56c6b7a;
reg [fgallag_WDTH -1:0] I9034255c2128aa8c4d707bf003a57e86, I2adb86feb263103c1419d34eb9b8ae4e;
reg [fgallag_WDTH -1:0] Ia9bc32f3ef4f4681782fec452e572cf2, I733561ae7e5600d8275667457f2ea151;
reg [fgallag_WDTH -1:0] I9791a65b490a63c3c201409a30b86199, I4db74afe0a9f15f643d8295051f762c0;
reg [fgallag_WDTH -1:0] Id5297cb2f91d5b3e67c4bd97a8c05401, Id194460b74adf4856635d5c432ea772f;
reg [fgallag_WDTH -1:0] Ibc826b606b10904061b2666eb204469e, Ifc1dfcb0afd77d1a01bbb54da77a5f70;
reg [fgallag_WDTH -1:0] I06dabbc9dc6fb6b8fa517e188ee74208, I0cec4bb6f8f736beea5fd2dc57310432;
reg [fgallag_WDTH -1:0] I4d3607d7cd13b86ae4a22bebaf65ef0e, If878a4e87d963261e36cde448d6c3bbc;
reg [fgallag_WDTH -1:0] Ia974eebd7b7563b2f0822f538c13a911, I2d28d468beee8a809ece79a2b7b07d27;
reg [fgallag_WDTH -1:0] I191470ccfa2c2838a34aceb571582bb4, I8b553bf742d14f23835e62aeade33413;
reg [fgallag_WDTH -1:0] I01714219c84cfbfd7ff940108ddbb6b3, Iacc099c63faabe7dda342eafe07e26d4;
reg [fgallag_WDTH -1:0] I118d11a015af5944d64290a46bf49c09, Ifc3d28213bc38fbcff2eb42ebc350c8a;
reg [fgallag_WDTH -1:0] Ib878ef5592b0bf1af247ede54fe13a45, I7fd466826e266237c64dd4010bf19ed8;
reg [fgallag_WDTH -1:0] I7686f623f51c5a9f8f3f8d143ed8bcb5, I5c42c7a5b8b8d73e5374eb00cf80f91b;
reg [fgallag_WDTH -1:0] I4d48fc8081756af036b8f1b1b9e56051, I2e4f341a2f112ba1df12c82183bd3566;
reg [fgallag_WDTH -1:0] Ia1d93d4bbc6b1e73dbb0c6c26d102f10, I757c6c719d8455faea81fa0901a2c15e;
reg [fgallag_WDTH -1:0] Ifb7d0d12a916fc3f2f9c0341f27ef53f, Ie146524ab065ed90500947d0e77f7e5e;
reg [fgallag_WDTH -1:0] I4ee596c96f91a18ef1ebb0ee6de285ae, I40fd0db59f8b8877f3f62b9b87e2892d;
reg [fgallag_WDTH -1:0] I5aeda0b5dc8459d86e9ab5082bf9fed8, I2c05c52719e300f911b6245928a40fb3;
reg [fgallag_WDTH -1:0] I7b6ff145fa076d152af672e0c3a062bc, I07acde143b8be8c4ec4e562a66562b58;
reg [fgallag_WDTH -1:0] I3929cfb9fb8795d4dd9f54f9c4a2fa02, I5d0ae3e1a3333e7dcc389a609644376a;
reg [fgallag_WDTH -1:0] If33f043047ad17b323733a201aa649da, I13b47a7b710051dde6ab5cae17f216d4;
reg [fgallag_WDTH -1:0] Icfb9314b47604c3b065ffdd5d9042682, I1c0174a95fd6b5322576907671acdd82;
reg [fgallag_WDTH -1:0] I5cd61f07b490ca79f1ec069ed2d47528, Ica09fab419a2bd1a966956988b6507b3;
reg [fgallag_WDTH -1:0] I1bace448ce54ae41e9e8d27acf548338, I27097218191d9ad8cd380a75b5b4d467;
reg [fgallag_WDTH -1:0] I692bf3f934f0ee8fbf02c7dce98f924c, I354ec2d3605e41d982076dcb7e32d2c1;
reg [fgallag_WDTH -1:0] Ifb3af535b42775dae1e0ade2d8bf79df, I14c93bdff35500174e3db5c18b48cb94;
reg [fgallag_WDTH -1:0] I569a621522dd636df609f60c1b22d7f7, I30084765c13a4c6a7514a16e3f45a9c2;
reg [fgallag_WDTH -1:0] Ic651187a36eb89eaf129a368af3474ee, I1f07b4c82c226595be454e07eed346ab;
reg [fgallag_WDTH -1:0] Ib120bd9cfec97e7956bb64f8e4527caf, I7401e0464789f88be2b661eb055bbdef;
reg [fgallag_WDTH -1:0] I41e452eee26c8ede812d3ca957488aec, Ia1e603a00bf98ee21caea749765ed341;
reg I7aa491e6301b27435c2dadebe447b43a ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 Ia6f93d7eab83c88b604f8a81a74c04e9 <= 'h0;
 Ice05aa8a4d2a062da9785286081fd024 <= 'h0;
 I6e41efdbe6eeb41b9c9b39e56f3d8b9c <= 'h0;
 Ibe53a3b8a9caa8643361263d463290c8 <= 'h0;
 Ifbcddebb5f791d2df0b2e7aa94a81c22 <= 'h0;
 I341146b894d9d94c2c803e6b6c464085 <= 'h0;
 Iccfcaba2f6129c8201cb97323a8e740a <= 'h0;
 I850f7b404a1ab022498350d9ef0cbdc2 <= 'h0;
 Ie88f3ca2bc79208be9385225a7ad7268 <= 'h0;
 If4137d66b193970e9ae89b8e1b00e8ca <= 'h0;
 I877047b00cef1f6a938ed9915215e203 <= 'h0;
 Ic9e529e5e428a666bf6bcf2041969d1e <= 'h0;
 I2e8ce46a773bcf5f2c3129441a267af4 <= 'h0;
 Ie734c46bfea46055c73a2642b3f8a7da <= 'h0;
 Id980a518f6b9c84062f5bd7d6f57472f <= 'h0;
 I8901003e5fb9f89fddb0fa87dc5b2d05 <= 'h0;
 Ia5402393b456807ca5fee0ecb219c7d9 <= 'h0;
 I41d38680c5aca0364ef9c716cd4525e7 <= 'h0;
 I03ee8c787b49b08c0a5a503bd28fcca5 <= 'h0;
 Id85bac587e9c200406f0aecafbaf3dd5 <= 'h0;
 Ibb5dbc2fc80aca18dbaa13b7ecdb6c20 <= 'h0;
 I9b5df9c23c9a2aaa14a99abd110075cb <= 'h0;
 Ic00f5a4dfdbbf58316107417ccc6bb74 <= 'h0;
 Ic208118fb71fea311016edcb1203407d <= 'h0;
 Ib3d96f215fc42ace8fddda8c64afbc05 <= 'h0;
 Ie304d02670ae74fb93fb42328d43079e <= 'h0;
 I1a875fdb7e3681839eeb5fdb8c6b47c3 <= 'h0;
 I85c6964245f5e3423ddfcae7ae864429 <= 'h0;
 Idd3396a16fde9c928bfd71f9b05b98bf <= 'h0;
 I3a124ec3bd01d433c39ecbfd0b153d74 <= 'h0;
 I7be57c1f60b38d43d0fe2c02175aeef5 <= 'h0;
 I886a56b1cae34e1860e4cd2c28606a45 <= 'h0;
 I4dfc6b1e7b358ad6a32f6682e487d962 <= 'h0;
 I4c60daf9c53a50f2a228ca9ad0d75115 <= 'h0;
 I5fa487af5385cb6dcd0bac274a2b2261 <= 'h0;
 If3024e217350078f9a06275cc31b6699 <= 'h0;
 Ifb39ced2cc4424e46be38af68161181a <= 'h0;
 I17934cad1385024244ce8bd07b709db0 <= 'h0;
 Ie43b90c9bb7dcb76f116c75615df246b <= 'h0;
 I7f095ecd42b65b1781e2290db664a73d <= 'h0;
 I4d7c79dc1c72745d5750cac86454beb8 <= 'h0;
 I00c66baa19546590a542100f8883d4ab <= 'h0;
 I97293ec9139e6e252c554d9f26619f06 <= 'h0;
 I067a46089f564be32860d44b3c69af1a <= 'h0;
 Ib11764f9c254c7ddf0782d0cccae0067 <= 'h0;
 Ic63385ac292f30c59ab2ad6f8b7d8903 <= 'h0;
 I5d3f02e43c3a9ab32c9769c1cf45ec6c <= 'h0;
 I968edb5f5a70a3d391db21db00dafe78 <= 'h0;
 I59ad05479adc69422b7e06e4507a8f7a <= 'h0;
 I3755b61b6fb958538b1b906a4ad1103d <= 'h0;
 I0ba5990e179758e1080a8407412a9a59 <= 'h0;
 I7562a62ae85c4676605b60594722a950 <= 'h0;
 I62c2ba2ded74107adfcbe43670718e65 <= 'h0;
 Ie43871350b062263474a7e0dbca850ce <= 'h0;
 I12d1f6ac4ef39cb76907b09745b4f8ad <= 'h0;
 If9b05209071a1c16ecce1c28f886ee1d <= 'h0;
 Iebb87060282934e67cd1e7e8493fcf20 <= 'h0;
 I22b235f6e6f0938fe2a026f91bfd72cf <= 'h0;
 I185299c78eca06f6174996089a2df4d5 <= 'h0;
 I90f70f8385f7d8fc69fe21f42d96eeeb <= 'h0;
 I5d03a9d2e8ca426a10005cf5a1689f4f <= 'h0;
 I1f30e3cf906aa5a09d71f23c5be461ba <= 'h0;
 I13069dca0bc85e00a513e9fe7562b346 <= 'h0;
 Ib69a5ff88f694a3cf18fa11fcccdd9c2 <= 'h0;
 If4b3a419df7ce8b8cd5f2b7a26e1a629 <= 'h0;
 I03b2bc96c0edf4f4c27ab02d8beda293 <= 'h0;
 Iddd38c69253e1ba79f6762c9e69857ad <= 'h0;
 I3437ae400dbe3a2eb99a65a263889bb6 <= 'h0;
 I0bb76633859552dc99f63b3c520037cc <= 'h0;
 Ifcb79d8780c0e5859fc885521a3a4070 <= 'h0;
 Ia43aac10d65d1661b3d7f9968c829c21 <= 'h0;
 I6ecfb2be423754892a663315c2c74440 <= 'h0;
 Ic9b31062ba9aedcda0f4c91e39fe1814 <= 'h0;
 Ie5ff9375515964757ffe821812ed8e73 <= 'h0;
 I5152ee18b04c8d038ead4817bc68fa57 <= 'h0;
 I606544d89b457531a204f0a9a061dc74 <= 'h0;
 If7bcb8673722495218ae395b5716c89a <= 'h0;
 I755d5c8837cace07fc3c0393a6ba2a43 <= 'h0;
 I2051dc0ec4b2e1de6e3308c6e0ae74bd <= 'h0;
 I9ff8a14d8788f2e0deb7a0c1f4d0fa0d <= 'h0;
 Id017562a43e853ec27712b3f8d449361 <= 'h0;
 I7c408398d6b1e91c00962636fbf59b83 <= 'h0;
 I53387cf352304840ccae53d5b5b153e7 <= 'h0;
 I6d483d27683d84d2309d756d36f43ae9 <= 'h0;
 I1c44630f8f2d9bf2a5df81f22a67ed43 <= 'h0;
 Ic7a0ea4cb5954db181b37e8072cf54fb <= 'h0;
 I591e5713ec07915309f4a588ea51a990 <= 'h0;
 Ibab6e2a97bd19438998b97780bdae17d <= 'h0;
 Icb868f4e4f276036478f3977e8d831a3 <= 'h0;
 I8dde06b1ca763ca0cdd273e440de86ab <= 'h0;
 I44049fcab453cba240bed48d89a664e5 <= 'h0;
 I4c6d3af7a2d1adb1f60b61a523dd9bff <= 'h0;
 I70d83e5081cd2c9051f9c6b8652462d7 <= 'h0;
 Id841c70607e96ab5144c91a573a771c7 <= 'h0;
 Ib9318ad9f3aa8b5fd8b8c59fe3bd1616 <= 'h0;
 I569eefbb2dbaf1e589f1cf1bc35721c7 <= 'h0;
 Id399e2be28090c81e93743f1bfe00347 <= 'h0;
 I04b7604f3936be2c49deb140a0d1eae5 <= 'h0;
 I23d474402240b1761c2f9d785cd2973b <= 'h0;
 Ia5bbbcb8956d08a529457d6ca2c38ebc <= 'h0;
 I116f8968c4a02e2a22a8ea4eb5dd3951 <= 'h0;
 I1ebdf4675d0986c912c52af538ac358d <= 'h0;
 I92cd919b7b5b4ca8984668bfbdb43d3b <= 'h0;
 Ibdecc8406ba4102713fde4a51206403f <= 'h0;
 Ie79b340519a003c4388b90a3d8fac445 <= 'h0;
 I719e56962c59071b4783ff87e554a37e <= 'h0;
 Id2a6a7580c31d450f8c78217e8997f7e <= 'h0;
 I74f0171925c0986fe140602b09a0caf2 <= 'h0;
 I5e9bef3789fd851fb793bea78beef829 <= 'h0;
 I0f3062a73289917dc123b87666bdad07 <= 'h0;
 I238a8e826a1d8f069455ae0163d508f2 <= 'h0;
 Iedd0e164003fd9532945df51a5408307 <= 'h0;
 Ib8a70644d197140114eacd4c9612dd77 <= 'h0;
 Ib171958fe2af1d20130ca83b668af768 <= 'h0;
 I80d67b47c44a3b424d1ed4c8e357c265 <= 'h0;
 Iaa9183f11cd736e6271b9e6259a807a7 <= 'h0;
 I1f2ac0b753cee68f5e984de8994f2f0d <= 'h0;
 I495ac3abe6643625add1aeef4776b39e <= 'h0;
 I4c8185fc93a069b6fa81b3936de2b4b0 <= 'h0;
 Ib05eddf67c2a5797e8e0e733fca4328b <= 'h0;
 I8f8316a85f64267a15f99a0b47db5f08 <= 'h0;
 I69116a38d209590270e61cfe9d2e56d5 <= 'h0;
 I713819fe0cf6d54393d9cd5a32a37807 <= 'h0;
 I811d183d31135919e65f87250c0ba456 <= 'h0;
 I8a99662ff2d2b8f153d6d9359b88eff5 <= 'h0;
 Ib246205f26dd43b9d1fa057a2179e4b2 <= 'h0;
 I972077c6595b44e3113b0d7a925aa913 <= 'h0;
 Idde043a5721004c3904eb2b55031e7c1 <= 'h0;
 Iebfd00d9a2a6e39e6fc73f95c4f29539 <= 'h0;
 I3e10f0cc7d257acf63a5ca7a0cb9c7cf <= 'h0;
 I62895b1265f950882fc5fb770dafd51d <= 'h0;
 I9f890d3f6b5edfbf106d59df07cb1b68 <= 'h0;
 Icd6b85be80234c06eaeaf1347ebabb38 <= 'h0;
 I1e9047545567e723fa101ab94dffa45f <= 'h0;
 Iea7a223f22fb02e29871f500b61fa205 <= 'h0;
 Ida8637c3dd298410093697077abad3e0 <= 'h0;
 Ic767ff5ab4bfc377cf1b7bae10b42d3e <= 'h0;
 Ieafe43b66027e5b192cdd5fe25977f4c <= 'h0;
 I41d92f30c38301789ac4155986c2a634 <= 'h0;
 I5c4bedc45aa3faab29c3547e29c6db68 <= 'h0;
 I1bf648fa37015e2997a689769881149c <= 'h0;
 I4f38b0092062a40f0bd68bbe8911f248 <= 'h0;
 I74c408ce157c47049698b52949d1fd38 <= 'h0;
 I3ed597f1774bf9274566cb5fc7dbbdc5 <= 'h0;
 I8d111345e29debfc7addbb913d4e9054 <= 'h0;
 I8d19b379f6693601f18ea748bbbadf9b <= 'h0;
 I68521e797f1f404e6a190855b1a322f1 <= 'h0;
 I5ecffa51c73d64359ba32c2cf56c6b7a <= 'h0;
 I2adb86feb263103c1419d34eb9b8ae4e <= 'h0;
 I733561ae7e5600d8275667457f2ea151 <= 'h0;
 I4db74afe0a9f15f643d8295051f762c0 <= 'h0;
 Id194460b74adf4856635d5c432ea772f <= 'h0;
 Ifc1dfcb0afd77d1a01bbb54da77a5f70 <= 'h0;
 I0cec4bb6f8f736beea5fd2dc57310432 <= 'h0;
 If878a4e87d963261e36cde448d6c3bbc <= 'h0;
 I2d28d468beee8a809ece79a2b7b07d27 <= 'h0;
 I8b553bf742d14f23835e62aeade33413 <= 'h0;
 Iacc099c63faabe7dda342eafe07e26d4 <= 'h0;
 Ifc3d28213bc38fbcff2eb42ebc350c8a <= 'h0;
 I7fd466826e266237c64dd4010bf19ed8 <= 'h0;
 I5c42c7a5b8b8d73e5374eb00cf80f91b <= 'h0;
 I2e4f341a2f112ba1df12c82183bd3566 <= 'h0;
 I757c6c719d8455faea81fa0901a2c15e <= 'h0;
 Ie146524ab065ed90500947d0e77f7e5e <= 'h0;
 I40fd0db59f8b8877f3f62b9b87e2892d <= 'h0;
 I2c05c52719e300f911b6245928a40fb3 <= 'h0;
 I07acde143b8be8c4ec4e562a66562b58 <= 'h0;
 I5d0ae3e1a3333e7dcc389a609644376a <= 'h0;
 I13b47a7b710051dde6ab5cae17f216d4 <= 'h0;
 I1c0174a95fd6b5322576907671acdd82 <= 'h0;
 Ica09fab419a2bd1a966956988b6507b3 <= 'h0;
 I27097218191d9ad8cd380a75b5b4d467 <= 'h0;
 I354ec2d3605e41d982076dcb7e32d2c1 <= 'h0;
 I14c93bdff35500174e3db5c18b48cb94 <= 'h0;
 I30084765c13a4c6a7514a16e3f45a9c2 <= 'h0;
 I1f07b4c82c226595be454e07eed346ab <= 'h0;
 I7401e0464789f88be2b661eb055bbdef <= 'h0;
 Ia1e603a00bf98ee21caea749765ed341 <= 'h0;
 I7aa491e6301b27435c2dadebe447b43a <= 'h0;
end
else
begin
 Ia6f93d7eab83c88b604f8a81a74c04e9 <=  I9c9ab24ecd80ca61b89534e3e5adfca8;
 Ice05aa8a4d2a062da9785286081fd024 <=  Ie92d645c17dda47f594bc34b0937caac;
 I6e41efdbe6eeb41b9c9b39e56f3d8b9c <=  Ieb8b25a5f6d3cc4cead3f3845234d1d3;
 Ibe53a3b8a9caa8643361263d463290c8 <=  Ibcbdbe8034a373448800d1b745cb5849;
 Ifbcddebb5f791d2df0b2e7aa94a81c22 <=  Ibd0769c69670150d8263d9873cbf668f;
 I341146b894d9d94c2c803e6b6c464085 <=  I2010cff1e77f9706d8c659482f51c898;
 Iccfcaba2f6129c8201cb97323a8e740a <=  I4183447a1a1727e91b0fcabb9bec1963;
 I850f7b404a1ab022498350d9ef0cbdc2 <=  I780bea956f609c6f3cd0ffd126f99316;
 Ie88f3ca2bc79208be9385225a7ad7268 <=  I349cff38817dd1607e798b9a2ae6fb8b;
 If4137d66b193970e9ae89b8e1b00e8ca <=  I3ff605a8af8eceb2c055e842e6208958;
 I877047b00cef1f6a938ed9915215e203 <=  Ib53b2b0d39dbe6d09f51e0af27e5986f;
 Ic9e529e5e428a666bf6bcf2041969d1e <=  I343242367c13febc05ee63f57dd4f754;
 I2e8ce46a773bcf5f2c3129441a267af4 <=  Ibde6749f31c571c5209a8b36c1c8f4da;
 Ie734c46bfea46055c73a2642b3f8a7da <=  Ib735324969bc744cc0ab8c2b3a7c5561;
 Id980a518f6b9c84062f5bd7d6f57472f <=  If53ed28774233bca87090e799465e3a5;
 I8901003e5fb9f89fddb0fa87dc5b2d05 <=  Ib5017be08e079fe946c365fc01461d11;
 Ia5402393b456807ca5fee0ecb219c7d9 <=  I0f24b1ca1d272d4971cde83a2acfe5ac;
 I41d38680c5aca0364ef9c716cd4525e7 <=  I1d1f2f5dd46b3f89c5a614ebad298d13;
 I03ee8c787b49b08c0a5a503bd28fcca5 <=  I09dbcf2140141aaa400ad52408f8ab41;
 Id85bac587e9c200406f0aecafbaf3dd5 <=  I8315726dd19b5074a78796ee704d7108;
 Ibb5dbc2fc80aca18dbaa13b7ecdb6c20 <=  Idb03654ee570200d2fe82907af7095d7;
 I9b5df9c23c9a2aaa14a99abd110075cb <=  I9a5f25915425b586c1c3979240ff1a54;
 Ic00f5a4dfdbbf58316107417ccc6bb74 <=  I259241ceeda0568e6c10162cd43ca1dc;
 Ic208118fb71fea311016edcb1203407d <=  I66d1b07d77d2fe21d535920b30e176ff;
 Ib3d96f215fc42ace8fddda8c64afbc05 <=  I135dcccb8e63f697fe4559b964322345;
 Ie304d02670ae74fb93fb42328d43079e <=  Ic37c4058485edfc0ca4f12fd7a97bf93;
 I1a875fdb7e3681839eeb5fdb8c6b47c3 <=  I1400488e51bbe6c921439713342d39f8;
 I85c6964245f5e3423ddfcae7ae864429 <=  Iaa8359974e7a41f754b38d6a232c5e72;
 Idd3396a16fde9c928bfd71f9b05b98bf <=  Ie99b9c10b4b5208374b9f4ba1bd3eeab;
 I3a124ec3bd01d433c39ecbfd0b153d74 <=  I54462091230adebf4bf4ec0cea25e374;
 I7be57c1f60b38d43d0fe2c02175aeef5 <=  Iba9e737dd791a2ee966dbf6958339d65;
 I886a56b1cae34e1860e4cd2c28606a45 <=  Ib205f5f9a6005baa465f1b254e4014d0;
 I4dfc6b1e7b358ad6a32f6682e487d962 <=  I5ea13e282884d2343e8fdbe17d7ee058;
 I4c60daf9c53a50f2a228ca9ad0d75115 <=  I6d8ed091d5f44b3b49e8b0eb63f0d106;
 I5fa487af5385cb6dcd0bac274a2b2261 <=  I4109473d968250506e17f8227bc55d06;
 If3024e217350078f9a06275cc31b6699 <=  Ia7da78b0d37028fcd34d3d39c7e36596;
 Ifb39ced2cc4424e46be38af68161181a <=  I034454a1608fbde69fffb6b28e685f9f;
 I17934cad1385024244ce8bd07b709db0 <=  I6e487d671a19855fd1eae42664d9c57f;
 Ie43b90c9bb7dcb76f116c75615df246b <=  Ib49b6b6895bd7200dc9e026584bea017;
 I7f095ecd42b65b1781e2290db664a73d <=  I220ce4284bf6adf0e46cf524b04a0e1b;
 I4d7c79dc1c72745d5750cac86454beb8 <=  I64586e3b7241a57c2e887b651819c7f9;
 I00c66baa19546590a542100f8883d4ab <=  Ifad0bf7a3d7d334b5f8ea0d1a973fd39;
 I97293ec9139e6e252c554d9f26619f06 <=  If060b99963382d16c1f779faf00a7128;
 I067a46089f564be32860d44b3c69af1a <=  Ie80ad5b1c3c4046c80e6cb96ee51e5c0;
 Ib11764f9c254c7ddf0782d0cccae0067 <=  I4fe400daeacdfbebafcdf7e753af2787;
 Ic63385ac292f30c59ab2ad6f8b7d8903 <=  I5c1ec1001d1ea61ab7198336742ed99d;
 I5d3f02e43c3a9ab32c9769c1cf45ec6c <=  If50cfdca6c9b8000665da2513244ff24;
 I968edb5f5a70a3d391db21db00dafe78 <=  I4367feaf57687befa18bc6a902573bb9;
 I59ad05479adc69422b7e06e4507a8f7a <=  I8f2820928683d8d88d41b80a9d9832dd;
 I3755b61b6fb958538b1b906a4ad1103d <=  Id980002a738b3ab2a4c2ccb9d232d141;
 I0ba5990e179758e1080a8407412a9a59 <=  Ib1db1798d076dc0a6fa322c47e0ac062;
 I7562a62ae85c4676605b60594722a950 <=  Iba73f7b76a2e16d7d84cfbab4473143d;
 I62c2ba2ded74107adfcbe43670718e65 <=  Iad0a6e20283bbf4bd4114a0c70c0685e;
 Ie43871350b062263474a7e0dbca850ce <=  Ic772211084626d2ed3ddc4f32b467c6c;
 I12d1f6ac4ef39cb76907b09745b4f8ad <=  Ifcba38a9a6ca0931ba9d86396f257929;
 If9b05209071a1c16ecce1c28f886ee1d <=  I3ae9dbf37dbadabaf8a56188eae40288;
 Iebb87060282934e67cd1e7e8493fcf20 <=  Iae4d59e569911a81bb653cdb58c65137;
 I22b235f6e6f0938fe2a026f91bfd72cf <=  I9b12cb33d0f37813bd735c14d8be517e;
 I185299c78eca06f6174996089a2df4d5 <=  Ifab01268c2a1f0385dc4b18a9d488321;
 I90f70f8385f7d8fc69fe21f42d96eeeb <=  Ie0f0a8cf008e6a10d1698c11c380df97;
 I5d03a9d2e8ca426a10005cf5a1689f4f <=  I99aa62ad841c5bd5b1f2b6758d046784;
 I1f30e3cf906aa5a09d71f23c5be461ba <=  I3fc64e5c431cd64d48f3cc5c9c86f342;
 I13069dca0bc85e00a513e9fe7562b346 <=  I65a139ae2fa69f57c3a8ed35e00e29ae;
 Ib69a5ff88f694a3cf18fa11fcccdd9c2 <=  I628bc7c30b5e896c2b8f4af752b44637;
 If4b3a419df7ce8b8cd5f2b7a26e1a629 <=  I5c7ed27126a8097481ab5f966867783b;
 I03b2bc96c0edf4f4c27ab02d8beda293 <=  I686481757183441e45d85fece1a7b514;
 Iddd38c69253e1ba79f6762c9e69857ad <=  I10929316643f6670bedc63e77b293c97;
 I3437ae400dbe3a2eb99a65a263889bb6 <=  Ia66d818d01365175f416a4de87a281bb;
 I0bb76633859552dc99f63b3c520037cc <=  I7711386635a1760e7976d0947e0a5f8a;
 Ifcb79d8780c0e5859fc885521a3a4070 <=  I4b2cc8ae58d2fb89bd9095b2bb688cbe;
 Ia43aac10d65d1661b3d7f9968c829c21 <=  Ied1035a697824a18281435fe2b7f1f56;
 I6ecfb2be423754892a663315c2c74440 <=  I3e9ecaf8da044766c57685a1065ce10a;
 Ic9b31062ba9aedcda0f4c91e39fe1814 <=  Ibebda2f9816088ea15cd5b4f555c5d33;
 Ie5ff9375515964757ffe821812ed8e73 <=  I6043631f93e2c514d5ed6e86beffa7c6;
 I5152ee18b04c8d038ead4817bc68fa57 <=  Ibc084904fb63bb24102789357ce2cd76;
 I606544d89b457531a204f0a9a061dc74 <=  I9e82413dca68de150b81bd27ab180980;
 If7bcb8673722495218ae395b5716c89a <=  I4992c306a07d2e104a72dfcc37968e8c;
 I755d5c8837cace07fc3c0393a6ba2a43 <=  I637c0445b26879a0fb9d7d94baef55e4;
 I2051dc0ec4b2e1de6e3308c6e0ae74bd <=  I3f1f9cecc45287a2c9487c04d8430b5b;
 I9ff8a14d8788f2e0deb7a0c1f4d0fa0d <=  Ife3d2f48786c2e11f7c4f8b4a7bb829e;
 Id017562a43e853ec27712b3f8d449361 <=  I0a019e2861b41f395bd12b43cd978e59;
 I7c408398d6b1e91c00962636fbf59b83 <=  I34fcd098fa2b426f98542121dae204fc;
 I53387cf352304840ccae53d5b5b153e7 <=  I8c9a0911720c403f2794fa5662a31207;
 I6d483d27683d84d2309d756d36f43ae9 <=  I11af377ea2ae07f2249042a6daeef846;
 I1c44630f8f2d9bf2a5df81f22a67ed43 <=  Ib5d6d77cf92f29c1b498252859ec19ff;
 Ic7a0ea4cb5954db181b37e8072cf54fb <=  I1d6100bd00e7e46af792dd99286391a5;
 I591e5713ec07915309f4a588ea51a990 <=  Ia6e85ec8c498ed70cb4a4e01bf8d1530;
 Ibab6e2a97bd19438998b97780bdae17d <=  Icc6d40c383e5580bbac65b6c77da6528;
 Icb868f4e4f276036478f3977e8d831a3 <=  Id939e83f81205a66485908e0bba8504d;
 I8dde06b1ca763ca0cdd273e440de86ab <=  Ie709765eec241ae95c588fbfed18a87e;
 I44049fcab453cba240bed48d89a664e5 <=  I497fb247a6572f689aea3e595e657fdb;
 I4c6d3af7a2d1adb1f60b61a523dd9bff <=  I659b78a601b47941441dc1debcae4d46;
 I70d83e5081cd2c9051f9c6b8652462d7 <=  Ibed2d1ab1707ca759a8b09a5147a4268;
 Id841c70607e96ab5144c91a573a771c7 <=  I23c058e418bad060fb1404b248782705;
 Ib9318ad9f3aa8b5fd8b8c59fe3bd1616 <=  I95f73f2e7a5268d25f4fcaa53339c2fc;
 I569eefbb2dbaf1e589f1cf1bc35721c7 <=  I90b927c01ca8d69239141958db410c54;
 Id399e2be28090c81e93743f1bfe00347 <=  I79c64b98cdd4f4a1b41ddd2480c5d62a;
 I04b7604f3936be2c49deb140a0d1eae5 <=  I76071439d501dfac67b1355c33f04c79;
 I23d474402240b1761c2f9d785cd2973b <=  I3bed56f31105c1dd5524f2e04a6cdc0f;
 Ia5bbbcb8956d08a529457d6ca2c38ebc <=  I1ca06bac6a4d082efeed13d0448630fb;
 I116f8968c4a02e2a22a8ea4eb5dd3951 <=  Iefd7ba660203932e953d509b10032e4d;
 I1ebdf4675d0986c912c52af538ac358d <=  I76b3bd4ded426c469b208f83f7bb1781;
 I92cd919b7b5b4ca8984668bfbdb43d3b <=  I36261da4cc2946a22e80fb6f2a394753;
 Ibdecc8406ba4102713fde4a51206403f <=  Iaa84b434bf0040f25a2dd6af77d90df4;
 Ie79b340519a003c4388b90a3d8fac445 <=  I1a314b0ac2b2897b23d2e9fd3e5e63f0;
 I719e56962c59071b4783ff87e554a37e <=  I64eff7490d835e24cf4e5f4d0c60e18e;
 Id2a6a7580c31d450f8c78217e8997f7e <=  I95c886a9726c33f2a8f2f9413c9486cb;
 I74f0171925c0986fe140602b09a0caf2 <=  Ie2fbf1593b8aa394377ccc4ef0f705b6;
 I5e9bef3789fd851fb793bea78beef829 <=  I124a5e6d2c3103fbb4699cc2f7528a48;
 I0f3062a73289917dc123b87666bdad07 <=  I3625276282d727c6510f5123ee467e73;
 I238a8e826a1d8f069455ae0163d508f2 <=  I771e25faed091d437e00dae0e66d088b;
 Iedd0e164003fd9532945df51a5408307 <=  Iad7a84f48832522261c3495844b19dde;
 Ib8a70644d197140114eacd4c9612dd77 <=  I8de675a8e37ed2b30a82e49ff6d510a0;
 Ib171958fe2af1d20130ca83b668af768 <=  I4bbc70e0a3a56eeb62af73e6c80006b4;
 I80d67b47c44a3b424d1ed4c8e357c265 <=  I5c97bebf3cd2472e43ae7312d3956bb5;
 Iaa9183f11cd736e6271b9e6259a807a7 <=  I527847fbb55900e97761446b030ed540;
 I1f2ac0b753cee68f5e984de8994f2f0d <=  Ie707c8b057532a88aff15ca43d1a4cef;
 I495ac3abe6643625add1aeef4776b39e <=  I41708d131f34ee41b74f571661e751c6;
 I4c8185fc93a069b6fa81b3936de2b4b0 <=  I410af2866a81357ed84738c1800ee8e2;
 Ib05eddf67c2a5797e8e0e733fca4328b <=  Iae78b53a85d3b3441bb251688c85fe66;
 I8f8316a85f64267a15f99a0b47db5f08 <=  I1c4646eab74db4876187e2e87d861e4d;
 I69116a38d209590270e61cfe9d2e56d5 <=  Idb04b139376a9fd83c6f921b02c31849;
 I713819fe0cf6d54393d9cd5a32a37807 <=  I64c0c3c0d18d18ed62b2b2910930f8a0;
 I811d183d31135919e65f87250c0ba456 <=  I0c622446a77fe077062fd87448e11fec;
 I8a99662ff2d2b8f153d6d9359b88eff5 <=  Ie69cbbb6131f04ccf84db28990b4dbdd;
 Ib246205f26dd43b9d1fa057a2179e4b2 <=  Id0b467dbeaa2b30126ed60489530e29f;
 I972077c6595b44e3113b0d7a925aa913 <=  Idac7b0bec594eccd74ac2d944da4484e;
 Idde043a5721004c3904eb2b55031e7c1 <=  I4ddb027f246fb2b145bba7b01687d39b;
 Iebfd00d9a2a6e39e6fc73f95c4f29539 <=  I754ff7341b379de55d5facc6fcc9f874;
 I3e10f0cc7d257acf63a5ca7a0cb9c7cf <=  Ia7a71696b5ebed6c80cafb33a031626e;
 I62895b1265f950882fc5fb770dafd51d <=  I542db58e949d7d1c542c075005fb065c;
 I9f890d3f6b5edfbf106d59df07cb1b68 <=  I28aaa9370cb22a81b7c8d20fe7e1d347;
 Icd6b85be80234c06eaeaf1347ebabb38 <=  If4abfdcd468d4d98db5f32bb99303035;
 I1e9047545567e723fa101ab94dffa45f <=  Idfc14e592719d57828f8e6dc2130e270;
 Iea7a223f22fb02e29871f500b61fa205 <=  Ia51b4598ba3f6c128ffcd421a3ba7309;
 Ida8637c3dd298410093697077abad3e0 <=  Iee935e25f9fe5c7844bb0c0490cbb90f;
 Ic767ff5ab4bfc377cf1b7bae10b42d3e <=  I05d0b3631f8501ecafcbb321c15be5f1;
 Ieafe43b66027e5b192cdd5fe25977f4c <=  I7ea9adf8dba141eef7a08d76105580ec;
 I41d92f30c38301789ac4155986c2a634 <=  Ifa4cd939b137dc050f675a493546ddf6;
 I5c4bedc45aa3faab29c3547e29c6db68 <=  I7a6215a05dd8dbdcb421d7df535c5b67;
 I1bf648fa37015e2997a689769881149c <=  Ibd0c06d4190a37b90c51d562c6019551;
 I4f38b0092062a40f0bd68bbe8911f248 <=  I75b4b57cf9d7400feec38e037c948352;
 I74c408ce157c47049698b52949d1fd38 <=  I14a4e51be5aa98fa28cc4740e6446747;
 I3ed597f1774bf9274566cb5fc7dbbdc5 <=  I43196769a96d15dd03318e43b48a6b4d;
 I8d111345e29debfc7addbb913d4e9054 <=  I8494b9c75594140fabc1158bacf4438a;
 I8d19b379f6693601f18ea748bbbadf9b <=  I931bf44a358d9fd91d31aa78d3e16312;
 I68521e797f1f404e6a190855b1a322f1 <=  I5355f3939098f1ae0aa0f254b8e7e163;
 I5ecffa51c73d64359ba32c2cf56c6b7a <=  I6228ab1c737aec5845684c0eff41dac4;
 I2adb86feb263103c1419d34eb9b8ae4e <=  I9034255c2128aa8c4d707bf003a57e86;
 I733561ae7e5600d8275667457f2ea151 <=  Ia9bc32f3ef4f4681782fec452e572cf2;
 I4db74afe0a9f15f643d8295051f762c0 <=  I9791a65b490a63c3c201409a30b86199;
 Id194460b74adf4856635d5c432ea772f <=  Id5297cb2f91d5b3e67c4bd97a8c05401;
 Ifc1dfcb0afd77d1a01bbb54da77a5f70 <=  Ibc826b606b10904061b2666eb204469e;
 I0cec4bb6f8f736beea5fd2dc57310432 <=  I06dabbc9dc6fb6b8fa517e188ee74208;
 If878a4e87d963261e36cde448d6c3bbc <=  I4d3607d7cd13b86ae4a22bebaf65ef0e;
 I2d28d468beee8a809ece79a2b7b07d27 <=  Ia974eebd7b7563b2f0822f538c13a911;
 I8b553bf742d14f23835e62aeade33413 <=  I191470ccfa2c2838a34aceb571582bb4;
 Iacc099c63faabe7dda342eafe07e26d4 <=  I01714219c84cfbfd7ff940108ddbb6b3;
 Ifc3d28213bc38fbcff2eb42ebc350c8a <=  I118d11a015af5944d64290a46bf49c09;
 I7fd466826e266237c64dd4010bf19ed8 <=  Ib878ef5592b0bf1af247ede54fe13a45;
 I5c42c7a5b8b8d73e5374eb00cf80f91b <=  I7686f623f51c5a9f8f3f8d143ed8bcb5;
 I2e4f341a2f112ba1df12c82183bd3566 <=  I4d48fc8081756af036b8f1b1b9e56051;
 I757c6c719d8455faea81fa0901a2c15e <=  Ia1d93d4bbc6b1e73dbb0c6c26d102f10;
 Ie146524ab065ed90500947d0e77f7e5e <=  Ifb7d0d12a916fc3f2f9c0341f27ef53f;
 I40fd0db59f8b8877f3f62b9b87e2892d <=  I4ee596c96f91a18ef1ebb0ee6de285ae;
 I2c05c52719e300f911b6245928a40fb3 <=  I5aeda0b5dc8459d86e9ab5082bf9fed8;
 I07acde143b8be8c4ec4e562a66562b58 <=  I7b6ff145fa076d152af672e0c3a062bc;
 I5d0ae3e1a3333e7dcc389a609644376a <=  I3929cfb9fb8795d4dd9f54f9c4a2fa02;
 I13b47a7b710051dde6ab5cae17f216d4 <=  If33f043047ad17b323733a201aa649da;
 I1c0174a95fd6b5322576907671acdd82 <=  Icfb9314b47604c3b065ffdd5d9042682;
 Ica09fab419a2bd1a966956988b6507b3 <=  I5cd61f07b490ca79f1ec069ed2d47528;
 I27097218191d9ad8cd380a75b5b4d467 <=  I1bace448ce54ae41e9e8d27acf548338;
 I354ec2d3605e41d982076dcb7e32d2c1 <=  I692bf3f934f0ee8fbf02c7dce98f924c;
 I14c93bdff35500174e3db5c18b48cb94 <=  Ifb3af535b42775dae1e0ade2d8bf79df;
 I30084765c13a4c6a7514a16e3f45a9c2 <=  I569a621522dd636df609f60c1b22d7f7;
 I1f07b4c82c226595be454e07eed346ab <=  Ic651187a36eb89eaf129a368af3474ee;
 I7401e0464789f88be2b661eb055bbdef <=  Ib120bd9cfec97e7956bb64f8e4527caf;
 Ia1e603a00bf98ee21caea749765ed341 <=  I41e452eee26c8ede812d3ca957488aec;
 I7aa491e6301b27435c2dadebe447b43a <=  I99ba3451537a2876c9f585f72911bc4f;
end
