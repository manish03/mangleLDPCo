reg [fgallag_WDTH -1:0] fgallag0x00004_0, fgallag0x00004_0_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_1, fgallag0x00004_1_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_2, fgallag0x00004_2_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_3, fgallag0x00004_3_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_4, fgallag0x00004_4_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_5, fgallag0x00004_5_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_6, fgallag0x00004_6_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_7, fgallag0x00004_7_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_8, fgallag0x00004_8_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_9, fgallag0x00004_9_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_10, fgallag0x00004_10_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_11, fgallag0x00004_11_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_12, fgallag0x00004_12_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_13, fgallag0x00004_13_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_14, fgallag0x00004_14_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_15, fgallag0x00004_15_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_16, fgallag0x00004_16_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_17, fgallag0x00004_17_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_18, fgallag0x00004_18_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_19, fgallag0x00004_19_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_20, fgallag0x00004_20_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_21, fgallag0x00004_21_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_22, fgallag0x00004_22_q;
reg [fgallag_WDTH -1:0] fgallag0x00004_23, fgallag0x00004_23_q;
reg start_d_fgallag0x00004_q ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 fgallag0x00004_0_q <= 'h0;
 fgallag0x00004_1_q <= 'h0;
 fgallag0x00004_2_q <= 'h0;
 fgallag0x00004_3_q <= 'h0;
 fgallag0x00004_4_q <= 'h0;
 fgallag0x00004_5_q <= 'h0;
 fgallag0x00004_6_q <= 'h0;
 fgallag0x00004_7_q <= 'h0;
 fgallag0x00004_8_q <= 'h0;
 fgallag0x00004_9_q <= 'h0;
 fgallag0x00004_10_q <= 'h0;
 fgallag0x00004_11_q <= 'h0;
 fgallag0x00004_12_q <= 'h0;
 fgallag0x00004_13_q <= 'h0;
 fgallag0x00004_14_q <= 'h0;
 fgallag0x00004_15_q <= 'h0;
 fgallag0x00004_16_q <= 'h0;
 fgallag0x00004_17_q <= 'h0;
 fgallag0x00004_18_q <= 'h0;
 fgallag0x00004_19_q <= 'h0;
 fgallag0x00004_20_q <= 'h0;
 fgallag0x00004_21_q <= 'h0;
 fgallag0x00004_22_q <= 'h0;
 fgallag0x00004_23_q <= 'h0;
 start_d_fgallag0x00004_q <= 'h0;
end
else
begin
 fgallag0x00004_0_q <=  fgallag0x00004_0;
 fgallag0x00004_1_q <=  fgallag0x00004_1;
 fgallag0x00004_2_q <=  fgallag0x00004_2;
 fgallag0x00004_3_q <=  fgallag0x00004_3;
 fgallag0x00004_4_q <=  fgallag0x00004_4;
 fgallag0x00004_5_q <=  fgallag0x00004_5;
 fgallag0x00004_6_q <=  fgallag0x00004_6;
 fgallag0x00004_7_q <=  fgallag0x00004_7;
 fgallag0x00004_8_q <=  fgallag0x00004_8;
 fgallag0x00004_9_q <=  fgallag0x00004_9;
 fgallag0x00004_10_q <=  fgallag0x00004_10;
 fgallag0x00004_11_q <=  fgallag0x00004_11;
 fgallag0x00004_12_q <=  fgallag0x00004_12;
 fgallag0x00004_13_q <=  fgallag0x00004_13;
 fgallag0x00004_14_q <=  fgallag0x00004_14;
 fgallag0x00004_15_q <=  fgallag0x00004_15;
 fgallag0x00004_16_q <=  fgallag0x00004_16;
 fgallag0x00004_17_q <=  fgallag0x00004_17;
 fgallag0x00004_18_q <=  fgallag0x00004_18;
 fgallag0x00004_19_q <=  fgallag0x00004_19;
 fgallag0x00004_20_q <=  fgallag0x00004_20;
 fgallag0x00004_21_q <=  fgallag0x00004_21;
 fgallag0x00004_22_q <=  fgallag0x00004_22;
 fgallag0x00004_23_q <=  fgallag0x00004_23;
 start_d_fgallag0x00004_q <=  start_d_fgallag0x00003_q;
end
