reg [fgallag_WDTH -1:0] I67f92596363d7abd702880c8dd319453, I03b14329c0d52c7997914a8d9ab65fed;
reg [fgallag_WDTH -1:0] I58dc37dd8f90b2815ebae43223ff2268, I63a4e0a46ca3426e2cb066ad3bfc245d;
reg [fgallag_WDTH -1:0] Ic5c9b0ef750a107380673521819d09e5, Ie21703557f53d7bf9cf79a7f6c1d5958;
reg [fgallag_WDTH -1:0] I6d82716e87b1ac554c6ff5e4169afe0b, I3a7b809a0160dee33125934243952cdc;
reg [fgallag_WDTH -1:0] I64fc488e4651b1cde21e870d2528613c, I1cb33fdd3dac4dda0b25adbab30d2913;
reg [fgallag_WDTH -1:0] Ice7c81f4524a3e2a6ec0b6e7d76fe9b6, Ia6905a32e1257061364dd1249fa76bf2;
reg [fgallag_WDTH -1:0] If1b3191923af5d433e5d97adf41bd97f, Id2b87d69ba4c78cf41a7be349397ad5e;
reg [fgallag_WDTH -1:0] If2cca0ade959a72defe62fb3eef484e4, I7d9d74dbceb047ad0c76322038fbf229;
reg [fgallag_WDTH -1:0] Ida8b253166cc056c54916e14755c6aa6, I856e4e862c70da83553a3dba9edea1ab;
reg [fgallag_WDTH -1:0] If1ac872a756deb15fa93f38bc63700c3, Iaf42178313f7b4aa6ce6090ecbf2b3b6;
reg [fgallag_WDTH -1:0] Ia8342322e4b86c946f8a133fc284bd4f, Id7a56c8135dad1fd457d336f7a632436;
reg [fgallag_WDTH -1:0] I316bb23418efb56e676cc0a58e8f0e19, I2ffc40e4b0cc841bd3c8d7519fc4512a;
reg [fgallag_WDTH -1:0] Ib659aa347010e749163015d2457712b7, I20c0389215371104437ef298cb12b3c4;
reg [fgallag_WDTH -1:0] Id87f3e882b2fb1c5af8b4134c83dff16, Ie4e1b20f36ecda5d4d917a241ef2a1fd;
reg [fgallag_WDTH -1:0] I0eda2f2f507535ab778d59c7ce193447, Icf120a29648cb8af4bae9e4343f13a40;
reg [fgallag_WDTH -1:0] If36a4176048d1fec4e9646d016b5a33b, I1e317164e9010fb6755c65adda38ea2a;
reg [fgallag_WDTH -1:0] Id3ffa72548f440a0e3a90db8b5ff1c39, I0f5a57095bb2bbf99b71f04a19e2c38f;
reg [fgallag_WDTH -1:0] Ic36450e12061ae80189b6f16d1cab329, Ib52869a26824ee42fff6262100e1ebe5;
reg [fgallag_WDTH -1:0] Iec0fe238288bd4b3f41ddec347477271, I61ff69ca863e90ffc9118f12c5aa3b14;
reg [fgallag_WDTH -1:0] Iff515d269a292258ff61605083324963, Iad3702f89b5505a20193d89537b49edc;
reg [fgallag_WDTH -1:0] I13b529dfc9f09f5208d2df5a91e4eabe, I08f41ede762b72d92816c6dff8e074f9;
reg [fgallag_WDTH -1:0] If5686d7de8ada834d078111dd1557853, I0d0befb35bf5e3529b47e296923360d6;
reg [fgallag_WDTH -1:0] I4393932a40ca1c79aa95d652d504c5f6, I912919c7cfae1b4827ca945a92a5310c;
reg [fgallag_WDTH -1:0] Ia4abb71881c5f95a1a30badf83a0a567, Icd7b7d17911094c9fa48fc5906968dcd;
reg I64ddd9e95d971d161174a6dd0c3d2fbe ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I03b14329c0d52c7997914a8d9ab65fed <= 'h0;
 I63a4e0a46ca3426e2cb066ad3bfc245d <= 'h0;
 Ie21703557f53d7bf9cf79a7f6c1d5958 <= 'h0;
 I3a7b809a0160dee33125934243952cdc <= 'h0;
 I1cb33fdd3dac4dda0b25adbab30d2913 <= 'h0;
 Ia6905a32e1257061364dd1249fa76bf2 <= 'h0;
 Id2b87d69ba4c78cf41a7be349397ad5e <= 'h0;
 I7d9d74dbceb047ad0c76322038fbf229 <= 'h0;
 I856e4e862c70da83553a3dba9edea1ab <= 'h0;
 Iaf42178313f7b4aa6ce6090ecbf2b3b6 <= 'h0;
 Id7a56c8135dad1fd457d336f7a632436 <= 'h0;
 I2ffc40e4b0cc841bd3c8d7519fc4512a <= 'h0;
 I20c0389215371104437ef298cb12b3c4 <= 'h0;
 Ie4e1b20f36ecda5d4d917a241ef2a1fd <= 'h0;
 Icf120a29648cb8af4bae9e4343f13a40 <= 'h0;
 I1e317164e9010fb6755c65adda38ea2a <= 'h0;
 I0f5a57095bb2bbf99b71f04a19e2c38f <= 'h0;
 Ib52869a26824ee42fff6262100e1ebe5 <= 'h0;
 I61ff69ca863e90ffc9118f12c5aa3b14 <= 'h0;
 Iad3702f89b5505a20193d89537b49edc <= 'h0;
 I08f41ede762b72d92816c6dff8e074f9 <= 'h0;
 I0d0befb35bf5e3529b47e296923360d6 <= 'h0;
 I912919c7cfae1b4827ca945a92a5310c <= 'h0;
 Icd7b7d17911094c9fa48fc5906968dcd <= 'h0;
 I64ddd9e95d971d161174a6dd0c3d2fbe <= 'h0;
end
else
begin
 I03b14329c0d52c7997914a8d9ab65fed <=  I67f92596363d7abd702880c8dd319453;
 I63a4e0a46ca3426e2cb066ad3bfc245d <=  I58dc37dd8f90b2815ebae43223ff2268;
 Ie21703557f53d7bf9cf79a7f6c1d5958 <=  Ic5c9b0ef750a107380673521819d09e5;
 I3a7b809a0160dee33125934243952cdc <=  I6d82716e87b1ac554c6ff5e4169afe0b;
 I1cb33fdd3dac4dda0b25adbab30d2913 <=  I64fc488e4651b1cde21e870d2528613c;
 Ia6905a32e1257061364dd1249fa76bf2 <=  Ice7c81f4524a3e2a6ec0b6e7d76fe9b6;
 Id2b87d69ba4c78cf41a7be349397ad5e <=  If1b3191923af5d433e5d97adf41bd97f;
 I7d9d74dbceb047ad0c76322038fbf229 <=  If2cca0ade959a72defe62fb3eef484e4;
 I856e4e862c70da83553a3dba9edea1ab <=  Ida8b253166cc056c54916e14755c6aa6;
 Iaf42178313f7b4aa6ce6090ecbf2b3b6 <=  If1ac872a756deb15fa93f38bc63700c3;
 Id7a56c8135dad1fd457d336f7a632436 <=  Ia8342322e4b86c946f8a133fc284bd4f;
 I2ffc40e4b0cc841bd3c8d7519fc4512a <=  I316bb23418efb56e676cc0a58e8f0e19;
 I20c0389215371104437ef298cb12b3c4 <=  Ib659aa347010e749163015d2457712b7;
 Ie4e1b20f36ecda5d4d917a241ef2a1fd <=  Id87f3e882b2fb1c5af8b4134c83dff16;
 Icf120a29648cb8af4bae9e4343f13a40 <=  I0eda2f2f507535ab778d59c7ce193447;
 I1e317164e9010fb6755c65adda38ea2a <=  If36a4176048d1fec4e9646d016b5a33b;
 I0f5a57095bb2bbf99b71f04a19e2c38f <=  Id3ffa72548f440a0e3a90db8b5ff1c39;
 Ib52869a26824ee42fff6262100e1ebe5 <=  Ic36450e12061ae80189b6f16d1cab329;
 I61ff69ca863e90ffc9118f12c5aa3b14 <=  Iec0fe238288bd4b3f41ddec347477271;
 Iad3702f89b5505a20193d89537b49edc <=  Iff515d269a292258ff61605083324963;
 I08f41ede762b72d92816c6dff8e074f9 <=  I13b529dfc9f09f5208d2df5a91e4eabe;
 I0d0befb35bf5e3529b47e296923360d6 <=  If5686d7de8ada834d078111dd1557853;
 I912919c7cfae1b4827ca945a92a5310c <=  I4393932a40ca1c79aa95d652d504c5f6;
 Icd7b7d17911094c9fa48fc5906968dcd <=  Ia4abb71881c5f95a1a30badf83a0a567;
 I64ddd9e95d971d161174a6dd0c3d2fbe <=  I4da12bc20380296febc560ba65f58a8e;
end
