//`include "GF2_LDPC_fgallag_0x00004_assign_inc.sv"
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00000] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00000] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00001] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00001] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00002] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00003] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00002] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00004] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00005] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00003] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00006] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00007] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00004] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00008] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00009] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00005] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0000a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0000b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00006] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0000c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0000d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00007] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0000e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0000f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00008] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00010] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00011] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00009] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00012] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00013] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00014] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00015] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00016] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00017] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00018] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00019] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0001a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0001b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0001c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0001d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0001e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0001f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00010] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00020] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00021] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00011] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00022] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00023] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00012] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00024] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00025] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00013] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00026] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00027] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00014] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00028] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00029] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00015] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0002a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0002b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00016] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0002c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0002d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00017] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0002e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0002f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00018] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00030] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00031] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00019] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00032] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00033] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00034] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00035] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00036] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00037] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00038] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00039] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0003a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0003b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0003c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0003d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0003e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0003f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00020] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00040] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00041] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00021] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00042] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00043] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00022] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00044] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00045] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00023] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00046] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00047] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00024] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00048] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00049] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00025] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0004a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0004b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00026] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0004c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0004d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00027] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0004e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0004f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00028] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00050] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00051] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00029] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00052] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00053] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00054] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00055] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00056] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00057] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00058] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00059] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0005a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0005b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0005c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0005d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0005e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0005f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00030] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00060] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00061] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00031] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00062] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00063] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00032] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00064] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00065] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00033] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00066] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00067] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00034] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00068] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00069] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00035] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0006a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0006b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00036] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0006c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0006d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00037] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0006e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0006f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00038] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00070] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00071] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00039] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00072] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00073] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00074] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00075] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00076] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00077] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00078] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00079] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0007a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0007b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0007c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0007d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0007e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0007f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00040] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00080] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00081] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00041] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00082] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00083] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00042] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00084] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00085] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00043] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00086] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00087] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00044] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00088] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00089] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00045] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0008a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0008b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00046] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0008c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0008d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00047] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0008e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0008f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00048] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00090] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00091] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00049] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00092] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00093] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00094] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00095] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00096] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00097] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00098] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00099] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0009a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0009b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0009c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0009d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0009e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0009f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00050] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000a0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000a1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00051] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000a2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000a3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00052] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000a4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000a5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00053] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000a6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000a7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00054] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000a8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000a9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00055] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000aa] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ab] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00056] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ac] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ad] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00057] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ae] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000af] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00058] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000b0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000b1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00059] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000b2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000b3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000b4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000b5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000b6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000b7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000b8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000b9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ba] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000bb] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000bc] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000bd] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000be] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000bf] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00060] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000c0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000c1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00061] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000c2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000c3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00062] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000c4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000c5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00063] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000c6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000c7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00064] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000c8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000c9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00065] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ca] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000cb] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00066] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000cc] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000cd] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00067] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ce] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000cf] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00068] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000d0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000d1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00069] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000d2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000d3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000d4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000d5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000d6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000d7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000d8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000d9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000da] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000db] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000dc] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000dd] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000de] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000df] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00070] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000e0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000e1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00071] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000e2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000e3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00072] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000e4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000e5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00073] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000e6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000e7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00074] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000e8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000e9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00075] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ea] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000eb] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00076] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ec] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ed] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00077] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ee] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ef] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00078] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000f0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000f1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00079] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000f2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000f3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000f4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000f5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000f6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000f7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000f8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000f9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000fa] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000fb] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000fc] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000fd] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000fe] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h000ff] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00080] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00100] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00101] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00081] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00102] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00103] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00082] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00104] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00105] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00083] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00106] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00107] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00084] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00108] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00109] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00085] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0010a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0010b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00086] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0010c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0010d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00087] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0010e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0010f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00088] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00110] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00111] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00089] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00112] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00113] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00114] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00115] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00116] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00117] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00118] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00119] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0011a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0011b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0011c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0011d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0011e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0011f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00090] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00120] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00121] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00091] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00122] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00123] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00092] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00124] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00125] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00093] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00126] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00127] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00094] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00128] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00129] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00095] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0012a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0012b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00096] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0012c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0012d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00097] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0012e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0012f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00098] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00130] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00131] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00099] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00132] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00133] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00134] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00135] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00136] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00137] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00138] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00139] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0013a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0013b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0013c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0013d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0013e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0013f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a0] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00140] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00141] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a1] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00142] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00143] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a2] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00144] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00145] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a3] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00146] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00147] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a4] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00148] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00149] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a5] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0014a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0014b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a6] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0014c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0014d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a7] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0014e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0014f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a8] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00150] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00151] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a9] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00152] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00153] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000aa] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00154] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00155] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ab] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00156] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00157] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ac] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00158] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00159] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ad] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0015a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0015b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ae] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0015c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0015d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000af] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0015e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0015f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b0] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00160] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00161] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b1] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00162] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00163] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b2] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00164] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00165] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b3] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00166] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00167] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b4] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00168] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00169] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b5] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0016a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0016b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b6] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0016c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0016d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b7] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0016e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0016f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b8] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00170] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00171] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b9] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00172] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00173] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ba] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00174] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00175] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000bb] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00176] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00177] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000bc] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00178] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00179] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000bd] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0017a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0017b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000be] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0017c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0017d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000bf] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0017e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0017f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c0] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00180] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00181] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c1] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00182] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00183] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c2] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00184] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00185] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c3] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00186] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00187] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c4] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00188] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00189] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c5] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0018a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0018b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c6] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0018c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0018d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c7] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0018e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0018f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c8] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00190] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00191] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c9] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00192] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00193] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ca] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00194] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00195] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000cb] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00196] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00197] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000cc] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00198] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00199] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000cd] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0019a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0019b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ce] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0019c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0019d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000cf] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0019e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0019f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d0] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001a0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001a1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d1] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001a2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001a3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d2] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001a4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001a5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d3] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001a6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001a7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d4] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001a8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001a9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d5] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001aa] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ab] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d6] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ac] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ad] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d7] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ae] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001af] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d8] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001b0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001b1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d9] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001b2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001b3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000da] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001b4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001b5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000db] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001b6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001b7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000dc] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001b8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001b9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000dd] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ba] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001bb] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000de] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001bc] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001bd] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000df] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001be] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001bf] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e0] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001c0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001c1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e1] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001c2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001c3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e2] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001c4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001c5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e3] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001c6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001c7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e4] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001c8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001c9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e5] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ca] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001cb] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e6] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001cc] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001cd] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e7] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ce] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001cf] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e8] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001d0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001d1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e9] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001d2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001d3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ea] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001d4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001d5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000eb] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001d6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001d7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ec] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001d8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001d9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ed] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001da] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001db] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ee] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001dc] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001dd] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ef] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001de] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001df] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f0] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001e0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001e1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f1] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001e2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001e3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f2] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001e4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001e5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f3] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001e6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001e7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f4] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001e8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001e9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f5] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ea] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001eb] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f6] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ec] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ed] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f7] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ee] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ef] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f8] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001f0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001f1] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f9] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001f2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001f3] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000fa] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001f4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001f5] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000fb] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001f6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001f7] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000fc] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001f8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001f9] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000fd] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001fa] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001fb] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000fe] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001fc] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001fd] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ff] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001fe] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h001ff] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00100] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00200] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00201] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00101] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00202] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00203] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00102] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00204] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00205] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00103] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00206] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00207] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00104] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00208] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00209] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00105] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0020a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0020b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00106] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0020c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0020d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00107] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0020e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0020f] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00108] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00210] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00211] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00109] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00212] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00213] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00214] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00215] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00216] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00217] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00218] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00219] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0021a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0021b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0021c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0021d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0021e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0021f] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00110] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00220] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00111] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00222] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00223] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00112] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00224] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00225] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00113] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00226] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00227] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00114] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00228] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00229] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00115] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0022a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0022b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00116] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0022c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0022d] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00117] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0022e] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00118] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00230] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00231] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00119] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00232] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00233] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00234] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00235] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00236] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00237] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00238] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0023a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0023b] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0023c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0023d] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0023e] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00120] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00240] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00241] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00121] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00242] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00243] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00122] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00244] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00245] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00123] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00246] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00124] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00248] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00249] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00125] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0024a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0024b] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00126] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0024c] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00127] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0024e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0024f] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00128] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00250] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00129] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00252] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00253] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00254] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00255] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00256] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00258] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00259] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0025a] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012e] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0025c] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0025d] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012f] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0025e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0025f] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00130] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00260] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00131] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00262] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00263] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00132] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00264] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00133] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00266] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00267] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00134] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00268] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00135] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0026a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0026b] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00136] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0026c] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00137] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0026e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0026f] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00138] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00270] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00139] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00272] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00273] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00274] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00276] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00277] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00278] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0027a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0027b] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0027c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0027e] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00140] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00280] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00281] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00141] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00282] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00142] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00284] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00285] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00143] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00286] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00144] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00288] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00145] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0028a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0028b] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00146] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0028c] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00147] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0028e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0028f] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00148] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00290] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00149] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00292] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014a] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00294] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00295] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00296] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00298] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0029a] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0029b] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0029c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0029e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00150] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00151] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00152] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002a4] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00153] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002a6] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002a7] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00154] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00155] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002aa] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00156] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002ac] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002ad] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00157] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00158] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002b0] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00159] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002b2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002b3] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0015a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0015b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0015c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002b8] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0015d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002ba] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002bb] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0015e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0015f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002be] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00160] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002c0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002c1] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00161] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00162] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00163] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002c6] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00164] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002c8] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002c9] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00165] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00166] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00167] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00168] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002d0] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00169] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002d2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002d3] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0016a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0016b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0016c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002d8] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0016d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002da] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002db] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0016e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0016f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00170] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00171] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002e2] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00172] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002e4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002e5] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00173] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00174] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00175] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00176] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00177] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002ee] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00178] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002f0] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002f1] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00179] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0017a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0017b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0017c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002f8] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0017d] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002fa] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002fb] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0017e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0017f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h002fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00180] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00300] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00181] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00302] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00182] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00304] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00183] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00306] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00184] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00308] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00309] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00185] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0030a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00186] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0030c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00187] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0030e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00188] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00310] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00189] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00312] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0018a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00314] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0018b] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00316] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00317] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0018c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00318] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0018d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0031a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0018e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0031c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0018f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0031e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00190] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00320] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00191] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00322] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00192] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00324] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00193] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00326] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00327] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00194] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00328] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00195] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0032a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00196] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0032c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00197] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0032e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00198] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00330] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00199] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00332] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0019a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00334] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0019b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00336] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0019c] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00338] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00339] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0019d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0033a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0019e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0033c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0019f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0033e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00340] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00342] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00344] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00346] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00348] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0034a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0034c] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a7] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0034e] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0034f] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00350] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00352] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00354] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00356] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00358] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0035a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0035c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0035e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00360] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00362] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00364] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00366] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b4] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00368] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00369] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0036a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0036c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0036e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00370] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00372] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00374] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00376] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00378] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0037a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0037c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0037e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00380] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00382] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00384] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00386] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c4] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00388] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00389] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0038a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0038c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0038e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00390] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00392] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00394] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00396] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00398] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0039a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0039c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0039e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003b0] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d9] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003b2] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003b3] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003f2] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001fa] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003f4] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003f5] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h003fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00200] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00400] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00201] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00402] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00202] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00404] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00203] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00406] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00204] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00408] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00205] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0040a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00206] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0040c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00207] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0040e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00208] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00410] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00209] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00412] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0020a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00414] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0020b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00416] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0020c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00418] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0020d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0041a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0020e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0041c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0020f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0041e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00210] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00420] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00211] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00422] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00212] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00424] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00213] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00426] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00214] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00428] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00215] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0042a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00216] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0042c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00217] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0042e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00218] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00430] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00219] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00432] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0021a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00434] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0021b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00436] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0021c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00438] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0021d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0043a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0021e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0043c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0021f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0043e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00220] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00440] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00221] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00442] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00222] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00444] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00223] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00446] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00224] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00448] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00225] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0044a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00226] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0044c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00227] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0044e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00228] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00450] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00229] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00452] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0022a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00454] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0022b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00456] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0022c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00458] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0022d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0045a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0022e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0045c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0022f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0045e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00230] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00460] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00231] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00462] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00232] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00464] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00233] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00466] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00234] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00468] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00235] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0046a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00236] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0046c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00237] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0046e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00238] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00470] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00239] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00472] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0023a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00474] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0023b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00476] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0023c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00478] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0023d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0047a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0023e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0047c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0023f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0047e] ;
//end
//always_comb begin
              Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00240] = 
          (!fgallag_sel['h00004]) ? 
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00480] : //%
                       I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00481] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00241] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00482] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00242] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00484] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00243] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00486] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00244] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00488] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00245] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0048a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00246] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0048c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00247] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0048e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00248] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00490] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00249] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00492] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0024a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00494] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0024b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00496] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0024c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00498] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0024d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0049a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0024e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0049c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0024f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0049e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00250] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00251] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00252] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00253] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00254] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00255] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00256] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00257] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00258] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00259] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0025a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0025b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0025c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0025d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0025e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0025f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00260] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00261] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00262] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00263] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00264] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00265] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00266] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00267] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00268] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00269] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0026a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0026b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0026c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0026d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0026e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0026f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00270] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00271] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00272] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00273] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00274] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00275] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00276] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00277] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00278] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00279] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0027a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0027b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0027c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0027d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0027e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0027f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h004fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00280] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00500] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00281] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00502] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00282] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00504] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00283] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00506] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00284] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00508] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00285] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0050a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00286] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0050c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00287] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0050e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00288] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00510] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00289] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00512] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0028a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00514] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0028b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00516] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0028c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00518] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0028d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0051a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0028e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0051c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0028f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0051e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00290] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00520] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00291] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00522] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00292] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00524] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00293] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00526] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00294] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00528] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00295] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0052a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00296] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0052c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00297] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0052e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00298] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00530] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00299] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00532] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0029a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00534] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0029b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00536] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0029c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00538] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0029d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0053a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0029e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0053c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0029f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0053e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00540] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00542] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00544] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00546] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00548] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0054a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0054c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0054e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00550] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00552] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00554] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00556] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00558] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0055a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0055c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0055e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00560] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00562] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00564] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00566] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00568] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0056a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0056c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0056e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00570] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00572] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00574] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00576] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00578] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0057a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0057c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0057e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00580] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00582] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00584] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00586] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00588] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0058a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0058c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0058e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00590] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00592] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00594] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00596] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00598] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0059a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0059c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0059e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h005fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00300] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00600] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00301] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00602] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00302] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00604] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00303] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00606] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00304] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00608] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00305] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0060a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00306] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0060c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00307] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0060e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00308] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00610] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00309] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00612] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0030a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00614] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0030b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00616] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0030c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00618] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0030d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0061a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0030e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0061c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0030f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0061e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00310] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00620] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00311] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00622] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00312] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00624] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00313] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00626] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00314] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00628] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00315] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0062a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00316] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0062c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00317] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0062e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00318] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00630] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00319] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00632] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0031a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00634] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0031b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00636] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0031c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00638] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0031d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0063a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0031e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0063c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0031f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0063e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00320] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00640] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00321] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00642] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00322] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00644] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00323] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00646] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00324] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00648] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00325] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0064a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00326] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0064c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00327] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0064e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00328] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00650] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00329] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00652] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0032a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00654] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0032b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00656] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0032c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00658] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0032d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0065a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0032e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0065c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0032f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0065e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00330] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00660] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00331] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00662] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00332] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00664] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00333] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00666] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00334] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00668] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00335] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0066a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00336] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0066c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00337] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0066e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00338] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00670] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00339] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00672] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0033a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00674] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0033b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00676] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0033c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00678] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0033d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0067a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0033e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0067c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0033f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0067e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00340] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00680] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00341] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00682] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00342] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00684] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00343] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00686] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00344] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00688] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00345] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0068a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00346] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0068c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00347] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0068e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00348] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00690] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00349] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00692] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0034a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00694] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0034b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00696] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0034c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00698] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0034d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0069a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0034e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0069c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0034f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0069e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00350] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00351] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00352] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00353] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00354] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00355] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00356] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00357] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00358] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00359] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0035a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0035b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0035c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0035d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0035e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0035f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00360] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00361] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00362] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00363] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00364] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00365] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00366] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00367] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00368] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00369] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0036a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0036b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0036c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0036d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0036e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0036f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00370] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00371] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00372] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00373] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00374] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00375] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00376] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00377] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00378] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00379] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0037a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0037b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0037c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0037d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0037e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0037f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h006fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00380] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00700] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00381] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00702] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00382] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00704] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00383] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00706] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00384] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00708] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00385] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0070a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00386] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0070c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00387] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0070e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00388] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00710] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00389] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00712] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0038a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00714] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0038b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00716] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0038c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00718] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0038d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0071a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0038e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0071c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0038f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0071e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00390] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00720] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00391] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00722] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00392] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00724] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00393] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00726] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00394] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00728] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00395] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0072a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00396] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0072c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00397] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0072e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00398] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00730] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00399] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00732] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0039a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00734] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0039b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00736] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0039c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00738] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0039d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0073a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0039e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0073c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0039f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0073e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00740] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00742] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00744] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00746] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00748] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0074a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0074c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0074e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00750] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00752] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00754] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00756] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00758] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0075a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0075c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0075e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00760] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00762] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00764] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00766] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00768] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0076a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0076c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0076e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00770] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00772] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00774] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00776] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00778] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0077a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0077c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0077e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00780] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00782] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00784] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00786] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00788] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0078a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0078c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0078e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00790] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00792] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00794] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00796] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00798] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0079a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0079c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0079e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h007fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00400] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00800] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00401] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00802] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00402] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00804] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00403] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00806] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00404] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00808] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00405] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0080a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00406] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0080c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00407] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0080e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00408] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00810] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00409] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00812] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0040a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00814] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0040b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00816] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0040c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00818] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0040d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0081a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0040e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0081c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0040f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0081e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00410] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00820] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00411] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00822] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00412] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00824] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00413] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00826] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00414] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00828] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00415] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0082a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00416] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0082c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00417] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0082e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00418] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00830] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00419] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00832] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0041a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00834] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0041b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00836] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0041c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00838] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0041d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0083a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0041e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0083c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0041f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0083e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00420] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00840] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00421] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00842] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00422] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00844] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00423] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00846] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00424] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00848] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00425] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0084a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00426] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0084c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00427] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0084e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00428] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00850] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00429] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00852] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0042a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00854] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0042b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00856] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0042c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00858] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0042d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0085a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0042e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0085c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0042f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0085e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00430] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00860] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00431] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00862] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00432] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00864] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00433] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00866] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00434] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00868] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00435] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0086a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00436] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0086c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00437] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0086e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00438] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00870] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00439] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00872] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0043a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00874] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0043b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00876] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0043c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00878] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0043d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0087a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0043e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0087c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0043f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0087e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00440] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00880] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00441] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00882] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00442] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00884] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00443] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00886] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00444] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00888] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00445] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0088a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00446] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0088c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00447] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0088e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00448] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00890] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00449] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00892] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0044a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00894] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0044b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00896] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0044c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00898] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0044d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0089a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0044e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0089c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0044f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0089e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00450] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00451] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00452] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00453] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00454] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00455] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00456] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00457] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00458] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00459] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0045a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0045b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0045c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0045d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0045e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0045f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00460] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00461] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00462] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00463] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00464] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00465] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00466] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00467] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00468] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00469] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0046a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0046b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0046c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0046d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0046e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0046f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00470] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00471] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00472] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00473] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00474] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00475] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00476] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00477] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00478] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00479] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0047a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0047b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0047c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0047d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0047e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0047f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h008fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00480] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00900] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00481] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00902] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00482] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00904] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00483] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00906] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00484] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00908] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00485] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0090a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00486] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0090c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00487] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0090e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00488] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00910] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00489] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00912] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0048a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00914] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0048b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00916] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0048c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00918] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0048d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0091a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0048e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0091c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0048f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0091e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00490] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00920] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00491] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00922] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00492] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00924] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00493] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00926] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00494] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00928] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00495] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0092a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00496] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0092c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00497] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0092e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00498] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00930] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00499] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00932] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0049a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00934] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0049b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00936] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0049c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00938] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0049d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0093a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0049e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0093c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0049f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0093e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00940] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00942] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00944] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00946] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00948] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0094a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0094c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0094e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00950] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00952] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00954] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00956] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00958] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0095a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0095c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0095e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00960] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00962] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00964] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00966] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00968] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0096a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0096c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0096e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00970] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00972] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00974] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00976] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00978] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0097a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0097c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0097e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00980] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00982] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00984] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00986] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00988] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0098a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0098c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0098e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00990] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00992] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00994] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00996] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00998] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0099a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0099c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0099e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h009fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00500] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00501] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00502] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00503] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00504] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00505] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00506] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00507] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00508] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00509] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0050a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0050b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0050c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0050d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0050e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0050f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00510] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00511] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00512] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00513] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00514] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00515] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00516] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00517] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00518] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00519] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0051a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0051b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0051c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0051d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0051e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0051f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00520] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00521] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00522] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00523] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00524] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00525] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00526] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00527] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00528] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00529] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0052a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0052b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0052c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0052d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0052e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0052f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00530] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00531] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00532] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00533] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00534] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00535] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00536] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00537] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00538] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00539] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0053a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0053b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0053c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0053d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0053e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0053f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00540] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00541] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00542] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00543] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00544] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00545] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00546] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00547] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00548] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00549] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0054a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0054b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0054c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0054d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0054e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0054f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00a9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00550] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00551] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00552] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00553] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00554] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00555] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00556] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00557] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00558] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ab0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00559] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ab2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0055a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ab4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0055b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ab6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0055c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ab8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0055d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0055e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00abc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0055f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00abe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00560] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ac0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00561] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ac2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00562] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ac4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00563] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ac6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00564] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ac8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00565] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00566] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00acc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00567] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ace] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00568] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ad0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00569] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ad2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0056a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ad4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0056b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ad6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0056c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ad8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0056d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ada] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0056e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00adc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0056f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ade] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00570] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ae0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00571] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ae2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00572] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ae4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00573] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ae6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00574] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ae8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00575] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00576] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00577] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00aee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00578] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00af0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00579] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00af2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0057a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00af4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0057b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00af6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0057c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00af8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0057d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00afa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0057e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00afc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0057f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00afe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00580] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00581] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00582] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00583] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00584] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00585] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00586] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00587] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00588] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00589] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0058a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0058b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0058c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0058d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0058e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0058f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00590] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00591] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00592] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00593] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00594] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00595] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00596] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00597] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00598] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00599] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0059a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0059b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0059c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0059d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0059e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0059f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00b9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ba0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ba2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ba4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ba6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ba8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00baa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00be0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00be2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00be4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00be6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00be8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00bfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00600] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00601] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00602] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00603] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00604] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00605] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00606] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00607] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00608] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00609] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0060a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0060b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0060c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0060d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0060e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0060f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00610] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00611] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00612] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00613] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00614] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00615] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00616] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00617] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00618] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00619] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0061a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0061b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0061c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0061d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0061e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0061f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00620] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00621] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00622] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00623] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00624] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00625] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00626] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00627] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00628] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00629] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0062a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0062b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0062c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0062d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0062e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0062f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00630] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00631] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00632] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00633] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00634] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00635] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00636] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00637] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00638] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00639] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0063a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0063b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0063c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0063d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0063e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0063f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00640] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00641] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00642] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00643] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00644] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00645] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00646] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00647] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00648] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00649] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0064a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0064b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0064c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0064d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0064e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0064f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00c9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00650] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ca0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00651] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ca2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00652] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ca4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00653] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ca6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00654] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ca8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00655] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00caa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00656] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00657] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00658] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00659] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0065a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0065b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0065c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0065d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0065e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0065f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00660] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00661] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00662] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00663] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00664] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00665] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00666] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ccc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00667] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00668] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00669] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0066a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0066b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0066c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0066d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0066e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0066f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00670] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ce0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00671] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ce2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00672] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ce4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00673] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ce6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00674] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ce8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00675] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00676] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00677] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00678] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00679] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0067a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0067b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0067c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0067d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0067e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0067f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00cfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00680] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00681] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00682] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00683] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00684] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00685] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00686] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00687] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00688] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00689] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0068a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0068b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0068c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0068d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0068e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0068f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00690] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00691] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00692] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00693] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00694] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00695] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00696] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00697] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00698] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00699] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0069a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0069b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0069c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0069d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0069e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0069f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00d9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00da0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00da2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00da4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00da6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00da8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00daa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00db0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00db2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00db4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00db6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00db8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ddc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00de0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00de2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00de4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00de6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00de8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00df0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00df2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00df4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00df6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00df8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00dfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00700] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00701] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00702] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00703] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00704] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00705] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00706] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00707] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00708] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00709] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0070a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0070b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0070c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0070d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0070e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0070f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00710] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00711] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00712] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00713] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00714] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00715] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00716] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00717] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00718] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00719] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0071a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0071b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0071c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0071d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0071e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0071f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00720] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00721] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00722] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00723] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00724] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00725] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00726] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00727] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00728] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00729] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0072a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0072b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0072c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0072d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0072e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0072f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00730] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00731] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00732] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00733] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00734] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00735] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00736] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00737] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00738] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00739] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0073a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0073b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0073c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0073d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0073e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0073f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00740] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00741] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00742] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00743] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00744] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00745] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00746] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00747] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00748] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00749] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0074a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0074b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0074c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0074d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0074e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0074f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00e9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00750] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ea0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00751] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ea2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00752] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ea4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00753] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ea6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00754] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ea8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00755] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00756] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00757] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00758] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00759] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0075a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0075b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0075c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0075d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0075e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ebc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0075f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ebe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00760] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ec0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00761] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ec2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00762] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ec4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00763] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ec6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00764] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ec8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00765] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00766] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ecc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00767] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ece] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00768] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ed0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00769] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ed2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0076a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ed4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0076b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ed6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0076c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ed8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0076d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0076e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00edc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0076f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ede] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00770] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ee0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00771] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ee2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00772] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ee4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00773] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ee6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00774] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ee8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00775] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00776] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00777] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00eee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00778] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ef0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00779] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ef2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0077a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ef4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0077b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ef6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0077c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ef8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0077d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00efa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0077e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00efc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0077f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00efe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00780] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00781] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00782] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00783] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00784] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00785] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00786] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00787] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00788] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00789] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0078a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0078b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0078c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0078d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0078e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0078f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00790] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00791] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00792] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00793] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00794] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00795] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00796] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00797] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00798] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00799] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0079a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0079b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0079c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0079d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0079e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0079f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00f9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00faa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fe0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fe2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fe4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fe6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fe8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00fee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ff0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ff2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ff4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ff6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ff8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ffa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ffc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h00ffe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00800] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01000] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00801] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01002] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00802] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01004] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00803] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01006] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00804] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01008] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00805] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0100a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00806] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0100c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00807] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0100e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00808] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01010] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00809] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01012] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0080a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01014] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0080b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01016] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0080c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01018] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0080d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0101a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0080e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0101c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0080f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0101e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00810] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01020] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00811] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01022] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00812] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01024] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00813] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01026] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00814] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01028] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00815] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0102a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00816] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0102c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00817] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0102e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00818] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01030] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00819] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01032] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0081a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01034] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0081b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01036] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0081c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01038] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0081d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0103a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0081e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0103c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0081f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0103e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00820] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01040] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00821] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01042] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00822] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01044] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00823] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01046] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00824] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01048] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00825] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0104a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00826] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0104c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00827] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0104e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00828] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01050] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00829] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01052] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0082a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01054] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0082b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01056] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0082c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01058] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0082d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0105a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0082e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0105c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0082f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0105e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00830] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01060] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00831] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01062] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00832] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01064] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00833] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01066] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00834] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01068] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00835] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0106a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00836] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0106c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00837] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0106e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00838] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01070] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00839] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01072] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0083a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01074] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0083b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01076] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0083c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01078] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0083d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0107a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0083e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0107c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0083f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0107e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00840] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01080] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00841] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01082] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00842] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01084] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00843] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01086] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00844] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01088] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00845] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0108a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00846] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0108c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00847] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0108e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00848] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01090] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00849] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01092] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0084a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01094] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0084b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01096] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0084c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01098] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0084d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0109a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0084e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0109c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0084f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0109e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00850] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00851] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00852] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00853] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00854] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00855] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00856] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00857] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00858] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00859] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0085a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0085b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0085c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0085d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0085e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0085f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00860] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00861] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00862] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00863] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00864] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00865] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00866] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00867] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00868] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00869] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0086a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0086b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0086c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0086d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0086e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0086f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00870] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00871] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00872] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00873] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00874] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00875] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00876] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00877] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00878] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00879] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0087a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0087b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0087c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0087d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0087e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0087f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h010fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00880] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01100] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00881] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01102] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00882] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01104] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00883] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01106] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00884] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01108] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00885] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0110a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00886] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0110c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00887] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0110e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00888] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01110] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00889] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01112] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0088a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01114] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0088b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01116] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0088c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01118] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0088d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0111a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0088e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0111c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0088f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0111e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00890] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01120] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00891] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01122] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00892] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01124] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00893] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01126] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00894] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01128] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00895] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0112a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00896] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0112c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00897] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0112e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00898] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01130] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00899] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01132] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0089a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01134] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0089b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01136] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0089c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01138] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0089d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0113a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0089e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0113c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0089f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0113e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01140] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01142] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01144] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01146] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01148] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0114a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0114c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0114e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01150] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01152] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01154] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01156] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01158] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0115a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0115c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0115e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01160] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01162] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01164] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01166] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01168] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0116a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0116c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0116e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01170] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01172] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01174] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01176] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01178] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0117a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0117c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0117e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01180] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01182] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01184] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01186] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01188] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0118a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0118c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0118e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01190] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01192] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01194] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01196] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01198] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0119a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0119c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0119e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h011fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00900] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01200] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00901] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01202] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00902] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01204] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00903] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01206] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00904] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01208] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00905] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0120a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00906] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0120c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00907] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0120e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00908] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01210] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00909] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01212] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0090a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01214] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0090b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01216] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0090c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01218] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0090d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0121a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0090e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0121c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0090f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0121e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00910] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01220] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00911] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01222] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00912] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01224] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00913] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01226] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00914] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01228] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00915] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0122a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00916] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0122c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00917] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0122e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00918] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01230] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00919] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01232] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0091a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01234] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0091b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01236] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0091c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01238] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0091d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0123a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0091e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0123c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0091f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0123e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00920] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01240] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00921] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01242] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00922] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01244] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00923] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01246] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00924] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01248] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00925] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0124a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00926] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0124c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00927] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0124e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00928] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01250] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00929] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01252] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0092a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01254] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0092b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01256] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0092c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01258] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0092d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0125a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0092e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0125c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0092f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0125e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00930] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01260] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00931] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01262] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00932] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01264] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00933] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01266] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00934] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01268] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00935] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0126a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00936] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0126c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00937] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0126e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00938] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01270] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00939] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01272] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0093a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01274] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0093b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01276] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0093c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01278] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0093d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0127a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0093e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0127c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0093f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0127e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00940] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01280] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00941] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01282] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00942] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01284] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00943] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01286] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00944] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01288] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00945] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0128a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00946] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0128c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00947] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0128e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00948] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01290] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00949] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01292] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0094a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01294] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0094b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01296] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0094c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01298] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0094d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0129a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0094e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0129c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0094f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0129e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00950] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00951] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00952] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00953] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00954] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00955] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00956] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00957] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00958] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00959] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0095a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0095b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0095c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0095d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0095e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0095f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00960] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00961] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00962] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00963] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00964] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00965] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00966] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00967] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00968] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00969] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0096a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0096b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0096c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0096d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0096e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0096f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00970] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00971] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00972] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00973] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00974] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00975] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00976] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00977] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00978] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00979] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0097a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0097b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0097c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0097d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0097e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0097f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h012fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00980] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01300] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00981] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01302] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00982] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01304] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00983] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01306] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00984] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01308] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00985] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0130a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00986] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0130c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00987] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0130e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00988] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01310] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00989] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01312] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0098a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01314] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0098b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01316] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0098c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01318] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0098d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0131a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0098e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0131c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0098f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0131e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00990] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01320] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00991] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01322] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00992] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01324] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00993] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01326] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00994] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01328] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00995] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0132a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00996] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0132c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00997] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0132e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00998] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01330] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00999] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01332] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0099a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01334] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0099b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01336] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0099c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01338] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0099d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0133a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0099e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0133c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0099f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0133e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01340] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01342] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01344] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01346] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01348] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0134a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0134c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0134e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01350] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01352] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01354] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01356] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01358] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0135a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0135c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0135e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01360] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01362] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01364] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01366] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01368] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0136a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0136c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0136e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01370] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01372] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01374] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01376] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01378] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0137a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0137c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0137e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01380] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01382] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01384] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01386] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01388] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0138a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0138c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0138e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01390] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01392] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01394] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01396] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01398] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0139a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0139c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0139e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h013fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01400] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01402] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01404] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01406] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01408] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0140a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0140c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0140e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01410] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01412] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01414] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01416] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01418] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0141a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0141c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0141e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01420] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01422] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01424] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01426] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01428] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0142a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0142c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0142e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01430] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01432] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01434] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01436] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01438] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0143a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0143c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0143e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01440] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01442] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01444] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01446] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01448] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0144a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0144c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0144e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01450] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01452] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01454] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01456] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01458] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0145a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0145c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0145e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01460] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01462] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01464] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01466] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01468] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0146a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0146c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0146e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01470] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01472] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01474] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01476] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01478] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0147a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0147c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0147e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01480] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01482] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01484] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01486] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01488] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0148a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0148c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0148e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01490] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01492] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01494] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01496] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01498] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0149a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0149c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0149e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h014fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01500] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01502] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01504] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01506] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01508] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0150a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0150c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0150e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01510] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01512] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01514] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01516] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01518] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0151a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0151c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0151e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01520] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01522] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01524] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01526] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01528] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0152a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0152c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0152e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01530] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01532] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01534] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01536] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01538] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0153a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0153c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0153e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01540] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01542] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01544] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01546] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01548] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0154a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0154c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0154e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01550] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01552] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aaa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01554] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01556] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01558] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0155a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0155c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aaf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0155e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01560] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01562] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01564] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01566] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01568] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0156a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0156c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0156e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01570] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01572] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01574] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00abb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01576] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00abc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01578] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00abd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0157a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00abe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0157c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00abf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0157e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01580] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01582] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01584] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01586] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01588] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0158a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0158c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0158e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01590] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01592] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01594] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00acb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01596] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00acc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01598] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00acd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0159a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ace] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0159c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00acf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0159e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ada] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00adb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00adc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00add] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ade] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00adf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aeb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00afa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00afb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00afc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00afd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00afe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h015fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01600] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01602] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01604] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01606] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01608] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0160a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0160c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0160e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01610] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01612] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01614] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01616] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01618] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0161a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0161c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0161e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01620] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01622] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01624] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01626] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01628] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0162a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0162c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0162e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01630] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01632] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01634] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01636] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01638] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0163a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0163c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0163e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01640] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01642] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01644] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01646] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01648] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0164a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0164c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0164e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01650] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01652] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01654] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01656] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01658] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0165a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0165c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0165e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01660] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01662] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01664] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01666] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01668] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0166a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0166c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0166e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01670] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01672] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01674] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01676] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01678] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0167a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0167c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0167e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01680] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01682] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01684] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01686] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01688] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0168a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0168c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0168e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01690] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01692] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01694] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01696] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01698] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0169a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0169c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0169e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h016fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01700] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01702] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01704] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01706] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01708] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0170a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0170c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0170e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01710] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01712] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01714] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01716] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01718] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0171a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0171c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0171e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01720] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01722] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01724] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01726] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01728] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0172a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0172c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0172e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01730] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01732] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01734] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01736] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01738] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0173a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0173c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0173e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01740] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01742] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01744] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01746] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01748] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0174a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0174c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0174e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01750] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01752] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00baa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01754] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01756] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01758] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0175a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0175c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00baf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0175e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01760] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01762] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01764] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01766] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01768] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0176a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0176c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0176e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01770] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01772] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01774] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01776] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01778] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0177a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0177c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0177e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01780] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01782] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01784] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01786] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01788] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0178a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0178c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0178e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01790] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01792] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01794] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01796] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01798] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0179a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0179c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0179e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00beb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h017fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01800] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01802] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01804] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01806] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01808] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0180a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0180c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0180e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01810] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01812] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01814] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01816] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01818] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0181a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0181c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0181e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01820] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01822] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01824] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01826] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01828] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0182a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0182c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0182e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01830] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01832] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01834] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01836] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01838] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0183a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0183c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0183e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01840] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01842] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01844] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01846] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01848] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0184a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0184c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0184e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01850] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01852] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01854] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01856] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01858] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0185a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0185c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0185e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01860] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01862] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01864] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01866] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01868] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0186a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0186c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0186e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01870] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01872] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01874] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01876] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01878] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0187a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0187c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0187e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01880] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01882] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01884] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01886] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01888] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0188a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0188c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0188e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01890] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01892] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01894] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01896] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01898] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0189a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0189c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0189e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h018fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01900] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01902] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01904] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01906] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01908] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0190a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0190c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0190e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01910] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01912] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01914] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01916] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01918] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0191a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0191c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0191e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01920] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01922] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01924] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01926] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01928] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0192a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0192c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0192e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01930] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01932] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01934] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01936] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01938] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0193a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0193c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0193e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01940] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01942] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01944] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01946] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01948] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0194a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0194c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0194e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01950] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01952] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00caa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01954] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01956] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01958] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0195a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0195c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00caf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0195e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01960] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01962] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01964] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01966] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01968] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0196a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0196c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0196e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01970] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01972] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01974] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01976] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01978] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0197a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0197c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0197e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01980] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01982] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01984] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01986] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01988] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0198a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0198c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0198e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01990] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01992] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01994] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ccb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01996] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ccc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01998] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ccd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0199a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0199c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ccf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0199e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ceb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ced] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h019fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01a9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ab0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ab2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ab4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ab6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ab8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01abc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01abe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ac0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ac2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ac4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ac6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ac8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01acc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ace] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ad0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ad2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ad4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ad6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ad8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ada] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01adc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ade] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ae0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ae2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ae4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ae6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ae8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01aee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01af0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01af2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01af4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01af6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01af8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01afa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01afc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01afe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00daa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00daf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01b9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ba0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ba2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ba4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ba6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ba8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01baa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ddb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ddc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ddd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ddf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00deb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ded] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00def] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01be0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01be2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01be4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01be6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01be8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01bfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01c9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ca0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ca2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ca4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ca6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ca8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01caa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ccc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ce0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ce2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ce4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ce6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ce8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01cfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eaa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ead] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eaf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ebb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ebc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ebd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ebe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ebf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ecb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ecc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ecd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ece] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ecf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01d9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01da0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01da2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01da4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01da6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01da8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01daa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01db0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01db2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01db4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00edb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01db6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00edc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01db8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00edd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ede] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00edf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eeb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ddc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01de0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01de2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01de4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01de6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01de8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01df0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01df2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00efa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01df4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00efb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01df6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00efc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01df8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00efd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00efe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01dfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01e9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ea0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ea2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ea4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ea6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ea8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ebc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ebe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ec0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ec2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ec4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ec6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ec8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ecc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ece] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ed0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ed2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ed4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ed6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ed8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01edc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ede] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ee0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ee2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ee4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ee6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ee8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01eee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ef0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ef2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ef4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ef6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ef8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01efa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01efc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01efe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00faa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00faf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01f9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01faa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00feb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fe0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fe2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fe4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fe6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fe8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01fee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ff0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ff2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ffa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ff4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ffb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ff6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ffc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ff8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ffd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ffa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ffe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ffc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h01ffe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01000] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02000] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01001] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02002] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01002] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02004] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01003] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02006] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01004] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02008] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01005] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0200a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01006] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0200c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01007] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0200e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01008] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02010] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01009] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02012] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0100a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02014] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0100b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02016] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0100c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02018] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0100d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0201a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0100e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0201c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0100f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0201e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01010] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02020] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01011] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02022] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01012] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02024] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01013] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02026] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01014] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02028] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01015] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0202a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01016] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0202c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01017] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0202e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01018] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02030] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01019] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02032] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0101a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02034] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0101b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02036] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0101c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02038] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0101d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0203a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0101e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0203c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0101f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0203e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01020] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02040] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01021] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02042] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01022] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02044] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01023] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02046] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01024] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02048] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01025] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0204a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01026] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0204c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01027] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0204e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01028] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02050] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01029] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02052] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0102a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02054] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0102b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02056] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0102c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02058] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0102d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0205a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0102e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0205c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0102f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0205e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01030] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02060] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01031] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02062] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01032] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02064] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01033] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02066] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01034] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02068] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01035] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0206a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01036] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0206c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01037] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0206e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01038] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02070] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01039] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02072] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0103a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02074] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0103b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02076] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0103c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02078] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0103d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0207a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0103e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0207c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0103f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0207e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01040] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02080] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01041] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02082] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01042] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02084] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01043] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02086] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01044] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02088] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01045] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0208a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01046] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0208c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01047] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0208e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01048] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02090] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01049] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02092] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0104a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02094] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0104b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02096] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0104c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02098] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0104d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0209a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0104e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0209c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0104f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0209e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01050] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01051] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01052] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01053] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01054] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01055] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01056] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01057] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01058] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01059] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0105a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0105b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0105c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0105d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0105e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0105f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01060] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01061] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01062] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01063] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01064] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01065] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01066] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01067] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01068] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01069] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0106a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0106b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0106c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0106d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0106e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0106f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01070] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01071] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01072] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01073] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01074] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01075] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01076] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01077] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01078] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01079] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0107a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0107b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0107c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0107d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0107e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0107f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h020fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01080] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02100] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01081] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02102] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01082] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02104] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01083] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02106] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01084] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02108] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01085] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0210a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01086] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0210c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01087] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0210e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01088] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02110] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01089] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02112] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0108a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02114] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0108b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02116] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0108c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02118] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0108d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0211a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0108e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0211c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0108f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0211e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01090] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02120] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01091] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02122] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01092] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02124] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01093] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02126] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01094] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02128] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01095] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0212a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01096] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0212c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01097] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0212e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01098] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02130] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01099] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02132] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0109a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02134] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0109b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02136] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0109c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02138] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0109d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0213a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0109e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0213c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0109f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0213e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02140] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02142] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02144] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02146] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02148] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0214a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0214c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0214e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02150] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02152] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02154] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02156] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02158] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0215a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0215c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0215e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02160] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02162] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02164] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02166] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02168] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0216a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0216c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0216e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02170] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02172] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02174] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02176] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02178] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0217a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0217c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0217e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02180] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02182] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02184] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02186] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02188] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0218a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0218c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0218e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02190] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02192] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02194] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02196] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02198] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0219a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0219c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0219e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h021fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01100] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02200] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01101] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02202] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01102] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02204] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01103] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02206] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01104] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02208] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01105] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0220a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01106] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0220c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01107] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0220e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01108] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02210] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01109] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02212] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0110a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02214] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0110b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02216] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0110c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02218] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0110d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0221a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0110e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0221c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0110f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0221e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01110] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02220] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01111] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02222] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01112] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02224] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01113] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02226] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01114] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02228] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01115] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0222a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01116] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0222c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01117] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0222e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01118] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02230] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01119] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02232] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0111a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02234] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0111b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02236] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0111c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02238] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0111d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0223a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0111e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0223c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0111f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0223e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01120] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02240] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01121] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02242] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01122] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02244] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01123] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02246] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01124] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02248] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01125] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0224a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01126] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0224c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01127] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0224e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01128] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02250] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01129] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02252] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0112a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02254] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0112b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02256] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0112c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02258] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0112d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0225a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0112e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0225c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0112f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0225e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01130] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02260] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01131] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02262] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01132] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02264] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01133] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02266] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01134] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02268] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01135] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0226a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01136] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0226c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01137] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0226e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01138] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02270] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01139] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02272] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0113a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02274] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0113b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02276] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0113c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02278] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0113d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0227a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0113e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0227c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0113f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0227e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01140] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02280] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01141] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02282] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01142] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02284] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01143] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02286] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01144] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02288] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01145] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0228a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01146] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0228c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01147] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0228e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01148] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02290] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01149] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02292] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0114a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02294] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0114b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02296] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0114c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02298] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0114d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0229a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0114e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0229c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0114f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0229e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01150] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01151] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01152] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01153] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01154] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01155] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01156] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01157] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01158] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01159] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0115a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0115b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0115c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0115d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0115e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0115f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01160] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01161] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01162] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01163] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01164] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01165] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01166] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01167] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01168] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01169] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0116a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0116b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0116c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0116d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0116e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0116f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01170] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01171] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01172] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01173] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01174] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01175] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01176] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01177] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01178] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01179] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0117a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0117b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0117c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0117d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0117e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0117f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h022fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01180] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02300] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01181] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02302] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01182] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02304] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01183] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02306] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01184] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02308] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01185] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0230a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01186] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0230c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01187] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0230e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01188] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02310] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01189] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02312] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0118a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02314] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0118b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02316] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0118c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02318] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0118d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0231a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0118e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0231c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0118f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0231e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01190] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02320] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01191] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02322] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01192] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02324] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01193] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02326] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01194] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02328] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01195] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0232a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01196] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0232c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01197] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0232e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01198] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02330] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01199] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02332] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0119a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02334] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0119b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02336] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0119c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02338] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0119d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0233a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0119e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0233c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0119f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0233e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02340] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02342] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02344] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02346] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02348] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0234a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0234c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0234e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02350] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02352] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02354] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02356] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02358] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0235a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0235c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0235e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02360] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02362] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02364] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02366] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02368] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0236a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0236c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0236e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02370] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02372] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02374] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02376] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02378] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0237a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0237c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0237e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02380] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02382] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02384] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02386] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02388] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0238a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0238c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0238e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02390] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02392] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02394] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02396] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02398] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0239a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0239c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0239e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h023fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01200] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02400] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01201] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02402] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01202] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02404] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01203] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02406] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01204] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02408] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01205] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0240a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01206] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0240c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01207] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0240e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01208] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02410] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01209] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02412] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0120a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02414] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0120b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02416] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0120c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02418] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0120d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0241a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0120e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0241c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0120f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0241e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01210] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02420] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01211] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02422] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01212] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02424] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01213] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02426] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01214] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02428] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01215] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0242a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01216] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0242c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01217] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0242e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01218] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02430] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01219] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02432] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0121a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02434] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0121b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02436] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0121c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02438] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0121d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0243a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0121e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0243c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0121f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0243e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01220] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02440] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01221] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02442] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01222] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02444] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01223] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02446] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01224] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02448] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01225] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0244a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01226] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0244c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01227] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0244e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01228] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02450] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01229] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02452] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0122a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02454] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0122b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02456] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0122c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02458] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0122d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0245a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0122e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0245c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0122f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0245e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01230] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02460] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01231] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02462] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01232] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02464] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01233] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02466] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01234] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02468] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01235] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0246a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01236] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0246c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01237] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0246e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01238] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02470] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01239] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02472] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0123a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02474] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0123b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02476] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0123c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02478] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0123d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0247a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0123e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0247c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0123f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0247e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01240] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02480] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01241] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02482] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01242] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02484] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01243] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02486] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01244] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02488] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01245] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0248a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01246] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0248c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01247] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0248e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01248] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02490] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01249] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02492] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0124a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02494] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0124b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02496] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0124c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02498] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0124d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0249a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0124e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0249c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0124f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0249e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01250] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01251] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01252] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01253] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01254] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01255] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01256] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01257] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01258] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01259] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0125a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0125b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0125c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0125d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0125e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0125f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01260] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01261] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01262] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01263] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01264] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01265] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01266] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01267] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01268] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01269] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0126a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0126b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0126c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0126d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0126e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0126f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01270] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01271] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01272] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01273] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01274] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01275] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01276] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01277] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01278] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01279] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0127a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0127b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0127c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0127d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0127e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0127f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h024fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01280] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02500] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01281] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02502] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01282] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02504] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01283] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02506] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01284] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02508] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01285] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0250a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01286] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0250c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01287] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0250e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01288] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02510] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01289] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02512] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0128a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02514] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0128b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02516] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0128c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02518] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0128d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0251a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0128e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0251c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0128f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0251e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01290] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02520] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01291] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02522] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01292] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02524] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01293] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02526] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01294] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02528] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01295] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0252a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01296] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0252c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01297] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0252e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01298] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02530] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01299] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02532] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0129a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02534] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0129b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02536] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0129c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02538] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0129d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0253a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0129e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0253c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0129f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0253e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02540] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02542] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02544] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02546] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02548] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0254a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0254c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0254e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02550] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02552] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02554] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02556] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02558] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0255a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0255c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0255e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02560] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02562] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02564] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02566] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02568] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0256a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0256c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0256e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02570] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02572] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02574] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02576] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02578] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0257a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0257c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0257e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02580] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02582] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02584] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02586] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02588] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0258a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0258c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0258e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02590] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02592] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02594] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02596] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02598] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0259a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0259c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0259e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h025fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01300] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02600] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01301] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02602] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01302] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02604] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01303] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02606] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01304] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02608] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01305] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0260a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01306] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0260c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01307] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0260e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01308] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02610] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01309] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02612] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0130a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02614] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0130b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02616] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0130c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02618] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0130d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0261a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0130e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0261c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0130f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0261e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01310] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02620] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01311] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02622] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01312] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02624] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01313] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02626] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01314] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02628] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01315] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0262a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01316] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0262c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01317] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0262e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01318] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02630] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01319] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02632] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0131a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02634] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0131b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02636] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0131c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02638] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0131d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0263a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0131e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0263c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0131f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0263e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01320] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02640] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01321] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02642] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01322] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02644] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01323] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02646] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01324] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02648] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01325] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0264a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01326] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0264c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01327] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0264e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01328] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02650] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01329] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02652] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0132a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02654] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0132b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02656] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0132c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02658] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0132d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0265a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0132e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0265c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0132f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0265e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01330] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02660] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01331] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02662] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01332] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02664] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01333] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02666] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01334] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02668] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01335] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0266a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01336] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0266c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01337] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0266e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01338] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02670] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01339] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02672] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0133a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02674] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0133b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02676] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0133c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02678] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0133d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0267a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0133e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0267c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0133f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0267e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01340] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02680] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01341] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02682] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01342] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02684] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01343] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02686] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01344] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02688] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01345] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0268a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01346] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0268c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01347] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0268e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01348] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02690] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01349] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02692] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0134a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02694] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0134b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02696] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0134c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02698] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0134d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0269a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0134e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0269c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0134f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0269e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01350] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01351] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01352] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01353] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01354] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01355] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01356] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01357] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01358] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01359] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0135a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0135b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0135c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0135d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0135e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0135f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01360] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01361] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01362] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01363] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01364] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01365] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01366] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01367] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01368] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01369] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0136a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0136b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0136c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0136d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0136e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0136f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01370] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01371] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01372] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01373] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01374] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01375] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01376] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01377] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01378] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01379] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0137a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0137b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0137c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0137d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0137e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0137f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h026fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01380] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02700] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01381] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02702] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01382] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02704] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01383] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02706] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01384] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02708] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01385] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0270a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01386] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0270c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01387] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0270e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01388] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02710] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01389] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02712] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0138a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02714] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0138b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02716] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0138c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02718] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0138d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0271a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0138e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0271c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0138f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0271e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01390] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02720] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01391] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02722] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01392] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02724] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01393] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02726] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01394] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02728] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01395] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0272a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01396] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0272c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01397] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0272e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01398] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02730] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01399] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02732] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0139a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02734] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0139b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02736] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0139c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02738] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0139d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0273a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0139e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0273c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0139f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0273e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02740] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02742] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02744] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02746] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02748] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0274a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0274c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0274e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02750] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02752] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02754] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02756] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02758] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0275a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0275c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0275e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02760] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02762] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02764] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02766] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02768] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0276a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0276c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0276e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02770] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02772] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02774] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02776] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02778] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0277a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0277c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0277e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02780] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02782] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02784] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02786] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02788] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0278a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0278c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0278e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02790] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02792] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02794] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02796] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02798] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0279a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0279c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0279e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h027fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01400] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02800] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01401] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02802] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01402] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02804] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01403] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02806] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01404] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02808] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01405] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0280a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01406] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0280c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01407] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0280e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01408] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02810] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01409] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02812] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0140a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02814] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0140b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02816] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0140c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02818] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0140d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0281a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0140e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0281c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0140f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0281e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01410] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02820] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01411] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02822] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01412] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02824] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01413] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02826] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01414] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02828] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01415] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0282a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01416] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0282c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01417] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0282e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01418] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02830] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01419] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02832] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0141a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02834] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0141b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02836] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0141c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02838] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0141d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0283a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0141e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0283c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0141f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0283e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01420] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02840] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01421] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02842] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01422] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02844] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01423] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02846] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01424] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02848] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01425] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0284a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01426] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0284c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01427] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0284e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01428] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02850] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01429] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02852] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0142a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02854] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0142b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02856] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0142c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02858] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0142d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0285a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0142e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0285c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0142f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0285e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01430] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02860] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01431] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02862] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01432] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02864] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01433] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02866] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01434] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02868] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01435] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0286a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01436] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0286c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01437] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0286e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01438] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02870] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01439] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02872] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0143a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02874] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0143b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02876] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0143c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02878] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0143d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0287a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0143e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0287c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0143f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0287e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01440] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02880] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01441] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02882] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01442] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02884] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01443] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02886] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01444] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02888] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01445] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0288a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01446] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0288c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01447] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0288e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01448] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02890] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01449] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02892] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0144a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02894] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0144b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02896] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0144c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02898] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0144d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0289a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0144e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0289c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0144f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0289e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01450] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01451] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01452] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01453] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01454] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01455] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01456] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01457] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01458] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01459] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0145a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0145b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0145c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0145d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0145e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0145f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01460] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01461] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01462] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01463] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01464] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01465] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01466] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01467] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01468] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01469] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0146a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0146b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0146c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0146d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0146e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0146f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01470] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01471] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01472] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01473] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01474] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01475] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01476] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01477] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01478] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01479] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0147a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0147b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0147c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0147d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0147e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0147f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h028fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01480] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02900] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01481] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02902] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01482] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02904] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01483] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02906] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01484] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02908] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01485] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0290a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01486] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0290c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01487] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0290e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01488] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02910] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01489] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02912] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0148a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02914] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0148b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02916] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0148c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02918] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0148d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0291a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0148e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0291c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0148f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0291e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01490] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02920] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01491] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02922] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01492] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02924] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01493] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02926] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01494] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02928] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01495] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0292a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01496] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0292c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01497] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0292e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01498] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02930] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01499] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02932] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0149a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02934] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0149b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02936] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0149c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02938] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0149d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0293a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0149e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0293c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0149f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0293e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02940] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02942] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02944] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02946] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02948] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0294a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0294c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0294e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02950] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02952] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02954] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02956] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02958] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0295a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0295c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0295e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02960] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02962] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02964] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02966] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02968] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0296a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0296c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0296e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02970] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02972] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02974] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02976] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02978] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0297a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0297c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0297e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02980] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02982] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02984] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02986] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02988] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0298a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0298c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0298e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02990] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02992] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02994] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02996] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02998] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0299a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0299c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0299e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h029fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01500] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01501] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01502] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01503] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01504] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01505] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01506] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01507] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01508] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01509] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0150a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0150b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0150c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0150d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0150e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0150f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01510] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01511] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01512] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01513] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01514] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01515] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01516] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01517] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01518] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01519] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0151a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0151b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0151c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0151d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0151e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0151f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01520] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01521] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01522] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01523] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01524] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01525] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01526] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01527] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01528] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01529] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0152a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0152b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0152c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0152d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0152e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0152f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01530] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01531] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01532] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01533] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01534] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01535] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01536] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01537] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01538] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01539] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0153a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0153b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0153c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0153d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0153e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0153f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01540] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01541] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01542] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01543] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01544] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01545] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01546] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01547] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01548] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01549] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0154a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0154b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0154c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0154d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0154e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0154f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02a9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01550] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01551] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01552] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01553] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01554] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01555] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01556] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01557] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01558] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ab0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01559] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ab2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0155a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ab4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0155b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ab6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0155c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ab8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0155d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0155e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02abc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0155f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02abe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01560] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ac0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01561] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ac2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01562] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ac4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01563] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ac6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01564] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ac8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01565] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01566] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02acc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01567] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ace] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01568] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ad0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01569] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ad2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0156a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ad4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0156b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ad6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0156c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ad8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0156d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ada] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0156e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02adc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0156f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ade] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01570] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ae0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01571] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ae2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01572] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ae4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01573] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ae6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01574] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ae8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01575] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01576] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01577] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02aee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01578] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02af0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01579] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02af2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0157a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02af4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0157b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02af6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0157c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02af8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0157d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02afa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0157e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02afc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0157f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02afe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01580] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01581] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01582] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01583] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01584] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01585] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01586] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01587] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01588] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01589] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0158a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0158b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0158c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0158d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0158e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0158f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01590] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01591] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01592] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01593] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01594] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01595] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01596] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01597] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01598] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01599] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0159a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0159b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0159c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0159d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0159e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0159f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02b9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ba0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ba2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ba4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ba6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ba8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02baa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02be0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02be2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02be4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02be6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02be8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02bfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01600] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01601] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01602] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01603] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01604] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01605] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01606] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01607] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01608] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01609] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0160a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0160b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0160c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0160d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0160e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0160f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01610] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01611] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01612] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01613] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01614] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01615] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01616] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01617] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01618] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01619] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0161a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0161b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0161c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0161d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0161e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0161f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01620] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01621] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01622] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01623] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01624] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01625] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01626] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01627] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01628] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01629] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0162a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0162b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0162c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0162d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0162e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0162f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01630] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01631] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01632] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01633] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01634] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01635] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01636] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01637] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01638] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01639] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0163a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0163b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0163c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0163d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0163e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0163f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01640] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01641] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01642] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01643] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01644] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01645] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01646] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01647] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01648] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01649] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0164a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0164b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0164c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0164d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0164e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0164f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02c9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01650] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ca0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01651] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ca2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01652] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ca4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01653] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ca6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01654] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ca8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01655] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02caa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01656] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01657] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01658] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01659] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0165a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0165b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0165c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0165d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0165e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0165f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01660] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01661] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01662] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01663] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01664] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01665] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01666] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ccc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01667] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01668] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01669] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0166a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0166b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0166c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0166d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0166e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0166f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01670] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ce0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01671] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ce2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01672] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ce4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01673] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ce6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01674] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ce8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01675] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01676] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01677] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01678] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01679] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0167a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0167b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0167c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0167d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0167e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0167f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02cfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01680] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01681] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01682] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01683] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01684] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01685] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01686] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01687] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01688] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01689] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0168a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0168b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0168c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0168d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0168e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0168f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01690] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01691] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01692] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01693] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01694] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01695] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01696] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01697] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01698] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01699] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0169a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0169b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0169c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0169d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0169e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0169f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02d9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02da0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02da2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02da4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02da6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02da8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02daa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02db0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02db2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02db4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02db6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02db8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ddc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02de0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02de2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02de4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02de6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02de8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02df0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02df2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02df4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02df6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02df8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02dfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01700] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01701] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01702] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01703] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01704] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01705] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01706] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01707] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01708] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01709] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0170a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0170b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0170c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0170d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0170e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0170f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01710] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01711] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01712] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01713] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01714] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01715] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01716] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01717] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01718] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01719] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0171a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0171b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0171c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0171d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0171e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0171f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01720] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01721] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01722] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01723] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01724] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01725] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01726] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01727] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01728] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01729] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0172a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0172b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0172c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0172d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0172e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0172f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01730] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01731] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01732] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01733] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01734] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01735] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01736] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01737] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01738] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01739] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0173a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0173b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0173c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0173d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0173e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0173f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01740] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01741] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01742] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01743] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01744] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01745] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01746] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01747] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01748] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01749] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0174a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0174b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0174c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0174d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0174e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0174f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02e9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01750] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ea0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01751] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ea2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01752] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ea4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01753] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ea6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01754] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ea8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01755] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01756] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01757] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01758] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01759] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0175a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0175b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0175c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0175d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0175e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ebc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0175f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ebe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01760] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ec0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01761] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ec2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01762] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ec4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01763] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ec6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01764] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ec8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01765] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01766] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ecc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01767] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ece] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01768] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ed0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01769] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ed2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0176a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ed4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0176b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ed6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0176c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ed8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0176d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0176e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02edc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0176f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ede] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01770] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ee0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01771] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ee2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01772] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ee4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01773] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ee6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01774] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ee8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01775] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01776] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01777] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02eee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01778] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ef0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01779] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ef2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0177a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ef4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0177b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ef6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0177c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ef8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0177d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02efa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0177e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02efc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0177f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02efe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01780] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01781] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01782] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01783] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01784] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01785] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01786] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01787] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01788] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01789] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0178a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0178b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0178c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0178d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0178e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0178f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01790] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01791] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01792] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01793] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01794] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01795] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01796] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01797] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01798] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01799] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0179a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0179b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0179c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0179d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0179e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0179f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02f9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02faa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fe0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fe2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fe4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fe6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fe8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02fee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ff0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ff2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ff4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ff6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ff8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ffa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ffc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h02ffe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01800] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03000] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01801] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03002] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01802] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03004] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01803] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03006] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01804] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03008] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01805] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0300a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01806] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0300c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01807] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0300e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01808] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03010] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01809] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03012] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0180a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03014] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0180b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03016] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0180c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03018] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0180d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0301a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0180e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0301c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0180f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0301e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01810] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03020] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01811] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03022] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01812] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03024] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01813] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03026] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01814] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03028] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01815] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0302a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01816] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0302c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01817] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0302e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01818] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03030] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01819] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03032] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0181a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03034] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0181b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03036] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0181c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03038] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0181d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0303a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0181e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0303c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0181f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0303e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01820] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03040] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01821] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03042] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01822] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03044] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01823] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03046] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01824] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03048] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01825] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0304a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01826] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0304c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01827] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0304e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01828] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03050] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01829] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03052] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0182a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03054] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0182b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03056] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0182c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03058] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0182d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0305a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0182e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0305c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0182f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0305e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01830] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03060] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01831] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03062] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01832] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03064] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01833] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03066] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01834] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03068] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01835] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0306a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01836] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0306c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01837] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0306e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01838] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03070] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01839] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03072] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0183a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03074] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0183b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03076] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0183c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03078] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0183d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0307a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0183e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0307c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0183f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0307e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01840] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03080] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01841] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03082] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01842] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03084] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01843] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03086] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01844] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03088] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01845] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0308a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01846] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0308c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01847] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0308e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01848] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03090] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01849] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03092] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0184a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03094] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0184b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03096] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0184c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03098] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0184d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0309a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0184e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0309c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0184f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0309e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01850] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01851] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01852] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01853] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01854] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01855] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01856] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01857] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01858] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01859] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0185a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0185b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0185c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0185d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0185e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0185f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01860] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01861] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01862] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01863] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01864] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01865] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01866] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01867] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01868] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01869] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0186a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0186b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0186c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0186d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0186e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0186f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01870] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01871] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01872] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01873] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01874] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01875] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01876] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01877] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01878] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01879] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0187a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0187b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0187c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0187d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0187e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0187f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h030fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01880] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03100] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01881] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03102] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01882] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03104] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01883] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03106] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01884] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03108] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01885] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0310a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01886] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0310c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01887] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0310e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01888] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03110] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01889] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03112] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0188a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03114] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0188b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03116] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0188c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03118] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0188d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0311a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0188e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0311c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0188f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0311e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01890] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03120] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01891] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03122] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01892] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03124] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01893] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03126] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01894] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03128] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01895] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0312a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01896] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0312c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01897] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0312e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01898] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03130] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01899] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03132] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0189a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03134] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0189b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03136] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0189c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03138] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0189d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0313a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0189e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0313c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0189f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0313e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03140] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03142] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03144] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03146] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03148] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0314a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0314c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0314e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03150] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03152] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03154] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03156] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03158] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0315a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0315c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0315e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03160] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03162] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03164] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03166] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03168] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0316a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0316c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0316e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03170] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03172] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03174] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03176] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03178] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0317a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0317c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0317e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03180] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03182] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03184] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03186] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03188] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0318a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0318c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0318e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03190] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03192] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03194] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03196] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03198] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0319a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0319c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0319e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h031fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01900] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03200] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01901] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03202] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01902] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03204] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01903] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03206] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01904] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03208] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01905] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0320a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01906] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0320c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01907] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0320e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01908] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03210] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01909] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03212] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0190a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03214] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0190b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03216] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0190c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03218] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0190d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0321a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0190e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0321c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0190f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0321e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01910] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03220] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01911] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03222] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01912] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03224] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01913] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03226] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01914] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03228] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01915] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0322a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01916] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0322c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01917] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0322e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01918] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03230] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01919] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03232] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0191a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03234] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0191b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03236] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0191c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03238] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0191d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0323a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0191e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0323c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0191f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0323e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01920] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03240] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01921] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03242] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01922] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03244] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01923] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03246] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01924] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03248] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01925] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0324a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01926] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0324c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01927] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0324e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01928] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03250] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01929] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03252] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0192a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03254] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0192b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03256] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0192c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03258] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0192d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0325a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0192e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0325c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0192f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0325e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01930] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03260] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01931] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03262] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01932] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03264] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01933] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03266] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01934] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03268] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01935] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0326a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01936] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0326c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01937] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0326e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01938] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03270] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01939] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03272] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0193a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03274] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0193b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03276] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0193c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03278] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0193d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0327a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0193e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0327c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0193f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0327e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01940] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03280] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01941] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03282] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01942] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03284] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01943] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03286] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01944] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03288] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01945] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0328a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01946] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0328c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01947] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0328e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01948] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03290] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01949] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03292] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0194a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03294] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0194b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03296] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0194c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03298] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0194d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0329a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0194e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0329c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0194f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0329e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01950] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01951] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01952] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01953] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01954] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01955] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01956] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01957] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01958] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01959] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0195a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0195b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0195c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0195d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0195e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0195f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01960] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01961] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01962] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01963] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01964] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01965] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01966] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01967] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01968] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01969] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0196a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0196b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0196c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0196d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0196e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0196f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01970] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01971] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01972] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01973] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01974] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01975] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01976] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01977] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01978] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01979] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0197a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0197b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0197c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0197d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0197e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0197f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h032fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01980] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03300] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01981] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03302] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01982] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03304] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01983] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03306] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01984] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03308] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01985] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0330a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01986] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0330c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01987] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0330e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01988] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03310] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01989] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03312] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0198a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03314] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0198b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03316] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0198c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03318] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0198d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0331a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0198e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0331c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0198f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0331e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01990] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03320] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01991] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03322] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01992] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03324] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01993] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03326] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01994] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03328] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01995] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0332a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01996] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0332c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01997] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0332e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01998] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03330] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01999] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03332] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0199a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03334] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0199b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03336] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0199c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03338] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0199d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0333a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0199e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0333c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0199f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0333e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03340] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03342] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03344] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03346] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03348] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0334a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0334c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0334e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03350] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03352] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03354] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03356] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03358] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0335a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0335c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0335e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03360] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03362] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03364] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03366] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03368] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0336a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0336c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0336e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03370] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03372] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03374] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03376] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03378] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0337a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0337c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0337e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03380] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03382] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03384] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03386] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03388] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0338a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0338c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0338e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03390] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03392] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03394] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03396] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03398] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0339a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0339c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0339e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h033fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03400] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03402] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03404] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03406] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03408] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0340a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0340c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0340e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03410] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03412] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03414] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03416] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03418] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0341a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0341c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0341e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03420] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03422] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03424] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03426] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03428] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0342a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0342c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0342e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03430] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03432] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03434] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03436] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03438] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0343a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0343c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0343e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03440] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03442] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03444] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03446] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03448] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0344a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0344c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0344e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03450] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03452] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03454] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03456] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03458] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0345a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0345c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0345e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03460] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03462] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03464] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03466] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03468] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0346a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0346c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0346e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03470] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03472] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03474] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03476] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03478] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0347a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0347c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0347e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03480] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03482] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03484] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03486] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03488] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0348a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0348c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0348e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03490] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03492] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03494] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03496] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03498] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0349a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0349c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0349e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h034fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03500] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03502] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03504] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03506] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03508] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0350a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0350c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0350e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03510] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03512] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03514] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03516] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03518] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0351a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0351c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0351e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03520] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03522] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03524] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03526] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03528] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0352a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0352c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0352e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03530] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03532] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03534] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03536] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03538] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0353a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0353c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0353e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03540] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03542] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03544] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03546] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03548] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0354a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0354c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0354e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03550] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03552] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aaa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03554] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03556] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03558] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0355a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0355c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aaf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0355e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03560] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03562] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03564] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03566] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03568] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0356a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0356c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0356e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03570] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03572] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03574] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01abb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03576] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01abc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03578] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01abd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0357a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01abe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0357c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01abf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0357e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03580] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03582] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03584] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03586] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03588] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0358a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0358c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0358e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03590] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03592] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03594] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01acb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03596] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01acc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03598] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01acd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0359a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ace] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0359c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01acf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0359e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ada] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01adb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01adc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01add] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ade] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01adf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aeb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01afa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01afb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01afc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01afd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01afe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h035fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03600] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03602] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03604] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03606] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03608] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0360a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0360c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0360e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03610] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03612] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03614] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03616] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03618] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0361a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0361c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0361e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03620] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03622] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03624] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03626] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03628] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0362a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0362c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0362e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03630] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03632] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03634] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03636] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03638] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0363a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0363c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0363e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03640] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03642] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03644] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03646] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03648] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0364a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0364c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0364e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03650] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03652] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03654] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03656] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03658] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0365a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0365c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0365e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03660] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03662] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03664] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03666] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03668] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0366a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0366c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0366e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03670] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03672] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03674] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03676] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03678] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0367a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0367c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0367e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03680] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03682] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03684] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03686] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03688] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0368a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0368c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0368e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03690] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03692] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03694] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03696] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03698] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0369a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0369c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0369e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h036fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03700] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03702] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03704] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03706] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03708] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0370a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0370c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0370e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03710] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03712] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03714] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03716] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03718] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0371a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0371c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0371e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03720] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03722] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03724] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03726] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03728] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0372a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0372c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0372e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03730] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03732] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03734] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03736] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03738] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0373a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0373c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0373e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03740] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03742] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03744] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03746] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03748] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0374a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0374c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0374e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03750] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03752] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01baa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03754] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03756] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03758] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0375a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0375c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01baf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0375e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03760] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03762] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03764] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03766] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03768] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0376a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0376c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0376e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03770] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03772] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03774] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03776] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03778] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0377a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0377c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0377e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03780] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03782] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03784] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03786] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03788] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0378a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0378c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0378e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03790] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03792] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03794] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03796] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03798] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0379a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0379c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0379e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01beb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h037fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03800] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03802] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03804] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03806] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03808] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0380a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0380c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0380e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03810] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03812] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03814] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03816] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03818] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0381a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0381c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0381e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03820] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03822] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03824] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03826] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03828] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0382a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0382c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0382e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03830] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03832] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03834] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03836] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03838] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0383a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0383c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0383e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03840] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03842] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03844] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03846] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03848] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0384a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0384c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0384e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03850] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03852] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03854] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03856] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03858] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0385a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0385c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0385e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03860] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03862] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03864] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03866] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03868] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0386a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0386c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0386e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03870] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03872] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03874] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03876] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03878] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0387a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0387c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0387e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03880] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03882] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03884] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03886] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03888] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0388a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0388c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0388e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03890] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03892] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03894] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03896] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03898] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0389a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0389c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0389e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h038fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03900] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03902] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03904] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03906] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03908] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0390a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0390c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0390e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03910] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03912] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03914] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03916] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03918] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0391a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0391c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0391e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03920] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03922] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03924] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03926] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03928] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0392a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0392c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0392e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03930] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03932] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03934] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03936] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03938] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0393a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0393c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0393e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03940] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03942] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03944] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03946] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03948] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0394a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0394c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0394e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03950] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03952] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01caa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03954] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03956] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03958] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0395a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0395c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01caf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0395e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03960] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03962] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03964] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03966] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03968] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0396a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0396c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0396e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03970] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03972] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03974] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03976] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03978] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0397a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0397c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0397e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03980] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03982] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03984] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03986] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03988] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0398a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0398c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0398e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03990] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03992] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03994] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ccb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03996] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ccc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03998] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ccd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0399a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0399c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ccf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0399e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ceb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ced] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h039fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03a9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ab0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ab2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ab4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ab6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ab8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03abc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03abe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ac0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ac2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ac4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ac6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ac8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03acc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ace] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ad0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ad2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ad4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ad6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ad8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ada] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03adc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ade] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ae0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ae2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ae4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ae6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ae8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03aee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03af0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03af2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03af4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03af6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03af8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03afa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03afc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03afe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01daa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01daf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03b9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ba0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ba2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ba4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ba6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ba8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03baa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ddb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ddc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ddd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ddf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01deb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ded] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01def] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03be0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03be2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03be4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03be6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03be8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03bfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03c9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ca0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ca2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ca4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ca6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ca8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03caa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ccc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ce0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ce2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ce4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ce6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ce8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03cfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eaa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ead] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eaf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ebb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ebc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ebd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ebe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ebf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ecb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ecc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ecd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ece] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ecf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03d9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03da0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03da2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03da4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03da6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03da8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03daa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03db0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03db2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03db4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01edb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03db6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01edc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03db8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01edd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ede] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01edf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eeb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ddc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03de0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03de2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03de4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03de6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03de8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03df0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03df2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01efa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03df4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01efb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03df6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01efc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03df8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01efd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01efe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03dfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03e9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ea0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ea2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ea4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ea6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ea8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ebc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ebe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ec0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ec2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ec4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ec6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ec8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ecc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ece] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ed0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ed2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ed4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ed6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ed8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03edc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ede] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ee0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ee2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ee4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ee6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ee8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03eee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ef0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ef2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ef4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ef6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ef8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03efa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03efc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03efe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01faa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01faf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03f9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03faa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01feb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fe0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fe2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fe4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fe6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fe8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03fee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ff0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ff2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ffa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ff4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ffb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ff6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ffc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ff8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ffd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ffa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ffe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ffc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h03ffe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02000] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04000] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02001] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04002] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02002] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04004] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02003] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04006] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02004] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04008] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02005] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0400a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02006] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0400c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02007] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0400e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02008] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04010] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02009] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04012] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0200a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04014] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0200b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04016] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0200c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04018] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0200d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0401a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0200e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0401c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0200f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0401e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02010] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04020] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02011] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04022] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02012] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04024] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02013] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04026] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02014] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04028] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02015] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0402a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02016] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0402c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02017] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0402e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02018] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04030] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02019] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04032] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0201a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04034] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0201b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04036] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0201c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04038] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0201d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0403a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0201e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0403c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0201f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0403e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02020] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04040] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02021] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04042] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02022] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04044] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02023] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04046] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02024] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04048] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02025] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0404a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02026] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0404c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02027] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0404e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02028] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04050] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02029] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04052] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0202a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04054] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0202b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04056] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0202c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04058] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0202d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0405a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0202e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0405c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0202f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0405e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02030] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04060] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02031] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04062] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02032] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04064] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02033] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04066] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02034] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04068] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02035] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0406a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02036] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0406c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02037] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0406e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02038] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04070] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02039] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04072] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0203a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04074] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0203b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04076] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0203c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04078] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0203d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0407a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0203e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0407c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0203f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0407e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02040] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04080] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02041] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04082] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02042] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04084] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02043] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04086] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02044] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04088] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02045] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0408a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02046] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0408c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02047] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0408e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02048] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04090] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02049] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04092] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0204a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04094] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0204b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04096] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0204c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04098] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0204d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0409a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0204e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0409c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0204f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0409e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02050] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02051] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02052] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02053] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02054] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02055] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02056] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02057] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02058] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02059] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0205a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0205b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0205c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0205d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0205e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0205f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02060] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02061] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02062] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02063] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02064] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02065] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02066] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02067] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02068] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02069] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0206a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0206b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0206c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0206d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0206e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0206f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02070] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02071] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02072] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02073] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02074] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02075] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02076] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02077] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02078] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02079] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0207a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0207b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0207c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0207d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0207e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0207f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h040fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02080] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04100] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02081] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04102] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02082] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04104] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02083] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04106] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02084] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04108] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02085] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0410a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02086] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0410c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02087] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0410e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02088] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04110] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02089] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04112] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0208a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04114] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0208b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04116] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0208c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04118] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0208d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0411a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0208e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0411c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0208f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0411e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02090] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04120] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02091] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04122] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02092] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04124] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02093] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04126] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02094] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04128] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02095] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0412a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02096] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0412c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02097] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0412e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02098] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04130] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02099] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04132] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0209a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04134] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0209b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04136] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0209c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04138] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0209d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0413a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0209e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0413c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0209f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0413e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04140] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04142] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04144] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04146] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04148] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0414a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0414c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0414e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04150] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04152] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04154] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04156] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04158] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0415a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0415c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0415e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04160] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04162] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04164] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04166] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04168] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0416a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0416c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0416e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04170] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04172] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04174] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04176] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04178] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0417a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0417c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0417e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04180] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04182] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04184] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04186] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04188] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0418a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0418c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0418e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04190] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04192] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04194] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04196] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04198] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0419a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0419c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0419e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h041fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02100] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04200] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02101] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04202] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02102] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04204] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02103] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04206] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02104] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04208] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02105] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0420a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02106] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0420c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02107] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0420e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02108] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04210] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02109] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04212] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0210a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04214] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0210b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04216] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0210c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04218] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0210d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0421a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0210e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0421c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0210f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0421e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02110] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04220] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02111] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04222] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02112] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04224] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02113] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04226] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02114] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04228] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02115] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0422a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02116] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0422c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02117] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0422e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02118] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04230] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02119] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04232] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0211a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04234] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0211b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04236] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0211c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04238] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0211d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0423a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0211e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0423c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0211f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0423e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02120] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04240] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02121] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04242] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02122] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04244] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02123] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04246] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02124] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04248] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02125] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0424a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02126] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0424c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02127] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0424e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02128] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04250] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02129] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04252] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0212a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04254] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0212b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04256] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0212c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04258] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0212d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0425a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0212e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0425c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0212f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0425e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02130] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04260] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02131] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04262] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02132] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04264] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02133] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04266] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02134] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04268] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02135] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0426a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02136] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0426c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02137] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0426e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02138] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04270] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02139] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04272] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0213a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04274] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0213b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04276] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0213c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04278] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0213d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0427a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0213e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0427c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0213f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0427e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02140] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04280] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02141] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04282] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02142] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04284] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02143] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04286] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02144] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04288] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02145] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0428a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02146] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0428c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02147] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0428e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02148] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04290] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02149] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04292] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0214a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04294] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0214b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04296] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0214c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04298] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0214d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0429a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0214e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0429c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0214f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0429e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02150] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02151] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02152] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02153] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02154] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02155] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02156] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02157] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02158] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02159] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0215a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0215b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0215c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0215d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0215e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0215f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02160] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02161] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02162] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02163] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02164] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02165] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02166] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02167] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02168] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02169] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0216a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0216b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0216c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0216d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0216e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0216f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02170] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02171] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02172] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02173] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02174] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02175] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02176] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02177] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02178] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02179] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0217a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0217b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0217c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0217d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0217e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0217f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h042fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02180] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04300] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02181] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04302] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02182] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04304] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02183] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04306] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02184] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04308] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02185] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0430a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02186] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0430c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02187] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0430e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02188] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04310] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02189] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04312] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0218a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04314] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0218b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04316] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0218c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04318] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0218d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0431a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0218e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0431c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0218f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0431e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02190] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04320] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02191] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04322] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02192] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04324] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02193] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04326] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02194] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04328] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02195] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0432a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02196] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0432c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02197] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0432e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02198] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04330] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02199] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04332] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0219a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04334] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0219b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04336] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0219c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04338] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0219d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0433a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0219e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0433c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0219f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0433e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04340] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04342] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04344] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04346] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04348] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0434a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0434c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0434e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04350] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04352] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04354] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04356] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04358] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0435a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0435c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0435e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04360] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04362] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04364] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04366] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04368] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0436a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0436c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0436e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04370] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04372] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04374] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04376] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04378] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0437a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0437c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0437e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04380] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04382] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04384] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04386] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04388] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0438a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0438c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0438e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04390] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04392] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04394] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04396] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04398] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0439a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0439c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0439e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h043fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02200] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04400] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02201] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04402] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02202] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04404] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02203] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04406] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02204] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04408] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02205] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0440a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02206] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0440c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02207] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0440e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02208] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04410] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02209] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04412] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0220a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04414] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0220b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04416] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0220c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04418] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0220d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0441a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0220e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0441c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0220f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0441e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02210] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04420] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02211] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04422] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02212] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04424] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02213] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04426] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02214] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04428] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02215] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0442a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02216] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0442c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02217] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0442e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02218] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04430] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02219] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04432] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0221a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04434] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0221b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04436] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0221c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04438] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0221d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0443a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0221e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0443c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0221f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0443e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02220] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04440] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02221] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04442] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02222] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04444] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02223] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04446] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02224] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04448] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02225] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0444a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02226] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0444c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02227] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0444e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02228] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04450] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02229] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04452] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0222a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04454] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0222b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04456] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0222c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04458] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0222d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0445a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0222e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0445c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0222f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0445e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02230] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04460] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02231] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04462] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02232] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04464] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02233] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04466] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02234] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04468] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02235] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0446a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02236] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0446c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02237] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0446e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02238] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04470] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02239] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04472] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0223a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04474] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0223b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04476] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0223c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04478] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0223d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0447a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0223e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0447c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0223f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0447e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02240] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04480] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02241] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04482] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02242] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04484] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02243] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04486] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02244] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04488] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02245] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0448a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02246] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0448c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02247] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0448e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02248] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04490] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02249] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04492] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0224a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04494] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0224b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04496] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0224c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04498] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0224d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0449a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0224e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0449c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0224f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0449e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02250] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02251] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02252] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02253] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02254] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02255] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02256] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02257] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02258] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02259] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0225a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0225b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0225c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0225d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0225e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0225f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02260] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02261] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02262] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02263] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02264] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02265] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02266] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02267] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02268] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02269] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0226a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0226b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0226c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0226d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0226e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0226f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02270] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02271] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02272] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02273] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02274] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02275] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02276] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02277] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02278] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02279] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0227a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0227b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0227c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0227d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0227e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0227f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h044fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02280] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04500] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02281] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04502] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02282] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04504] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02283] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04506] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02284] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04508] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02285] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0450a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02286] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0450c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02287] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0450e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02288] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04510] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02289] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04512] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0228a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04514] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0228b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04516] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0228c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04518] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0228d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0451a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0228e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0451c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0228f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0451e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02290] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04520] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02291] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04522] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02292] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04524] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02293] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04526] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02294] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04528] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02295] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0452a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02296] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0452c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02297] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0452e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02298] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04530] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02299] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04532] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0229a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04534] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0229b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04536] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0229c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04538] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0229d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0453a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0229e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0453c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0229f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0453e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04540] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04542] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04544] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04546] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04548] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0454a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0454c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0454e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04550] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04552] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04554] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04556] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04558] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0455a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0455c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0455e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04560] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04562] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04564] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04566] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04568] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0456a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0456c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0456e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04570] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04572] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04574] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04576] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04578] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0457a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0457c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0457e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04580] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04582] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04584] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04586] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04588] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0458a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0458c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0458e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04590] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04592] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04594] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04596] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04598] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0459a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0459c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0459e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h045fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02300] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04600] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02301] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04602] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02302] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04604] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02303] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04606] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02304] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04608] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02305] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0460a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02306] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0460c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02307] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0460e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02308] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04610] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02309] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04612] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0230a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04614] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0230b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04616] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0230c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04618] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0230d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0461a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0230e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0461c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0230f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0461e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02310] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04620] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02311] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04622] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02312] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04624] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02313] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04626] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02314] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04628] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02315] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0462a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02316] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0462c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02317] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0462e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02318] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04630] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02319] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04632] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0231a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04634] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0231b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04636] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0231c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04638] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0231d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0463a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0231e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0463c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0231f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0463e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02320] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04640] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02321] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04642] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02322] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04644] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02323] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04646] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02324] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04648] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02325] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0464a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02326] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0464c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02327] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0464e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02328] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04650] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02329] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04652] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0232a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04654] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0232b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04656] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0232c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04658] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0232d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0465a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0232e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0465c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0232f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0465e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02330] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04660] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02331] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04662] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02332] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04664] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02333] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04666] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02334] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04668] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02335] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0466a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02336] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0466c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02337] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0466e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02338] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04670] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02339] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04672] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0233a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04674] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0233b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04676] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0233c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04678] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0233d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0467a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0233e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0467c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0233f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0467e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02340] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04680] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02341] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04682] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02342] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04684] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02343] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04686] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02344] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04688] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02345] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0468a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02346] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0468c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02347] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0468e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02348] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04690] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02349] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04692] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0234a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04694] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0234b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04696] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0234c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04698] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0234d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0469a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0234e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0469c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0234f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0469e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02350] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02351] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02352] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02353] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02354] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02355] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02356] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02357] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02358] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02359] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0235a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0235b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0235c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0235d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0235e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0235f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02360] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02361] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02362] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02363] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02364] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02365] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02366] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02367] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02368] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02369] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0236a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0236b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0236c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0236d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0236e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0236f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02370] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02371] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02372] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02373] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02374] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02375] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02376] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02377] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02378] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02379] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0237a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0237b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0237c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0237d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0237e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0237f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h046fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02380] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04700] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02381] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04702] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02382] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04704] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02383] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04706] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02384] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04708] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02385] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0470a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02386] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0470c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02387] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0470e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02388] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04710] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02389] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04712] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0238a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04714] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0238b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04716] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0238c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04718] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0238d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0471a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0238e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0471c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0238f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0471e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02390] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04720] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02391] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04722] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02392] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04724] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02393] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04726] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02394] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04728] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02395] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0472a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02396] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0472c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02397] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0472e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02398] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04730] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02399] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04732] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0239a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04734] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0239b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04736] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0239c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04738] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0239d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0473a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0239e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0473c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0239f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0473e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04740] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04742] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04744] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04746] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04748] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0474a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0474c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0474e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04750] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04752] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04754] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04756] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04758] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0475a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0475c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0475e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04760] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04762] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04764] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04766] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04768] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0476a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0476c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0476e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04770] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04772] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04774] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04776] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04778] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0477a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0477c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0477e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04780] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04782] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04784] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04786] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04788] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0478a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0478c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0478e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04790] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04792] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04794] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04796] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04798] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0479a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0479c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0479e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h047fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02400] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04800] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02401] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04802] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02402] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04804] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02403] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04806] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02404] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04808] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02405] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0480a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02406] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0480c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02407] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0480e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02408] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04810] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02409] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04812] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0240a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04814] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0240b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04816] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0240c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04818] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0240d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0481a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0240e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0481c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0240f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0481e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02410] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04820] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02411] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04822] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02412] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04824] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02413] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04826] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02414] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04828] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02415] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0482a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02416] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0482c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02417] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0482e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02418] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04830] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02419] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04832] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0241a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04834] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0241b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04836] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0241c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04838] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0241d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0483a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0241e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0483c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0241f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0483e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02420] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04840] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02421] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04842] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02422] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04844] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02423] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04846] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02424] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04848] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02425] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0484a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02426] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0484c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02427] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0484e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02428] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04850] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02429] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04852] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0242a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04854] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0242b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04856] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0242c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04858] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0242d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0485a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0242e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0485c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0242f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0485e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02430] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04860] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02431] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04862] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02432] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04864] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02433] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04866] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02434] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04868] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02435] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0486a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02436] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0486c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02437] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0486e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02438] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04870] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02439] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04872] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0243a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04874] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0243b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04876] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0243c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04878] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0243d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0487a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0243e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0487c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0243f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0487e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02440] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04880] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02441] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04882] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02442] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04884] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02443] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04886] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02444] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04888] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02445] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0488a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02446] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0488c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02447] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0488e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02448] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04890] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02449] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04892] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0244a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04894] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0244b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04896] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0244c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04898] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0244d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0489a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0244e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0489c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0244f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0489e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02450] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02451] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02452] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02453] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02454] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02455] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02456] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02457] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02458] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02459] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0245a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0245b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0245c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0245d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0245e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0245f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02460] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02461] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02462] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02463] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02464] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02465] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02466] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02467] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02468] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02469] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0246a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0246b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0246c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0246d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0246e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0246f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02470] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02471] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02472] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02473] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02474] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02475] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02476] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02477] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02478] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02479] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0247a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0247b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0247c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0247d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0247e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0247f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h048fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02480] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04900] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02481] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04902] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02482] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04904] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02483] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04906] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02484] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04908] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02485] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0490a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02486] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0490c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02487] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0490e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02488] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04910] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02489] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04912] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0248a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04914] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0248b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04916] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0248c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04918] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0248d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0491a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0248e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0491c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0248f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0491e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02490] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04920] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02491] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04922] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02492] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04924] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02493] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04926] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02494] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04928] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02495] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0492a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02496] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0492c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02497] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0492e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02498] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04930] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02499] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04932] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0249a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04934] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0249b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04936] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0249c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04938] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0249d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0493a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0249e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0493c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0249f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0493e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04940] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04942] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04944] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04946] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04948] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0494a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0494c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0494e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04950] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04952] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04954] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04956] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04958] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0495a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0495c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0495e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04960] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04962] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04964] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04966] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04968] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0496a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0496c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0496e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04970] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04972] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04974] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04976] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04978] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0497a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0497c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0497e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04980] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04982] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04984] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04986] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04988] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0498a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0498c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0498e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04990] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04992] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04994] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04996] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04998] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0499a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0499c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0499e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h049fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02500] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02501] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02502] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02503] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02504] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02505] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02506] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02507] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02508] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02509] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0250a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0250b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0250c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0250d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0250e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0250f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02510] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02511] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02512] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02513] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02514] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02515] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02516] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02517] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02518] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02519] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0251a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0251b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0251c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0251d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0251e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0251f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02520] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02521] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02522] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02523] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02524] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02525] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02526] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02527] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02528] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02529] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0252a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0252b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0252c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0252d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0252e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0252f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02530] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02531] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02532] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02533] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02534] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02535] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02536] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02537] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02538] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02539] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0253a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0253b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0253c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0253d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0253e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0253f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02540] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02541] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02542] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02543] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02544] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02545] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02546] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02547] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02548] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02549] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0254a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0254b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0254c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0254d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0254e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0254f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04a9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02550] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02551] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02552] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02553] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02554] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02555] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02556] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02557] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02558] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ab0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02559] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ab2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0255a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ab4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0255b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ab6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0255c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ab8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0255d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0255e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04abc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0255f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04abe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02560] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ac0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02561] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ac2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02562] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ac4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02563] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ac6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02564] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ac8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02565] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02566] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04acc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02567] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ace] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02568] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ad0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02569] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ad2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0256a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ad4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0256b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ad6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0256c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ad8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0256d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ada] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0256e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04adc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0256f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ade] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02570] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ae0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02571] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ae2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02572] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ae4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02573] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ae6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02574] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ae8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02575] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02576] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02577] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04aee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02578] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04af0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02579] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04af2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0257a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04af4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0257b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04af6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0257c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04af8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0257d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04afa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0257e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04afc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0257f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04afe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02580] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02581] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02582] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02583] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02584] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02585] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02586] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02587] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02588] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02589] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0258a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0258b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0258c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0258d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0258e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0258f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02590] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02591] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02592] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02593] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02594] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02595] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02596] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02597] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02598] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02599] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0259a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0259b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0259c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0259d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0259e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0259f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04b9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ba0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ba2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ba4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ba6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ba8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04baa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04be0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04be2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04be4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04be6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04be8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04bfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02600] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02601] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02602] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02603] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02604] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02605] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02606] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02607] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02608] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02609] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0260a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0260b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0260c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0260d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0260e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0260f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02610] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02611] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02612] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02613] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02614] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02615] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02616] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02617] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02618] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02619] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0261a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0261b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0261c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0261d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0261e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0261f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02620] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02621] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02622] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02623] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02624] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02625] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02626] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02627] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02628] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02629] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0262a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0262b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0262c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0262d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0262e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0262f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02630] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02631] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02632] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02633] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02634] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02635] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02636] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02637] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02638] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02639] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0263a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0263b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0263c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0263d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0263e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0263f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02640] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02641] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02642] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02643] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02644] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02645] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02646] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02647] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02648] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02649] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0264a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0264b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0264c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0264d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0264e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0264f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04c9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02650] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ca0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02651] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ca2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02652] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ca4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02653] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ca6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02654] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ca8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02655] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04caa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02656] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02657] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02658] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02659] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0265a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0265b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0265c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0265d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0265e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0265f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02660] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02661] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02662] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02663] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02664] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02665] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02666] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ccc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02667] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02668] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02669] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0266a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0266b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0266c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0266d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0266e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0266f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02670] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ce0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02671] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ce2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02672] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ce4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02673] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ce6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02674] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ce8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02675] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02676] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02677] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02678] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02679] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0267a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0267b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0267c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0267d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0267e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0267f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04cfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02680] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02681] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02682] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02683] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02684] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02685] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02686] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02687] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02688] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02689] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0268a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0268b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0268c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0268d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0268e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0268f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02690] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02691] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02692] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02693] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02694] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02695] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02696] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02697] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02698] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02699] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0269a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0269b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0269c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0269d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0269e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0269f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04d9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04da0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04da2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04da4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04da6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04da8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04daa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04db0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04db2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04db4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04db6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04db8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ddc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04de0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04de2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04de4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04de6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04de8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04df0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04df2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04df4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04df6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04df8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04dfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02700] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02701] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02702] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02703] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02704] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02705] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02706] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02707] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02708] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02709] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0270a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0270b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0270c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0270d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0270e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0270f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02710] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02711] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02712] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02713] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02714] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02715] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02716] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02717] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02718] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02719] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0271a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0271b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0271c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0271d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0271e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0271f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02720] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02721] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02722] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02723] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02724] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02725] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02726] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02727] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02728] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02729] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0272a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0272b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0272c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0272d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0272e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0272f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02730] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02731] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02732] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02733] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02734] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02735] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02736] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02737] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02738] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02739] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0273a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0273b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0273c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0273d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0273e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0273f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02740] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02741] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02742] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02743] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02744] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02745] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02746] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02747] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02748] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02749] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0274a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0274b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0274c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0274d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0274e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0274f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04e9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02750] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ea0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02751] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ea2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02752] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ea4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02753] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ea6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02754] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ea8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02755] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02756] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02757] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02758] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02759] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0275a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0275b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0275c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0275d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0275e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ebc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0275f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ebe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02760] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ec0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02761] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ec2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02762] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ec4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02763] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ec6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02764] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ec8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02765] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02766] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ecc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02767] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ece] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02768] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ed0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02769] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ed2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0276a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ed4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0276b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ed6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0276c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ed8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0276d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0276e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04edc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0276f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ede] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02770] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ee0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02771] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ee2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02772] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ee4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02773] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ee6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02774] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ee8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02775] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02776] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02777] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04eee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02778] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ef0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02779] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ef2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0277a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ef4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0277b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ef6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0277c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ef8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0277d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04efa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0277e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04efc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0277f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04efe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02780] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02781] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02782] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02783] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02784] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02785] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02786] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02787] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02788] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02789] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0278a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0278b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0278c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0278d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0278e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0278f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02790] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02791] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02792] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02793] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02794] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02795] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02796] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02797] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02798] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02799] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0279a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0279b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0279c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0279d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0279e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0279f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04f9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04faa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fe0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fe2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fe4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fe6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fe8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04fee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ff0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ff2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ff4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ff6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ff8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ffa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ffc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h04ffe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02800] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05000] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02801] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05002] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02802] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05004] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02803] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05006] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02804] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05008] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02805] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0500a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02806] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0500c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02807] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0500e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02808] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05010] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02809] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05012] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0280a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05014] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0280b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05016] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0280c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05018] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0280d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0501a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0280e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0501c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0280f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0501e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02810] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05020] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02811] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05022] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02812] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05024] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02813] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05026] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02814] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05028] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02815] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0502a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02816] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0502c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02817] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0502e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02818] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05030] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02819] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05032] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0281a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05034] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0281b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05036] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0281c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05038] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0281d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0503a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0281e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0503c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0281f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0503e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02820] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05040] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02821] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05042] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02822] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05044] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02823] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05046] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02824] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05048] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02825] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0504a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02826] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0504c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02827] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0504e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02828] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05050] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02829] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05052] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0282a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05054] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0282b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05056] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0282c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05058] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0282d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0505a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0282e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0505c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0282f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0505e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02830] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05060] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02831] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05062] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02832] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05064] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02833] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05066] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02834] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05068] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02835] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0506a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02836] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0506c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02837] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0506e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02838] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05070] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02839] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05072] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0283a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05074] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0283b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05076] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0283c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05078] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0283d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0507a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0283e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0507c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0283f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0507e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02840] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05080] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02841] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05082] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02842] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05084] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02843] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05086] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02844] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05088] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02845] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0508a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02846] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0508c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02847] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0508e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02848] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05090] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02849] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05092] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0284a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05094] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0284b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05096] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0284c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05098] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0284d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0509a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0284e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0509c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0284f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0509e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02850] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02851] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02852] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02853] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02854] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02855] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02856] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02857] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02858] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02859] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0285a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0285b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0285c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0285d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0285e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0285f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02860] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02861] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02862] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02863] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02864] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02865] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02866] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02867] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02868] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02869] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0286a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0286b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0286c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0286d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0286e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0286f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02870] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02871] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02872] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02873] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02874] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02875] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02876] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02877] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02878] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02879] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0287a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0287b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0287c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0287d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0287e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0287f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h050fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02880] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05100] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02881] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05102] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02882] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05104] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02883] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05106] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02884] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05108] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02885] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0510a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02886] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0510c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02887] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0510e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02888] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05110] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02889] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05112] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0288a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05114] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0288b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05116] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0288c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05118] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0288d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0511a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0288e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0511c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0288f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0511e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02890] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05120] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02891] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05122] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02892] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05124] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02893] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05126] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02894] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05128] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02895] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0512a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02896] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0512c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02897] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0512e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02898] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05130] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02899] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05132] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0289a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05134] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0289b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05136] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0289c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05138] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0289d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0513a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0289e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0513c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0289f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0513e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05140] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05142] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05144] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05146] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05148] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0514a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0514c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0514e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05150] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05152] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05154] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05156] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05158] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0515a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0515c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0515e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05160] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05162] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05164] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05166] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05168] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0516a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0516c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0516e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05170] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05172] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05174] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05176] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05178] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0517a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0517c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0517e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05180] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05182] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05184] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05186] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05188] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0518a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0518c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0518e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05190] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05192] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05194] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05196] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05198] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0519a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0519c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0519e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h051fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02900] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05200] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02901] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05202] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02902] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05204] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02903] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05206] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02904] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05208] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02905] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0520a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02906] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0520c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02907] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0520e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02908] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05210] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02909] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05212] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0290a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05214] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0290b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05216] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0290c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05218] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0290d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0521a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0290e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0521c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0290f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0521e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02910] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05220] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02911] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05222] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02912] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05224] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02913] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05226] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02914] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05228] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02915] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0522a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02916] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0522c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02917] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0522e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02918] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05230] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02919] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05232] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0291a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05234] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0291b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05236] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0291c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05238] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0291d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0523a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0291e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0523c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0291f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0523e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02920] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05240] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02921] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05242] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02922] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05244] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02923] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05246] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02924] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05248] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02925] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0524a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02926] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0524c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02927] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0524e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02928] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05250] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02929] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05252] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0292a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05254] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0292b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05256] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0292c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05258] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0292d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0525a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0292e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0525c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0292f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0525e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02930] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05260] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02931] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05262] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02932] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05264] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02933] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05266] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02934] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05268] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02935] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0526a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02936] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0526c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02937] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0526e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02938] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05270] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02939] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05272] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0293a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05274] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0293b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05276] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0293c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05278] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0293d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0527a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0293e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0527c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0293f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0527e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02940] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05280] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02941] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05282] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02942] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05284] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02943] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05286] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02944] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05288] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02945] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0528a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02946] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0528c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02947] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0528e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02948] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05290] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02949] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05292] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0294a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05294] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0294b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05296] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0294c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05298] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0294d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0529a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0294e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0529c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0294f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0529e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02950] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02951] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02952] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02953] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02954] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02955] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02956] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02957] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02958] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02959] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0295a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0295b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0295c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0295d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0295e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0295f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02960] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02961] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02962] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02963] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02964] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02965] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02966] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02967] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02968] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02969] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0296a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0296b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0296c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0296d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0296e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0296f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02970] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02971] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02972] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02973] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02974] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02975] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02976] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02977] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02978] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02979] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0297a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0297b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0297c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0297d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0297e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0297f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h052fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02980] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05300] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02981] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05302] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02982] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05304] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02983] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05306] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02984] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05308] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02985] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0530a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02986] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0530c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02987] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0530e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02988] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05310] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02989] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05312] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0298a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05314] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0298b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05316] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0298c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05318] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0298d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0531a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0298e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0531c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0298f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0531e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02990] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05320] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02991] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05322] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02992] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05324] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02993] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05326] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02994] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05328] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02995] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0532a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02996] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0532c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02997] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0532e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02998] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05330] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02999] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05332] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0299a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05334] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0299b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05336] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0299c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05338] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0299d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0533a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0299e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0533c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0299f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0533e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05340] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05342] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05344] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05346] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05348] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0534a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0534c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0534e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05350] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05352] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05354] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05356] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05358] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0535a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0535c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0535e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05360] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05362] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05364] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05366] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05368] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0536a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0536c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0536e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05370] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05372] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05374] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05376] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05378] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0537a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0537c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0537e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05380] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05382] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05384] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05386] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05388] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0538a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0538c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0538e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05390] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05392] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05394] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05396] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05398] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0539a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0539c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0539e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h053fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05400] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05402] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05404] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05406] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05408] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0540a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0540c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0540e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05410] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05412] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05414] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05416] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05418] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0541a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0541c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0541e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05420] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05422] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05424] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05426] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05428] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0542a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0542c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0542e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05430] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05432] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05434] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05436] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05438] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0543a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0543c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0543e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05440] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05442] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05444] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05446] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05448] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0544a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0544c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0544e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05450] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05452] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05454] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05456] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05458] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0545a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0545c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0545e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05460] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05462] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05464] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05466] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05468] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0546a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0546c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0546e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05470] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05472] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05474] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05476] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05478] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0547a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0547c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0547e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05480] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05482] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05484] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05486] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05488] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0548a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0548c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0548e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05490] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05492] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05494] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05496] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05498] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0549a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0549c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0549e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h054fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05500] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05502] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05504] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05506] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05508] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0550a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0550c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0550e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05510] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05512] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05514] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05516] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05518] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0551a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0551c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0551e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05520] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05522] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05524] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05526] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05528] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0552a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0552c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0552e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05530] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05532] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05534] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05536] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05538] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0553a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0553c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0553e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05540] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05542] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05544] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05546] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05548] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0554a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0554c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0554e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05550] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05552] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aaa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05554] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05556] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05558] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0555a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0555c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aaf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0555e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05560] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05562] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05564] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05566] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05568] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0556a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0556c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0556e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05570] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05572] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05574] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02abb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05576] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02abc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05578] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02abd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0557a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02abe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0557c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02abf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0557e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05580] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05582] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05584] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05586] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05588] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0558a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0558c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0558e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05590] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05592] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05594] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02acb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05596] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02acc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05598] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02acd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0559a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ace] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0559c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02acf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0559e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ada] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02adb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02adc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02add] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ade] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02adf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aeb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02afa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02afb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02afc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02afd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02afe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h055fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05600] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05602] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05604] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05606] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05608] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0560a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0560c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0560e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05610] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05612] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05614] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05616] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05618] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0561a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0561c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0561e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05620] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05622] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05624] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05626] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05628] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0562a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0562c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0562e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05630] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05632] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05634] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05636] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05638] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0563a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0563c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0563e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05640] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05642] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05644] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05646] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05648] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0564a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0564c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0564e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05650] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05652] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05654] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05656] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05658] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0565a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0565c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0565e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05660] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05662] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05664] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05666] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05668] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0566a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0566c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0566e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05670] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05672] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05674] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05676] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05678] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0567a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0567c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0567e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05680] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05682] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05684] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05686] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05688] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0568a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0568c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0568e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05690] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05692] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05694] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05696] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05698] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0569a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0569c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0569e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h056fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05700] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05702] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05704] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05706] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05708] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0570a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0570c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0570e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05710] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05712] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05714] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05716] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05718] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0571a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0571c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0571e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05720] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05722] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05724] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05726] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05728] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0572a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0572c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0572e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05730] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05732] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05734] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05736] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05738] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0573a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0573c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0573e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05740] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05742] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05744] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05746] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05748] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0574a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0574c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0574e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05750] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05752] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02baa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05754] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05756] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05758] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0575a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0575c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02baf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0575e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05760] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05762] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05764] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05766] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05768] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0576a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0576c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0576e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05770] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05772] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05774] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05776] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05778] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0577a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0577c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0577e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05780] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05782] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05784] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05786] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05788] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0578a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0578c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0578e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05790] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05792] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05794] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05796] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05798] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0579a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0579c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0579e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02beb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h057fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05800] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05802] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05804] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05806] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05808] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0580a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0580c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0580e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05810] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05812] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05814] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05816] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05818] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0581a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0581c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0581e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05820] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05822] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05824] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05826] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05828] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0582a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0582c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0582e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05830] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05832] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05834] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05836] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05838] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0583a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0583c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0583e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05840] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05842] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05844] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05846] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05848] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0584a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0584c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0584e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05850] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05852] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05854] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05856] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05858] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0585a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0585c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0585e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05860] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05862] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05864] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05866] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05868] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0586a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0586c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0586e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05870] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05872] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05874] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05876] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05878] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0587a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0587c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0587e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05880] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05882] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05884] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05886] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05888] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0588a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0588c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0588e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05890] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05892] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05894] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05896] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05898] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0589a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0589c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0589e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h058fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05900] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05902] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05904] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05906] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05908] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0590a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0590c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0590e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05910] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05912] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05914] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05916] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05918] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0591a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0591c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0591e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05920] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05922] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05924] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05926] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05928] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0592a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0592c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0592e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05930] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05932] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05934] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05936] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05938] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0593a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0593c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0593e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05940] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05942] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05944] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05946] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05948] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0594a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0594c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0594e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05950] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05952] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02caa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05954] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05956] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05958] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0595a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0595c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02caf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0595e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05960] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05962] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05964] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05966] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05968] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0596a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0596c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0596e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05970] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05972] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05974] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05976] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05978] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0597a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0597c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0597e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05980] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05982] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05984] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05986] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05988] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0598a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0598c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0598e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05990] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05992] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05994] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ccb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05996] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ccc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05998] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ccd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0599a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0599c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ccf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0599e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ceb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ced] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h059fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05a9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ab0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ab2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ab4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ab6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ab8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05abc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05abe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ac0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ac2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ac4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ac6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ac8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05acc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ace] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ad0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ad2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ad4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ad6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ad8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ada] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05adc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ade] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ae0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ae2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ae4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ae6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ae8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05aee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05af0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05af2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05af4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05af6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05af8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05afa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05afc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05afe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02daa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02daf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05b9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ba0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ba2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ba4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ba6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ba8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05baa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ddb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ddc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ddd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ddf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02deb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ded] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02def] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05be0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05be2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05be4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05be6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05be8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05bfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05c9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ca0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ca2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ca4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ca6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ca8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05caa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ccc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ce0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ce2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ce4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ce6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ce8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05cfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eaa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ead] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eaf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ebb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ebc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ebd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ebe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ebf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ecb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ecc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ecd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ece] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ecf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05d9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05da0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05da2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05da4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05da6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05da8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05daa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05db0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05db2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05db4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02edb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05db6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02edc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05db8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02edd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ede] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02edf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eeb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ddc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05de0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05de2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05de4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05de6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05de8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05df0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05df2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02efa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05df4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02efb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05df6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02efc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05df8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02efd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02efe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05dfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05e9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ea0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ea2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ea4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ea6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ea8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ebc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ebe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ec0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ec2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ec4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ec6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ec8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ecc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ece] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ed0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ed2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ed4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ed6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ed8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05edc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ede] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ee0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ee2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ee4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ee6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ee8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05eee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ef0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ef2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ef4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ef6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ef8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05efa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05efc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05efe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02faa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02faf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05f9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05faa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02feb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fe0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fe2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fe4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fe6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fe8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05fee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ff0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ff2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ffa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ff4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ffb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ff6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ffc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ff8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ffd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ffa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ffe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ffc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h05ffe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03000] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06000] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03001] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06002] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03002] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06004] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03003] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06006] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03004] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06008] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03005] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0600a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03006] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0600c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03007] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0600e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03008] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06010] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03009] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06012] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0300a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06014] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0300b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06016] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0300c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06018] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0300d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0601a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0300e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0601c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0300f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0601e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03010] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06020] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03011] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06022] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03012] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06024] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03013] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06026] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03014] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06028] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03015] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0602a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03016] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0602c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03017] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0602e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03018] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06030] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03019] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06032] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0301a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06034] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0301b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06036] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0301c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06038] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0301d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0603a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0301e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0603c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0301f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0603e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03020] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06040] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03021] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06042] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03022] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06044] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03023] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06046] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03024] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06048] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03025] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0604a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03026] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0604c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03027] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0604e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03028] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06050] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03029] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06052] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0302a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06054] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0302b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06056] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0302c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06058] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0302d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0605a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0302e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0605c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0302f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0605e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03030] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06060] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03031] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06062] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03032] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06064] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03033] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06066] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03034] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06068] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03035] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0606a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03036] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0606c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03037] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0606e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03038] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06070] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03039] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06072] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0303a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06074] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0303b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06076] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0303c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06078] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0303d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0607a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0303e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0607c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0303f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0607e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03040] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06080] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03041] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06082] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03042] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06084] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03043] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06086] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03044] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06088] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03045] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0608a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03046] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0608c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03047] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0608e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03048] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06090] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03049] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06092] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0304a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06094] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0304b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06096] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0304c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06098] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0304d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0609a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0304e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0609c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0304f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0609e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03050] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03051] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03052] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03053] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03054] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03055] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03056] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03057] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03058] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03059] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0305a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0305b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0305c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0305d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0305e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0305f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03060] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03061] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03062] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03063] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03064] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03065] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03066] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03067] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03068] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03069] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0306a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0306b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0306c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0306d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0306e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0306f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03070] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03071] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03072] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03073] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03074] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03075] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03076] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03077] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03078] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03079] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0307a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0307b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0307c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0307d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0307e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0307f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h060fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03080] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06100] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03081] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06102] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03082] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06104] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03083] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06106] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03084] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06108] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03085] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0610a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03086] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0610c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03087] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0610e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03088] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06110] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03089] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06112] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0308a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06114] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0308b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06116] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0308c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06118] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0308d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0611a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0308e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0611c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0308f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0611e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03090] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06120] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03091] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06122] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03092] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06124] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03093] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06126] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03094] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06128] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03095] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0612a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03096] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0612c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03097] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0612e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03098] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06130] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03099] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06132] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0309a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06134] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0309b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06136] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0309c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06138] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0309d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0613a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0309e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0613c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0309f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0613e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06140] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06142] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06144] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06146] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06148] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0614a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0614c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0614e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06150] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06152] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06154] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06156] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06158] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0615a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0615c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0615e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06160] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06162] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06164] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06166] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06168] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0616a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0616c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0616e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06170] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06172] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06174] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06176] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06178] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0617a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0617c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0617e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06180] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06182] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06184] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06186] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06188] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0618a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0618c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0618e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06190] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06192] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06194] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06196] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06198] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0619a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0619c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0619e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h061fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03100] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06200] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03101] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06202] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03102] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06204] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03103] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06206] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03104] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06208] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03105] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0620a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03106] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0620c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03107] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0620e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03108] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06210] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03109] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06212] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0310a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06214] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0310b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06216] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0310c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06218] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0310d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0621a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0310e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0621c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0310f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0621e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03110] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06220] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03111] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06222] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03112] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06224] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03113] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06226] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03114] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06228] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03115] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0622a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03116] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0622c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03117] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0622e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03118] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06230] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03119] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06232] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0311a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06234] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0311b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06236] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0311c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06238] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0311d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0623a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0311e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0623c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0311f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0623e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03120] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06240] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03121] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06242] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03122] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06244] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03123] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06246] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03124] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06248] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03125] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0624a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03126] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0624c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03127] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0624e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03128] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06250] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03129] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06252] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0312a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06254] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0312b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06256] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0312c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06258] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0312d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0625a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0312e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0625c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0312f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0625e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03130] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06260] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03131] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06262] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03132] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06264] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03133] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06266] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03134] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06268] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03135] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0626a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03136] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0626c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03137] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0626e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03138] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06270] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03139] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06272] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0313a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06274] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0313b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06276] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0313c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06278] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0313d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0627a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0313e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0627c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0313f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0627e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03140] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06280] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03141] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06282] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03142] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06284] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03143] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06286] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03144] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06288] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03145] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0628a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03146] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0628c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03147] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0628e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03148] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06290] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03149] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06292] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0314a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06294] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0314b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06296] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0314c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06298] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0314d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0629a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0314e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0629c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0314f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0629e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03150] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03151] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03152] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03153] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03154] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03155] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03156] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03157] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03158] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03159] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0315a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0315b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0315c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0315d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0315e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0315f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03160] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03161] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03162] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03163] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03164] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03165] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03166] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03167] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03168] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03169] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0316a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0316b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0316c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0316d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0316e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0316f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03170] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03171] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03172] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03173] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03174] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03175] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03176] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03177] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03178] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03179] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0317a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0317b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0317c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0317d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0317e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0317f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h062fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03180] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06300] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03181] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06302] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03182] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06304] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03183] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06306] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03184] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06308] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03185] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0630a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03186] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0630c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03187] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0630e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03188] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06310] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03189] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06312] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0318a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06314] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0318b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06316] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0318c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06318] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0318d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0631a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0318e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0631c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0318f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0631e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03190] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06320] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03191] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06322] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03192] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06324] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03193] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06326] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03194] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06328] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03195] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0632a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03196] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0632c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03197] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0632e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03198] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06330] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03199] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06332] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0319a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06334] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0319b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06336] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0319c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06338] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0319d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0633a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0319e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0633c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0319f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0633e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06340] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06342] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06344] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06346] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06348] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0634a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0634c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0634e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06350] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06352] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06354] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06356] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06358] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0635a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0635c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0635e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06360] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06362] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06364] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06366] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06368] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0636a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0636c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0636e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06370] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06372] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06374] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06376] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06378] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0637a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0637c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0637e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06380] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06382] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06384] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06386] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06388] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0638a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0638c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0638e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06390] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06392] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06394] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06396] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06398] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0639a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0639c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0639e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h063fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03200] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06400] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03201] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06402] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03202] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06404] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03203] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06406] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03204] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06408] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03205] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0640a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03206] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0640c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03207] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0640e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03208] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06410] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03209] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06412] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0320a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06414] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0320b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06416] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0320c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06418] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0320d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0641a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0320e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0641c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0320f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0641e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03210] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06420] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03211] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06422] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03212] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06424] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03213] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06426] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03214] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06428] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03215] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0642a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03216] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0642c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03217] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0642e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03218] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06430] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03219] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06432] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0321a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06434] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0321b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06436] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0321c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06438] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0321d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0643a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0321e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0643c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0321f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0643e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03220] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06440] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03221] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06442] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03222] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06444] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03223] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06446] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03224] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06448] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03225] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0644a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03226] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0644c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03227] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0644e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03228] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06450] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03229] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06452] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0322a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06454] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0322b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06456] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0322c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06458] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0322d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0645a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0322e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0645c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0322f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0645e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03230] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06460] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03231] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06462] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03232] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06464] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03233] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06466] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03234] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06468] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03235] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0646a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03236] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0646c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03237] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0646e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03238] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06470] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03239] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06472] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0323a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06474] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0323b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06476] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0323c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06478] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0323d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0647a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0323e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0647c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0323f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0647e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03240] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06480] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03241] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06482] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03242] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06484] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03243] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06486] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03244] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06488] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03245] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0648a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03246] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0648c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03247] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0648e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03248] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06490] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03249] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06492] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0324a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06494] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0324b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06496] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0324c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06498] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0324d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0649a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0324e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0649c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0324f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0649e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03250] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03251] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03252] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03253] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03254] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03255] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03256] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03257] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03258] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03259] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0325a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0325b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0325c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0325d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0325e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0325f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03260] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03261] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03262] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03263] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03264] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03265] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03266] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03267] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03268] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03269] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0326a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0326b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0326c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0326d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0326e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0326f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03270] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03271] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03272] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03273] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03274] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03275] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03276] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03277] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03278] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03279] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0327a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0327b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0327c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0327d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0327e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0327f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h064fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03280] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06500] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03281] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06502] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03282] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06504] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03283] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06506] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03284] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06508] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03285] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0650a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03286] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0650c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03287] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0650e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03288] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06510] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03289] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06512] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0328a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06514] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0328b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06516] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0328c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06518] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0328d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0651a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0328e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0651c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0328f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0651e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03290] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06520] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03291] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06522] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03292] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06524] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03293] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06526] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03294] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06528] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03295] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0652a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03296] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0652c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03297] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0652e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03298] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06530] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03299] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06532] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0329a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06534] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0329b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06536] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0329c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06538] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0329d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0653a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0329e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0653c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0329f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0653e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06540] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06542] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06544] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06546] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06548] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0654a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0654c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0654e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06550] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06552] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06554] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06556] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06558] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0655a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0655c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0655e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06560] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06562] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06564] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06566] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06568] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0656a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0656c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0656e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06570] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06572] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06574] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06576] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06578] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0657a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0657c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0657e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06580] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06582] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06584] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06586] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06588] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0658a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0658c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0658e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06590] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06592] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06594] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06596] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06598] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0659a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0659c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0659e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h065fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03300] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06600] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03301] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06602] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03302] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06604] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03303] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06606] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03304] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06608] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03305] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0660a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03306] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0660c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03307] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0660e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03308] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06610] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03309] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06612] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0330a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06614] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0330b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06616] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0330c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06618] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0330d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0661a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0330e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0661c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0330f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0661e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03310] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06620] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03311] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06622] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03312] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06624] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03313] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06626] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03314] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06628] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03315] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0662a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03316] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0662c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03317] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0662e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03318] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06630] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03319] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06632] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0331a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06634] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0331b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06636] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0331c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06638] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0331d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0663a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0331e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0663c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0331f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0663e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03320] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06640] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03321] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06642] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03322] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06644] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03323] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06646] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03324] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06648] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03325] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0664a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03326] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0664c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03327] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0664e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03328] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06650] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03329] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06652] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0332a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06654] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0332b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06656] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0332c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06658] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0332d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0665a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0332e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0665c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0332f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0665e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03330] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06660] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03331] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06662] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03332] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06664] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03333] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06666] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03334] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06668] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03335] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0666a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03336] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0666c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03337] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0666e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03338] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06670] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03339] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06672] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0333a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06674] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0333b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06676] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0333c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06678] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0333d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0667a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0333e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0667c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0333f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0667e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03340] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06680] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03341] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06682] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03342] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06684] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03343] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06686] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03344] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06688] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03345] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0668a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03346] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0668c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03347] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0668e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03348] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06690] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03349] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06692] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0334a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06694] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0334b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06696] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0334c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06698] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0334d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0669a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0334e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0669c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0334f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0669e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03350] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03351] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03352] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03353] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03354] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03355] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03356] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03357] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03358] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03359] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0335a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0335b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0335c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0335d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0335e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0335f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03360] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03361] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03362] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03363] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03364] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03365] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03366] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03367] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03368] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03369] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0336a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0336b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0336c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0336d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0336e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0336f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03370] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03371] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03372] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03373] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03374] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03375] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03376] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03377] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03378] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03379] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0337a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0337b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0337c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0337d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0337e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0337f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h066fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03380] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06700] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03381] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06702] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03382] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06704] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03383] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06706] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03384] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06708] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03385] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0670a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03386] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0670c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03387] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0670e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03388] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06710] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03389] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06712] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0338a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06714] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0338b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06716] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0338c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06718] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0338d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0671a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0338e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0671c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0338f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0671e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03390] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06720] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03391] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06722] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03392] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06724] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03393] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06726] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03394] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06728] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03395] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0672a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03396] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0672c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03397] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0672e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03398] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06730] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03399] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06732] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0339a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06734] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0339b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06736] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0339c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06738] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0339d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0673a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0339e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0673c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0339f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0673e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06740] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06742] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06744] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06746] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06748] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0674a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0674c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0674e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06750] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06752] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06754] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06756] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06758] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0675a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0675c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0675e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06760] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06762] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06764] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06766] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06768] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0676a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0676c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0676e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06770] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06772] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06774] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06776] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06778] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0677a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0677c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0677e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06780] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06782] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06784] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06786] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06788] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0678a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0678c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0678e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06790] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06792] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06794] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06796] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06798] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0679a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0679c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0679e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h067fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03400] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06800] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03401] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06802] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03402] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06804] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03403] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06806] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03404] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06808] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03405] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0680a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03406] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0680c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03407] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0680e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03408] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06810] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03409] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06812] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0340a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06814] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0340b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06816] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0340c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06818] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0340d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0681a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0340e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0681c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0340f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0681e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03410] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06820] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03411] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06822] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03412] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06824] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03413] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06826] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03414] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06828] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03415] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0682a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03416] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0682c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03417] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0682e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03418] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06830] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03419] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06832] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0341a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06834] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0341b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06836] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0341c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06838] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0341d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0683a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0341e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0683c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0341f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0683e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03420] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06840] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03421] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06842] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03422] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06844] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03423] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06846] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03424] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06848] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03425] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0684a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03426] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0684c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03427] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0684e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03428] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06850] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03429] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06852] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0342a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06854] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0342b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06856] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0342c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06858] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0342d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0685a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0342e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0685c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0342f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0685e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03430] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06860] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03431] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06862] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03432] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06864] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03433] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06866] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03434] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06868] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03435] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0686a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03436] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0686c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03437] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0686e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03438] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06870] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03439] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06872] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0343a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06874] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0343b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06876] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0343c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06878] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0343d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0687a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0343e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0687c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0343f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0687e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03440] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06880] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03441] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06882] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03442] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06884] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03443] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06886] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03444] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06888] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03445] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0688a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03446] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0688c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03447] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0688e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03448] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06890] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03449] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06892] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0344a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06894] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0344b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06896] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0344c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06898] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0344d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0689a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0344e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0689c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0344f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0689e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03450] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03451] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03452] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03453] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03454] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03455] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03456] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03457] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03458] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03459] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0345a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0345b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0345c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0345d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0345e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0345f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03460] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03461] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03462] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03463] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03464] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03465] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03466] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03467] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03468] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03469] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0346a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0346b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0346c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0346d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0346e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0346f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03470] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03471] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03472] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03473] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03474] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03475] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03476] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03477] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03478] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03479] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0347a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0347b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0347c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0347d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0347e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0347f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h068fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03480] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06900] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03481] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06902] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03482] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06904] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03483] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06906] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03484] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06908] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03485] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0690a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03486] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0690c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03487] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0690e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03488] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06910] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03489] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06912] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0348a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06914] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0348b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06916] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0348c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06918] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0348d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0691a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0348e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0691c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0348f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0691e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03490] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06920] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03491] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06922] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03492] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06924] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03493] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06926] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03494] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06928] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03495] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0692a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03496] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0692c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03497] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0692e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03498] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06930] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03499] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06932] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0349a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06934] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0349b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06936] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0349c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06938] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0349d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0693a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0349e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0693c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0349f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0693e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06940] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06942] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06944] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06946] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06948] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0694a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0694c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0694e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06950] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06952] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06954] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06956] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06958] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0695a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0695c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0695e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06960] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06962] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06964] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06966] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06968] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0696a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0696c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0696e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06970] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06972] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06974] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06976] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06978] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0697a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0697c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0697e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06980] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06982] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06984] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06986] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06988] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0698a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0698c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0698e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06990] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06992] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06994] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06996] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06998] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0699a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0699c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0699e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h069fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03500] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03501] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03502] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03503] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03504] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03505] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03506] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03507] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03508] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03509] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0350a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0350b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0350c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0350d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0350e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0350f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03510] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03511] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03512] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03513] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03514] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03515] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03516] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03517] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03518] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03519] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0351a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0351b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0351c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0351d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0351e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0351f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03520] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03521] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03522] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03523] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03524] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03525] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03526] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03527] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03528] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03529] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0352a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0352b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0352c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0352d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0352e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0352f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03530] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03531] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03532] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03533] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03534] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03535] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03536] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03537] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03538] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03539] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0353a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0353b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0353c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0353d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0353e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0353f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03540] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03541] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03542] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03543] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03544] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03545] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03546] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03547] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03548] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03549] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0354a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0354b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0354c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0354d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0354e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0354f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06a9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03550] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03551] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03552] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03553] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03554] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03555] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03556] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03557] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03558] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ab0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03559] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ab2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0355a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ab4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0355b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ab6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0355c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ab8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0355d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0355e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06abc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0355f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06abe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03560] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ac0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03561] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ac2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03562] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ac4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03563] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ac6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03564] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ac8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03565] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03566] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06acc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03567] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ace] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03568] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ad0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03569] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ad2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0356a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ad4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0356b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ad6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0356c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ad8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0356d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ada] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0356e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06adc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0356f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ade] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03570] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ae0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03571] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ae2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03572] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ae4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03573] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ae6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03574] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ae8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03575] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03576] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03577] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06aee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03578] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06af0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03579] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06af2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0357a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06af4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0357b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06af6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0357c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06af8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0357d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06afa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0357e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06afc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0357f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06afe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03580] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03581] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03582] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03583] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03584] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03585] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03586] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03587] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03588] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03589] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0358a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0358b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0358c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0358d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0358e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0358f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03590] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03591] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03592] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03593] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03594] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03595] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03596] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03597] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03598] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03599] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0359a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0359b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0359c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0359d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0359e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0359f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06b9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ba0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ba2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ba4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ba6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ba8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06baa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06be0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06be2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06be4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06be6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06be8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06bfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03600] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03601] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03602] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03603] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03604] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03605] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03606] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03607] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03608] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03609] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0360a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0360b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0360c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0360d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0360e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0360f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03610] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03611] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03612] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03613] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03614] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03615] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03616] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03617] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03618] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03619] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0361a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0361b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0361c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0361d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0361e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0361f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03620] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03621] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03622] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03623] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03624] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03625] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03626] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03627] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03628] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03629] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0362a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0362b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0362c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0362d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0362e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0362f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03630] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03631] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03632] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03633] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03634] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03635] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03636] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03637] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03638] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03639] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0363a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0363b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0363c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0363d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0363e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0363f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03640] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03641] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03642] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03643] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03644] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03645] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03646] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03647] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03648] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03649] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0364a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0364b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0364c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0364d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0364e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0364f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06c9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03650] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ca0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03651] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ca2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03652] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ca4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03653] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ca6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03654] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ca8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03655] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06caa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03656] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03657] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03658] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03659] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0365a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0365b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0365c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0365d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0365e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0365f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03660] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03661] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03662] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03663] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03664] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03665] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03666] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ccc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03667] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03668] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03669] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0366a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0366b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0366c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0366d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0366e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0366f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03670] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ce0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03671] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ce2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03672] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ce4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03673] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ce6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03674] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ce8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03675] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03676] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03677] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03678] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03679] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0367a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0367b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0367c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0367d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0367e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0367f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06cfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03680] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03681] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03682] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03683] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03684] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03685] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03686] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03687] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03688] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03689] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0368a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0368b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0368c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0368d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0368e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0368f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03690] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03691] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03692] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03693] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03694] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03695] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03696] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03697] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03698] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03699] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0369a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0369b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0369c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0369d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0369e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0369f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06d9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06da0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06da2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06da4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06da6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06da8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06daa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06db0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06db2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06db4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06db6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06db8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ddc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06de0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06de2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06de4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06de6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06de8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06df0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06df2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06df4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06df6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06df8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06dfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03700] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03701] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03702] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03703] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03704] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03705] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03706] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03707] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03708] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03709] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0370a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0370b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0370c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0370d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0370e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0370f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03710] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03711] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03712] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03713] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03714] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03715] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03716] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03717] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03718] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03719] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0371a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0371b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0371c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0371d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0371e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0371f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03720] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03721] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03722] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03723] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03724] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03725] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03726] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03727] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03728] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03729] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0372a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0372b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0372c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0372d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0372e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0372f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03730] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03731] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03732] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03733] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03734] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03735] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03736] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03737] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03738] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03739] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0373a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0373b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0373c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0373d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0373e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0373f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03740] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03741] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03742] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03743] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03744] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03745] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03746] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03747] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03748] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03749] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0374a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0374b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0374c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0374d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0374e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0374f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06e9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03750] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ea0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03751] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ea2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03752] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ea4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03753] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ea6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03754] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ea8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03755] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03756] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03757] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03758] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03759] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0375a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0375b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0375c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0375d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0375e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ebc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0375f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ebe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03760] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ec0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03761] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ec2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03762] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ec4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03763] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ec6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03764] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ec8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03765] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03766] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ecc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03767] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ece] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03768] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ed0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03769] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ed2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0376a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ed4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0376b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ed6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0376c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ed8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0376d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0376e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06edc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0376f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ede] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03770] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ee0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03771] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ee2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03772] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ee4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03773] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ee6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03774] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ee8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03775] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03776] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03777] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06eee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03778] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ef0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03779] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ef2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0377a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ef4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0377b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ef6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0377c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ef8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0377d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06efa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0377e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06efc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0377f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06efe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03780] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03781] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03782] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03783] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03784] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03785] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03786] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03787] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03788] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03789] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0378a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0378b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0378c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0378d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0378e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0378f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03790] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03791] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03792] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03793] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03794] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03795] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03796] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03797] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03798] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03799] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0379a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0379b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0379c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0379d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0379e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0379f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06f9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06faa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fe0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fe2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fe4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fe6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fe8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06fee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ff0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ff2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ff4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ff6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ff8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ffa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ffc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h06ffe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03800] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07000] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03801] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07002] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03802] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07004] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03803] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07006] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03804] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07008] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03805] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0700a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03806] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0700c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03807] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0700e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03808] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07010] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03809] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07012] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0380a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07014] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0380b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07016] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0380c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07018] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0380d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0701a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0380e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0701c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0380f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0701e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03810] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07020] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03811] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07022] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03812] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07024] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03813] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07026] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03814] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07028] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03815] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0702a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03816] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0702c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03817] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0702e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03818] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07030] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03819] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07032] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0381a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07034] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0381b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07036] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0381c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07038] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0381d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0703a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0381e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0703c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0381f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0703e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03820] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07040] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03821] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07042] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03822] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07044] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03823] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07046] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03824] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07048] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03825] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0704a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03826] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0704c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03827] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0704e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03828] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07050] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03829] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07052] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0382a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07054] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0382b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07056] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0382c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07058] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0382d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0705a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0382e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0705c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0382f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0705e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03830] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07060] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03831] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07062] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03832] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07064] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03833] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07066] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03834] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07068] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03835] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0706a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03836] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0706c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03837] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0706e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03838] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07070] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03839] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07072] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0383a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07074] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0383b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07076] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0383c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07078] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0383d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0707a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0383e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0707c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0383f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0707e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03840] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07080] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03841] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07082] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03842] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07084] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03843] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07086] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03844] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07088] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03845] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0708a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03846] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0708c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03847] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0708e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03848] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07090] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03849] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07092] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0384a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07094] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0384b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07096] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0384c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07098] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0384d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0709a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0384e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0709c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0384f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0709e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03850] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03851] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03852] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03853] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03854] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03855] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03856] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03857] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03858] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03859] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0385a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0385b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0385c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0385d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0385e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0385f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03860] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03861] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03862] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03863] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03864] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03865] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03866] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03867] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03868] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03869] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0386a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0386b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0386c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0386d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0386e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0386f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03870] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03871] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03872] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03873] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03874] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03875] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03876] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03877] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03878] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03879] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0387a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0387b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0387c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0387d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0387e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0387f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h070fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03880] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07100] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03881] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07102] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03882] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07104] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03883] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07106] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03884] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07108] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03885] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0710a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03886] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0710c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03887] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0710e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03888] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07110] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03889] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07112] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0388a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07114] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0388b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07116] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0388c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07118] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0388d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0711a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0388e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0711c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0388f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0711e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03890] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07120] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03891] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07122] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03892] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07124] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03893] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07126] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03894] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07128] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03895] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0712a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03896] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0712c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03897] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0712e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03898] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07130] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03899] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07132] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0389a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07134] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0389b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07136] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0389c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07138] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0389d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0713a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0389e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0713c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0389f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0713e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07140] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07142] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07144] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07146] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07148] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0714a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0714c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0714e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07150] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07152] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07154] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07156] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07158] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0715a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0715c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0715e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07160] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07162] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07164] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07166] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07168] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0716a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0716c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0716e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07170] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07172] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07174] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07176] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07178] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0717a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0717c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0717e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07180] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07182] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07184] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07186] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07188] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0718a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0718c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0718e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07190] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07192] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07194] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07196] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07198] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0719a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0719c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0719e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h071fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03900] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07200] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03901] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07202] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03902] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07204] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03903] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07206] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03904] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07208] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03905] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0720a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03906] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0720c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03907] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0720e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03908] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07210] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03909] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07212] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0390a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07214] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0390b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07216] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0390c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07218] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0390d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0721a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0390e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0721c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0390f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0721e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03910] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07220] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03911] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07222] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03912] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07224] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03913] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07226] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03914] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07228] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03915] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0722a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03916] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0722c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03917] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0722e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03918] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07230] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03919] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07232] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0391a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07234] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0391b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07236] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0391c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07238] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0391d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0723a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0391e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0723c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0391f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0723e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03920] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07240] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03921] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07242] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03922] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07244] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03923] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07246] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03924] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07248] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03925] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0724a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03926] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0724c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03927] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0724e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03928] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07250] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03929] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07252] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0392a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07254] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0392b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07256] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0392c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07258] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0392d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0725a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0392e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0725c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0392f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0725e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03930] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07260] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03931] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07262] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03932] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07264] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03933] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07266] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03934] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07268] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03935] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0726a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03936] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0726c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03937] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0726e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03938] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07270] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03939] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07272] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0393a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07274] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0393b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07276] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0393c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07278] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0393d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0727a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0393e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0727c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0393f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0727e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03940] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07280] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03941] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07282] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03942] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07284] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03943] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07286] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03944] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07288] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03945] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0728a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03946] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0728c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03947] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0728e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03948] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07290] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03949] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07292] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0394a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07294] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0394b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07296] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0394c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07298] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0394d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0729a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0394e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0729c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0394f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0729e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03950] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03951] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03952] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03953] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03954] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03955] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03956] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03957] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03958] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03959] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0395a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0395b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0395c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0395d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0395e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0395f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03960] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03961] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03962] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03963] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03964] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03965] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03966] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03967] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03968] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03969] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0396a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0396b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0396c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0396d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0396e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0396f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03970] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03971] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03972] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03973] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03974] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03975] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03976] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03977] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03978] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03979] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0397a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0397b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0397c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0397d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0397e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0397f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h072fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03980] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07300] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03981] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07302] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03982] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07304] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03983] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07306] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03984] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07308] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03985] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0730a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03986] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0730c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03987] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0730e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03988] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07310] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03989] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07312] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0398a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07314] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0398b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07316] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0398c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07318] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0398d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0731a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0398e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0731c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0398f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0731e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03990] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07320] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03991] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07322] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03992] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07324] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03993] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07326] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03994] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07328] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03995] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0732a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03996] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0732c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03997] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0732e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03998] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07330] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03999] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07332] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0399a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07334] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0399b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07336] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0399c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07338] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0399d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0733a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0399e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0733c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0399f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0733e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07340] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07342] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07344] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07346] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07348] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0734a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0734c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0734e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07350] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07352] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039aa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07354] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07356] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07358] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0735a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0735c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039af] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0735e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07360] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07362] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07364] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07366] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07368] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0736a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0736c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0736e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07370] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07372] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07374] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039bb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07376] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039bc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07378] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039bd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0737a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039be] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0737c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039bf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0737e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07380] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07382] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07384] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07386] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07388] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0738a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0738c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0738e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07390] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07392] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07394] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039cb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07396] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039cc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07398] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039cd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0739a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0739c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039cf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0739e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039da] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039db] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039dc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039dd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039de] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039df] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039eb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039fa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039fb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039fc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039fd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039fe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h073fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07400] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07402] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07404] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07406] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07408] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0740a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0740c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0740e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07410] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07412] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07414] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07416] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07418] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0741a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0741c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0741e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07420] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07422] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07424] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07426] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07428] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0742a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0742c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0742e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07430] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07432] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07434] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07436] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07438] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0743a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0743c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0743e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07440] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07442] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07444] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07446] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07448] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0744a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0744c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0744e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07450] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07452] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07454] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07456] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07458] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0745a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0745c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0745e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07460] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07462] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07464] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07466] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07468] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0746a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0746c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0746e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07470] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07472] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07474] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07476] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07478] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0747a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0747c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0747e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07480] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07482] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07484] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07486] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07488] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0748a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0748c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0748e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07490] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07492] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07494] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07496] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07498] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0749a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0749c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0749e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h074fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07500] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07502] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07504] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07506] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07508] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0750a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0750c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0750e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07510] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07512] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07514] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07516] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07518] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0751a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0751c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0751e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07520] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07522] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07524] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07526] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07528] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0752a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0752c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0752e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07530] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07532] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07534] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07536] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07538] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0753a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0753c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0753e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07540] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07542] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07544] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07546] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07548] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0754a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0754c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0754e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07550] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07552] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aaa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07554] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07556] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07558] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0755a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0755c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aaf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0755e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07560] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07562] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07564] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07566] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07568] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0756a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0756c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0756e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07570] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07572] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07574] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03abb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07576] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03abc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07578] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03abd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0757a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03abe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0757c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03abf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0757e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07580] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07582] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07584] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07586] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07588] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0758a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0758c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0758e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07590] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07592] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07594] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03acb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07596] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03acc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07598] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03acd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0759a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ace] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0759c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03acf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0759e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ada] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03adb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03adc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03add] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ade] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03adf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aeb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03afa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03afb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03afc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03afd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03afe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h075fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07600] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07602] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07604] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07606] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07608] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0760a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0760c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0760e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07610] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07612] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07614] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07616] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07618] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0761a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0761c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0761e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07620] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07622] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07624] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07626] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07628] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0762a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0762c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0762e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07630] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07632] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07634] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07636] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07638] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0763a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0763c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0763e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07640] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07642] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07644] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07646] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07648] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0764a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0764c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0764e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07650] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07652] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07654] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07656] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07658] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0765a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0765c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0765e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07660] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07662] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07664] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07666] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07668] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0766a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0766c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0766e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07670] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07672] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07674] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07676] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07678] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0767a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0767c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0767e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07680] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07682] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07684] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07686] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07688] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0768a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0768c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0768e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07690] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07692] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07694] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07696] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07698] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0769a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0769c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0769e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h076fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07700] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07702] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07704] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07706] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07708] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0770a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0770c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0770e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07710] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07712] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07714] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07716] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07718] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0771a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0771c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0771e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07720] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07722] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07724] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07726] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07728] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0772a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0772c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0772e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07730] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07732] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07734] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07736] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07738] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0773a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0773c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0773e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07740] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07742] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07744] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07746] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07748] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0774a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0774c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0774e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07750] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07752] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03baa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07754] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07756] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07758] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0775a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0775c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03baf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0775e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07760] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07762] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07764] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07766] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07768] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0776a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0776c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0776e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07770] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07772] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07774] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07776] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07778] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0777a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0777c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0777e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07780] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07782] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07784] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07786] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07788] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0778a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0778c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0778e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07790] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07792] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07794] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07796] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07798] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0779a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0779c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0779e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03beb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h077fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07800] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07802] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07804] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07806] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07808] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0780a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0780c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0780e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07810] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07812] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07814] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07816] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07818] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0781a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0781c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0781e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07820] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07822] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07824] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07826] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07828] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0782a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0782c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0782e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07830] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07832] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07834] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07836] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07838] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0783a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0783c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0783e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07840] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07842] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07844] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07846] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07848] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0784a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0784c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0784e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07850] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07852] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07854] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07856] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07858] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0785a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0785c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0785e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07860] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07862] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07864] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07866] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07868] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0786a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0786c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0786e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07870] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07872] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07874] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07876] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07878] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0787a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0787c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0787e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07880] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07882] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07884] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07886] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07888] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0788a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0788c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0788e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07890] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07892] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07894] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07896] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07898] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0789a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0789c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0789e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h078fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07900] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07902] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07904] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07906] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07908] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0790a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0790c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0790e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07910] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07912] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07914] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07916] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07918] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0791a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0791c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0791e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07920] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07922] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07924] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07926] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07928] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0792a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0792c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0792e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07930] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07932] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07934] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07936] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07938] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0793a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0793c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0793e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07940] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07942] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07944] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07946] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07948] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0794a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0794c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0794e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07950] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07952] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03caa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07954] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07956] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07958] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0795a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0795c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03caf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0795e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07960] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07962] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07964] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07966] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07968] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0796a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0796c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0796e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07970] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07972] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07974] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07976] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07978] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0797a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0797c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0797e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07980] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07982] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07984] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07986] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07988] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0798a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0798c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0798e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07990] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07992] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07994] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ccb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07996] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ccc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07998] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ccd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0799a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0799c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ccf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h0799e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079a0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079a2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079a4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079a6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079a8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079aa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079ac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079ae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079b0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079b2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079b4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079b6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079b8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079ba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079bc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079be] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079c0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079c2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079c4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079c6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079c8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079ca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079cc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079ce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079d0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079d2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079d4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ceb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079d6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079d8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ced] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079da] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079dc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079de] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079e0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079e2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079e4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079e6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079e8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079ea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079ec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079ee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079f0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079f2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079f4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079f6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079f8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079fa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079fc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h079fe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07a9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ab0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ab2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ab4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ab6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ab8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07abc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07abe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ac0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ac2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ac4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ac6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ac8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07acc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ace] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ad0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ad2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ad4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ad6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ad8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ada] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07adc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ade] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ae0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ae2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ae4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ae6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ae8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07aee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07af0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07af2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07af4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07af6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07af8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07afa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07afc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07afe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03daa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03daf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07b9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ba0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ba2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ba4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ba6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ba8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07baa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ddb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ddc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ddd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ddf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03deb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ded] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03def] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07be0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07be2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07be4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07be6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07be8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dfa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dfb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dfc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dfd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dfe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07bfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07c9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ca0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ca2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ca4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ca6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ca8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07caa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ccc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ce0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ce2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ce4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ce6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ce8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cf0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cf2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cf4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cf6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cf8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07cfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eaa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ead] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eaf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ebb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ebc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ebd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ebe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ebf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ecb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ecc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ecd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ece] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ecf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07d9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07da0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07da2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07da4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07da6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07da8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07daa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07db0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07db2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07db4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03edb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07db6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03edc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07db8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03edd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ede] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03edf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eeb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ddc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07de0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07de2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07de4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07de6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07de8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07df0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07df2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03efa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07df4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03efb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07df6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03efc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07df8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03efd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dfa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03efe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dfc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07dfe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f00] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f01] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f02] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f03] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f04] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f05] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f06] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f07] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f08] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f09] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f0a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f0b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f0c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f0d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f0e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f0f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f10] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f11] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f12] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f13] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f14] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f15] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f16] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f17] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f18] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f19] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f1a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f1b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f1c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f1d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f1e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f1f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f20] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f21] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f22] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f23] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f24] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f25] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f26] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f27] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f28] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f29] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f2a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f2b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f2c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f2d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f2e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f2f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f30] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f31] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f32] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f33] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f34] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f35] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f36] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f37] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f38] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f39] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f3a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f3b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f3c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f3d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f3e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f3f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f40] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f41] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f42] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f43] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f44] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f45] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f46] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f47] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f48] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f49] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f4a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f4b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f4c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f4d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f4e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f4f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07e9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f50] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ea0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f51] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ea2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f52] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ea4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f53] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ea6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f54] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ea8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f55] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eaa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f56] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f57] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f58] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f59] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f5a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f5b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f5c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f5d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f5e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ebc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f5f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ebe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f60] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ec0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f61] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ec2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f62] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ec4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f63] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ec6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f64] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ec8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f65] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f66] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ecc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f67] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ece] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f68] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ed0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f69] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ed2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f6a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ed4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f6b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ed6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f6c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ed8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f6d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f6e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07edc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f6f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ede] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f70] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ee0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f71] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ee2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f72] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ee4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f73] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ee6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f74] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ee8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f75] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f76] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f77] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07eee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f78] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ef0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f79] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ef2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f7a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ef4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f7b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ef6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f7c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ef8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f7d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07efa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f7e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07efc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f7f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07efe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f80] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f00] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f81] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f02] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f82] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f04] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f83] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f06] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f84] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f08] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f85] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f0a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f86] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f0c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f87] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f0e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f88] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f10] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f89] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f12] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f8a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f14] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f8b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f16] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f8c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f18] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f8d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f1a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f8e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f1c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f8f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f1e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f90] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f20] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f91] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f22] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f92] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f24] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f93] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f26] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f94] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f28] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f95] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f2a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f96] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f2c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f97] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f2e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f98] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f30] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f99] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f32] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f9a] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f34] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f9b] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f36] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f9c] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f38] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f9d] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f3a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f9e] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f3c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f9f] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f3e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f40] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f42] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f44] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f46] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f48] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f4a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f4c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f4e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f50] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f52] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03faa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f54] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fab] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f56] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fac] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f58] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fad] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f5a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fae] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f5c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03faf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f5e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f60] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f62] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f64] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f66] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f68] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f6a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f6c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f6e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f70] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f72] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fba] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f74] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fbb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f76] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fbc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f78] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fbd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f7a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fbe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f7c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fbf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f7e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f80] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f82] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f84] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f86] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f88] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f8a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f8c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f8e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f90] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f92] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fca] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f94] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fcb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f96] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fcc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f98] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fcd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f9a] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fce] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f9c] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fcf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07f9e] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fa0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fa2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fa4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fa6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fa8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07faa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fac] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fae] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fb0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fb2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fda] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fb4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fdb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fb6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fdc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fb8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fdd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fba] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fde] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fbc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fdf] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fbe] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fc0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fc2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fc4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fc6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fc8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fca] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fcc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fce] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fd0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fd2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fea] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fd4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03feb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fd6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fec] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fd8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fed] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fda] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fee] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fdc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fef] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fde] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff0] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fe0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff1] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fe2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff2] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fe4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff3] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fe6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff4] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fe8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff5] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fea] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff6] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fec] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff7] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07fee] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff8] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ff0] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff9] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ff2] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ffa] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ff4] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ffb] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ff6] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ffc] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ff8] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ffd] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ffa] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ffe] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ffc] ;
//end
//always_comb begin // 
               Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fff] =  I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e['h07ffe] ;
//end
