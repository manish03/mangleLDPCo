parameter n_minus_m = 'd40;
parameter n_int = 'd208;
parameter m_int = 'd168;



parameter z_int = 'd4;



wire [n_int-1:n_int-m_int] Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c; 
wire Iab07a22132333dc82dfd2bb37d146a4afe639be50119ec29071aef525973c414;
assign Iab07a22132333dc82dfd2bb37d146a4afe639be50119ec29071aef525973c414 = 
        y_nr_in[5] ^ 
        y_nr_in[8] ^ 
        y_nr_in[14] ^ 
0; 



wire Iea6de604aaff37b3ef8fe79b4d320861d98645b7eabcc908f78968b998a90023;
assign Iea6de604aaff37b3ef8fe79b4d320861d98645b7eabcc908f78968b998a90023 = 
        y_nr_in[25] ^ 
        y_nr_in[37] ^ 
        y_nr_in[3] ^ 
0; 



wire I79564af2d1f960a0b996143407a5abe6fb627e52634b56529d4d7924ca7d687d;
assign I79564af2d1f960a0b996143407a5abe6fb627e52634b56529d4d7924ca7d687d = 
        y_nr_in[14] ^ 
        y_nr_in[17] ^ 
        y_nr_in[21] ^ 
0; 



wire I0d2cf4e6eef8eec4983f8c40142a8bf8a2ad8bb5c4e10b769d6b5710fec91903;
assign I0d2cf4e6eef8eec4983f8c40142a8bf8a2ad8bb5c4e10b769d6b5710fec91903 = 
        y_nr_in[26] ^ 
        y_nr_in[28] ^ 
        y_nr_in[32] ^ 
0; 



wire Ia31ac86371faab0167761f477dd9e1caa9f77ffa3df023c71820c0be8a855809;
assign Ia31ac86371faab0167761f477dd9e1caa9f77ffa3df023c71820c0be8a855809 = 
        y_nr_in[36] ^ 
        y_nr_in[1] ^ 
        y_nr_in[6] ^ 
0; 



wire I5a69a39df49748f6e56b592cd8fd289e66ca518769bc0ce68fbd1ce750a73cf5;
assign I5a69a39df49748f6e56b592cd8fd289e66ca518769bc0ce68fbd1ce750a73cf5 = 
        y_nr_in[12] ^ 
        y_nr_in[16] ^ 
        y_nr_in[32] ^ 
0; 



wire I46f5ea8015199f30dd79254a3dd0c0af5ae81e6963ab67aa8514881dd27ddd06;
assign I46f5ea8015199f30dd79254a3dd0c0af5ae81e6963ab67aa8514881dd27ddd06 = 
        y_nr_in[4] ^ 
        y_nr_in[10] ^ 
        y_nr_in[18] ^ 
0; 



wire Ida3af96cb68bdec0bafe8f371a9fbe67e45a145a33066d32da8dc3aa39fce8a3;
assign Ida3af96cb68bdec0bafe8f371a9fbe67e45a145a33066d32da8dc3aa39fce8a3 = 
        y_nr_in[20] ^ 
        y_nr_in[25] ^ 
        y_nr_in[30] ^ 
0; 



wire I74cd5c3fac22a70cb1e62c6a3c750e289f5b3d61a2532ac35248579d60f4873d;
assign I74cd5c3fac22a70cb1e62c6a3c750e289f5b3d61a2532ac35248579d60f4873d = 
        y_nr_in[34] ^ 
        y_nr_in[36] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[40] = 
Iab07a22132333dc82dfd2bb37d146a4afe639be50119ec29071aef525973c414 ^ 
Iea6de604aaff37b3ef8fe79b4d320861d98645b7eabcc908f78968b998a90023 ^ 
I79564af2d1f960a0b996143407a5abe6fb627e52634b56529d4d7924ca7d687d ^ 
I0d2cf4e6eef8eec4983f8c40142a8bf8a2ad8bb5c4e10b769d6b5710fec91903 ^ 
Ia31ac86371faab0167761f477dd9e1caa9f77ffa3df023c71820c0be8a855809 ^ 
I5a69a39df49748f6e56b592cd8fd289e66ca518769bc0ce68fbd1ce750a73cf5 ^ 
I46f5ea8015199f30dd79254a3dd0c0af5ae81e6963ab67aa8514881dd27ddd06 ^ 
Ida3af96cb68bdec0bafe8f371a9fbe67e45a145a33066d32da8dc3aa39fce8a3 ^ 
I74cd5c3fac22a70cb1e62c6a3c750e289f5b3d61a2532ac35248579d60f4873d ^ 
0; 



wire I1021f3960dc6d9dbead5d89ab46837450094ec1eb9995a54c3e035bc39b41e39;
assign I1021f3960dc6d9dbead5d89ab46837450094ec1eb9995a54c3e035bc39b41e39 = 
        y_nr_in[6] ^ 
        y_nr_in[9] ^ 
        y_nr_in[15] ^ 
0; 



wire I2c44abec3d29ee6fe5d6b31783f0aa93300b8534802a8a09b2a70d23719b743b;
assign I2c44abec3d29ee6fe5d6b31783f0aa93300b8534802a8a09b2a70d23719b743b = 
        y_nr_in[26] ^ 
        y_nr_in[38] ^ 
        y_nr_in[0] ^ 
0; 



wire Iad3150ccb063c396b66bffa8ffe6ed7034dd22e361d207954a4805775a4fb0ad;
assign Iad3150ccb063c396b66bffa8ffe6ed7034dd22e361d207954a4805775a4fb0ad = 
        y_nr_in[15] ^ 
        y_nr_in[18] ^ 
        y_nr_in[22] ^ 
0; 



wire I3b355fb597cfc8011e4fd3e31e10c5c2ceb948868606d39ae15ce5d5744d79a8;
assign I3b355fb597cfc8011e4fd3e31e10c5c2ceb948868606d39ae15ce5d5744d79a8 = 
        y_nr_in[27] ^ 
        y_nr_in[29] ^ 
        y_nr_in[33] ^ 
0; 



wire Ib156d16e1883853f9afe96b67e6067ff6ff3f63bc2766ab997ad153d57f7ad5a;
assign Ib156d16e1883853f9afe96b67e6067ff6ff3f63bc2766ab997ad153d57f7ad5a = 
        y_nr_in[37] ^ 
        y_nr_in[2] ^ 
        y_nr_in[7] ^ 
0; 



wire I0383243d7b7304219092aca387e7dcc02a3ed24cb8912177be8316c7f6fb7f25;
assign I0383243d7b7304219092aca387e7dcc02a3ed24cb8912177be8316c7f6fb7f25 = 
        y_nr_in[13] ^ 
        y_nr_in[17] ^ 
        y_nr_in[33] ^ 
0; 



wire I95c9f9357b036b5293f8475587502bb6c20b40d5144bdfb61b1912ce61206585;
assign I95c9f9357b036b5293f8475587502bb6c20b40d5144bdfb61b1912ce61206585 = 
        y_nr_in[5] ^ 
        y_nr_in[11] ^ 
        y_nr_in[19] ^ 
0; 



wire Ida8b63aa236a3a46d40657291702f887f60f1c648d85eb7d4b7e4c14699089cc;
assign Ida8b63aa236a3a46d40657291702f887f60f1c648d85eb7d4b7e4c14699089cc = 
        y_nr_in[21] ^ 
        y_nr_in[26] ^ 
        y_nr_in[31] ^ 
0; 



wire Ib8158ac56db5224bad0c42449015c8e3bcdae41a1cdc91dfb8a31edafe6f130a;
assign Ib8158ac56db5224bad0c42449015c8e3bcdae41a1cdc91dfb8a31edafe6f130a = 
        y_nr_in[35] ^ 
        y_nr_in[37] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[41] = 
I1021f3960dc6d9dbead5d89ab46837450094ec1eb9995a54c3e035bc39b41e39 ^ 
I2c44abec3d29ee6fe5d6b31783f0aa93300b8534802a8a09b2a70d23719b743b ^ 
Iad3150ccb063c396b66bffa8ffe6ed7034dd22e361d207954a4805775a4fb0ad ^ 
I3b355fb597cfc8011e4fd3e31e10c5c2ceb948868606d39ae15ce5d5744d79a8 ^ 
Ib156d16e1883853f9afe96b67e6067ff6ff3f63bc2766ab997ad153d57f7ad5a ^ 
I0383243d7b7304219092aca387e7dcc02a3ed24cb8912177be8316c7f6fb7f25 ^ 
I95c9f9357b036b5293f8475587502bb6c20b40d5144bdfb61b1912ce61206585 ^ 
Ida8b63aa236a3a46d40657291702f887f60f1c648d85eb7d4b7e4c14699089cc ^ 
Ib8158ac56db5224bad0c42449015c8e3bcdae41a1cdc91dfb8a31edafe6f130a ^ 
0; 



wire I14bcc7037579859fb0b78322d661a77583d6954f553bf1c312da3edfc4aea4d6;
assign I14bcc7037579859fb0b78322d661a77583d6954f553bf1c312da3edfc4aea4d6 = 
        y_nr_in[7] ^ 
        y_nr_in[10] ^ 
        y_nr_in[12] ^ 
0; 



wire Icb15408687f0a3019efd733726eccdc9cde4e2bc819c47c2a1259c7d20457388;
assign Icb15408687f0a3019efd733726eccdc9cde4e2bc819c47c2a1259c7d20457388 = 
        y_nr_in[27] ^ 
        y_nr_in[39] ^ 
        y_nr_in[1] ^ 
0; 



wire I4d1a5af2946924d8ab30ab7c3469aecf069b5ef7aebca19adb09c9076ce029c3;
assign I4d1a5af2946924d8ab30ab7c3469aecf069b5ef7aebca19adb09c9076ce029c3 = 
        y_nr_in[12] ^ 
        y_nr_in[19] ^ 
        y_nr_in[23] ^ 
0; 



wire Ie44d088557dea31d11e2ee8c893fd0e23048af601f482de92f5eb30196be2d10;
assign Ie44d088557dea31d11e2ee8c893fd0e23048af601f482de92f5eb30196be2d10 = 
        y_nr_in[24] ^ 
        y_nr_in[30] ^ 
        y_nr_in[34] ^ 
0; 



wire I2b23350d74b2188a4798cfbf7451eb61ef9f289796e0a83e0f026959946cb5d5;
assign I2b23350d74b2188a4798cfbf7451eb61ef9f289796e0a83e0f026959946cb5d5 = 
        y_nr_in[38] ^ 
        y_nr_in[3] ^ 
        y_nr_in[4] ^ 
0; 



wire Ief1a245cc840afe888b40f74314d5401197a4b1caacefca72781e5475b58351b;
assign Ief1a245cc840afe888b40f74314d5401197a4b1caacefca72781e5475b58351b = 
        y_nr_in[14] ^ 
        y_nr_in[18] ^ 
        y_nr_in[34] ^ 
0; 



wire I179125003da12b3a72a65fca1f1f568214da36fee73fb0ccc0834fc1414b5725;
assign I179125003da12b3a72a65fca1f1f568214da36fee73fb0ccc0834fc1414b5725 = 
        y_nr_in[6] ^ 
        y_nr_in[8] ^ 
        y_nr_in[16] ^ 
0; 



wire I12c5704853780c2806dcded4d1ed50c68a15c8076b28f799bebc5ef12152e03b;
assign I12c5704853780c2806dcded4d1ed50c68a15c8076b28f799bebc5ef12152e03b = 
        y_nr_in[22] ^ 
        y_nr_in[27] ^ 
        y_nr_in[28] ^ 
0; 



wire If61fb2374651687574f1c4cf226ba7095f37daffe5f379de72fce155400baf22;
assign If61fb2374651687574f1c4cf226ba7095f37daffe5f379de72fce155400baf22 = 
        y_nr_in[32] ^ 
        y_nr_in[38] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[42] = 
I14bcc7037579859fb0b78322d661a77583d6954f553bf1c312da3edfc4aea4d6 ^ 
Icb15408687f0a3019efd733726eccdc9cde4e2bc819c47c2a1259c7d20457388 ^ 
I4d1a5af2946924d8ab30ab7c3469aecf069b5ef7aebca19adb09c9076ce029c3 ^ 
Ie44d088557dea31d11e2ee8c893fd0e23048af601f482de92f5eb30196be2d10 ^ 
I2b23350d74b2188a4798cfbf7451eb61ef9f289796e0a83e0f026959946cb5d5 ^ 
Ief1a245cc840afe888b40f74314d5401197a4b1caacefca72781e5475b58351b ^ 
I179125003da12b3a72a65fca1f1f568214da36fee73fb0ccc0834fc1414b5725 ^ 
I12c5704853780c2806dcded4d1ed50c68a15c8076b28f799bebc5ef12152e03b ^ 
If61fb2374651687574f1c4cf226ba7095f37daffe5f379de72fce155400baf22 ^ 
0; 



wire I3e6bdfbaa1119c206b79fa1bd1482b00ec49e9faaf6fe9e6cc7a26d0e0cf5601;
assign I3e6bdfbaa1119c206b79fa1bd1482b00ec49e9faaf6fe9e6cc7a26d0e0cf5601 = 
        y_nr_in[4] ^ 
        y_nr_in[11] ^ 
        y_nr_in[13] ^ 
0; 



wire I65f788fc8443ed1153c2ec1b5043e0f11c4264879a28e67d456d0f7decdde271;
assign I65f788fc8443ed1153c2ec1b5043e0f11c4264879a28e67d456d0f7decdde271 = 
        y_nr_in[24] ^ 
        y_nr_in[36] ^ 
        y_nr_in[2] ^ 
0; 



wire I4ea77074b68c91fa0d20c29c36885a631cabcf530cf459379fec1a8f876cc4e0;
assign I4ea77074b68c91fa0d20c29c36885a631cabcf530cf459379fec1a8f876cc4e0 = 
        y_nr_in[13] ^ 
        y_nr_in[16] ^ 
        y_nr_in[20] ^ 
0; 



wire Idaa6056608bfae5be4c691c8236600735a7529cc581a0f3c8941fec85273f767;
assign Idaa6056608bfae5be4c691c8236600735a7529cc581a0f3c8941fec85273f767 = 
        y_nr_in[25] ^ 
        y_nr_in[31] ^ 
        y_nr_in[35] ^ 
0; 



wire If8110a0237ea795b56b187b217ebf3ab7960cbc72234624a4f80505ed600693d;
assign If8110a0237ea795b56b187b217ebf3ab7960cbc72234624a4f80505ed600693d = 
        y_nr_in[39] ^ 
        y_nr_in[0] ^ 
        y_nr_in[5] ^ 
0; 



wire I35f7038c24558f6a440829bc74531b01ee21dacbaf1606582e2d5919c1e64796;
assign I35f7038c24558f6a440829bc74531b01ee21dacbaf1606582e2d5919c1e64796 = 
        y_nr_in[15] ^ 
        y_nr_in[19] ^ 
        y_nr_in[35] ^ 
0; 



wire Iae14b788a61d774755daa8f1a666263d5bc53eaf1c340a98f2eeb3147e99ed11;
assign Iae14b788a61d774755daa8f1a666263d5bc53eaf1c340a98f2eeb3147e99ed11 = 
        y_nr_in[7] ^ 
        y_nr_in[9] ^ 
        y_nr_in[17] ^ 
0; 



wire I99da4d46716d5fc981448b5a4b0bf9ed7753abd84678a6d9e6551d95f6610aed;
assign I99da4d46716d5fc981448b5a4b0bf9ed7753abd84678a6d9e6551d95f6610aed = 
        y_nr_in[23] ^ 
        y_nr_in[24] ^ 
        y_nr_in[29] ^ 
0; 



wire I5060342870576d2e4bba1f9eea4fef4004116611da636b27d986b3da38ede3ff;
assign I5060342870576d2e4bba1f9eea4fef4004116611da636b27d986b3da38ede3ff = 
        y_nr_in[33] ^ 
        y_nr_in[39] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[43] = 
I3e6bdfbaa1119c206b79fa1bd1482b00ec49e9faaf6fe9e6cc7a26d0e0cf5601 ^ 
I65f788fc8443ed1153c2ec1b5043e0f11c4264879a28e67d456d0f7decdde271 ^ 
I4ea77074b68c91fa0d20c29c36885a631cabcf530cf459379fec1a8f876cc4e0 ^ 
Idaa6056608bfae5be4c691c8236600735a7529cc581a0f3c8941fec85273f767 ^ 
If8110a0237ea795b56b187b217ebf3ab7960cbc72234624a4f80505ed600693d ^ 
I35f7038c24558f6a440829bc74531b01ee21dacbaf1606582e2d5919c1e64796 ^ 
Iae14b788a61d774755daa8f1a666263d5bc53eaf1c340a98f2eeb3147e99ed11 ^ 
I99da4d46716d5fc981448b5a4b0bf9ed7753abd84678a6d9e6551d95f6610aed ^ 
I5060342870576d2e4bba1f9eea4fef4004116611da636b27d986b3da38ede3ff ^ 
0; 



wire I4ec3b7ee477264f3d1c336bd00d2fabb40f0116218727e3619709e1296468c24;
assign I4ec3b7ee477264f3d1c336bd00d2fabb40f0116218727e3619709e1296468c24 = 
        y_nr_in[5] ^ 
        y_nr_in[8] ^ 
        y_nr_in[14] ^ 
0; 



wire Ieceddce637e91b17dcdf72e43b0eeacc0af6b3c8983e8863316bf68711130abf;
assign Ieceddce637e91b17dcdf72e43b0eeacc0af6b3c8983e8863316bf68711130abf = 
        y_nr_in[25] ^ 
        y_nr_in[37] ^ 
        y_nr_in[40] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[44] = 
I4ec3b7ee477264f3d1c336bd00d2fabb40f0116218727e3619709e1296468c24 ^ 
Ieceddce637e91b17dcdf72e43b0eeacc0af6b3c8983e8863316bf68711130abf ^ 
0; 



wire Idcdd8b778353d44d370a1a3ebac9cda0d67cfe850715e86fdf4aa07c5711a951;
assign Idcdd8b778353d44d370a1a3ebac9cda0d67cfe850715e86fdf4aa07c5711a951 = 
        y_nr_in[6] ^ 
        y_nr_in[9] ^ 
        y_nr_in[15] ^ 
0; 



wire If21d6269cf0a04b6ab675023508e3e7df981656e5426ac641504f414efc97789;
assign If21d6269cf0a04b6ab675023508e3e7df981656e5426ac641504f414efc97789 = 
        y_nr_in[26] ^ 
        y_nr_in[38] ^ 
        y_nr_in[41] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[45] = 
Idcdd8b778353d44d370a1a3ebac9cda0d67cfe850715e86fdf4aa07c5711a951 ^ 
If21d6269cf0a04b6ab675023508e3e7df981656e5426ac641504f414efc97789 ^ 
0; 



wire I89d0a135e12a1d3e58ab85368e7b060daafc1fc9debfd29b3faffb2b94fcc86f;
assign I89d0a135e12a1d3e58ab85368e7b060daafc1fc9debfd29b3faffb2b94fcc86f = 
        y_nr_in[7] ^ 
        y_nr_in[10] ^ 
        y_nr_in[12] ^ 
0; 



wire I38239b6ab86f4ff40dff1abeb52aacc9694eba64eebab8322f0d15fca272c9d3;
assign I38239b6ab86f4ff40dff1abeb52aacc9694eba64eebab8322f0d15fca272c9d3 = 
        y_nr_in[27] ^ 
        y_nr_in[39] ^ 
        y_nr_in[42] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[46] = 
I89d0a135e12a1d3e58ab85368e7b060daafc1fc9debfd29b3faffb2b94fcc86f ^ 
I38239b6ab86f4ff40dff1abeb52aacc9694eba64eebab8322f0d15fca272c9d3 ^ 
0; 



wire I858df6bb38a70d9caf8b447cfe0dfbb9cb9bd24e9f42adc59d561e8e7425ef35;
assign I858df6bb38a70d9caf8b447cfe0dfbb9cb9bd24e9f42adc59d561e8e7425ef35 = 
        y_nr_in[4] ^ 
        y_nr_in[11] ^ 
        y_nr_in[13] ^ 
0; 



wire I3cbddc8bfb69bb229bbc8084504f4d2d9b07f3cdfa924d0cce6b3c57a8ad8307;
assign I3cbddc8bfb69bb229bbc8084504f4d2d9b07f3cdfa924d0cce6b3c57a8ad8307 = 
        y_nr_in[24] ^ 
        y_nr_in[36] ^ 
        y_nr_in[43] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[47] = 
I858df6bb38a70d9caf8b447cfe0dfbb9cb9bd24e9f42adc59d561e8e7425ef35 ^ 
I3cbddc8bfb69bb229bbc8084504f4d2d9b07f3cdfa924d0cce6b3c57a8ad8307 ^ 
0; 



wire I68ab23a12dceb8cda9709ed2a8e2988caa47f0fc29e1ff33f3b8940e4d5116ad;
assign I68ab23a12dceb8cda9709ed2a8e2988caa47f0fc29e1ff33f3b8940e4d5116ad = 
        y_nr_in[3] ^ 
        y_nr_in[14] ^ 
        y_nr_in[17] ^ 
0; 



wire I30de6e6f3e76be1eb1109eb87f7b26ddf13dc14903e3757353eb1280f5b16129;
assign I30de6e6f3e76be1eb1109eb87f7b26ddf13dc14903e3757353eb1280f5b16129 = 
        y_nr_in[21] ^ 
        y_nr_in[26] ^ 
        y_nr_in[28] ^ 
0; 



wire I4d4c5d7a5f9ec94d1944c9bc64c21e72de8d369c2175834ffc38f5dfe7f0ecbc;
assign I4d4c5d7a5f9ec94d1944c9bc64c21e72de8d369c2175834ffc38f5dfe7f0ecbc = 
        y_nr_in[32] ^ 
        y_nr_in[36] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[48] = 
I68ab23a12dceb8cda9709ed2a8e2988caa47f0fc29e1ff33f3b8940e4d5116ad ^ 
I30de6e6f3e76be1eb1109eb87f7b26ddf13dc14903e3757353eb1280f5b16129 ^ 
I4d4c5d7a5f9ec94d1944c9bc64c21e72de8d369c2175834ffc38f5dfe7f0ecbc ^ 
0; 



wire Ib60fade8c09d8680a36e5bf1a0284b796673a17e94a819251f2a71e15295fa3b;
assign Ib60fade8c09d8680a36e5bf1a0284b796673a17e94a819251f2a71e15295fa3b = 
        y_nr_in[0] ^ 
        y_nr_in[15] ^ 
        y_nr_in[18] ^ 
0; 



wire I9320ae9c560a5fa7618f9c1a2e0928bd597fae2df6bbcd0f016a3cbf53c7e5bd;
assign I9320ae9c560a5fa7618f9c1a2e0928bd597fae2df6bbcd0f016a3cbf53c7e5bd = 
        y_nr_in[22] ^ 
        y_nr_in[27] ^ 
        y_nr_in[29] ^ 
0; 



wire I4d8a658a9ee5bb4179af98ec2f44aa9aa3a913439259ed20bc954ed05507fe77;
assign I4d8a658a9ee5bb4179af98ec2f44aa9aa3a913439259ed20bc954ed05507fe77 = 
        y_nr_in[33] ^ 
        y_nr_in[37] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[49] = 
Ib60fade8c09d8680a36e5bf1a0284b796673a17e94a819251f2a71e15295fa3b ^ 
I9320ae9c560a5fa7618f9c1a2e0928bd597fae2df6bbcd0f016a3cbf53c7e5bd ^ 
I4d8a658a9ee5bb4179af98ec2f44aa9aa3a913439259ed20bc954ed05507fe77 ^ 
0; 



wire Ibdf7ebe201cc10bc9e3809cf2240498e771574655b7f896bbfad6ee92aca8a23;
assign Ibdf7ebe201cc10bc9e3809cf2240498e771574655b7f896bbfad6ee92aca8a23 = 
        y_nr_in[1] ^ 
        y_nr_in[12] ^ 
        y_nr_in[19] ^ 
0; 



wire Ia1e4adca904053c0bb484052b149e3294bb6eabdd7949a87ea22569021c731e7;
assign Ia1e4adca904053c0bb484052b149e3294bb6eabdd7949a87ea22569021c731e7 = 
        y_nr_in[23] ^ 
        y_nr_in[24] ^ 
        y_nr_in[30] ^ 
0; 



wire I6185cea71d367209dcbaaed784f980bccfce35299bf861aa3200942f49b0d02d;
assign I6185cea71d367209dcbaaed784f980bccfce35299bf861aa3200942f49b0d02d = 
        y_nr_in[34] ^ 
        y_nr_in[38] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[50] = 
Ibdf7ebe201cc10bc9e3809cf2240498e771574655b7f896bbfad6ee92aca8a23 ^ 
Ia1e4adca904053c0bb484052b149e3294bb6eabdd7949a87ea22569021c731e7 ^ 
I6185cea71d367209dcbaaed784f980bccfce35299bf861aa3200942f49b0d02d ^ 
0; 



wire Iaa7fcac337b655b01c8c08546d9e383ead46575b522ed4a4355628ba67ca4fb1;
assign Iaa7fcac337b655b01c8c08546d9e383ead46575b522ed4a4355628ba67ca4fb1 = 
        y_nr_in[2] ^ 
        y_nr_in[13] ^ 
        y_nr_in[16] ^ 
0; 



wire I23c894d4e3c2edc79f5908165fc3b87646e64d996e0ae4798d87a1d86e8726bd;
assign I23c894d4e3c2edc79f5908165fc3b87646e64d996e0ae4798d87a1d86e8726bd = 
        y_nr_in[20] ^ 
        y_nr_in[25] ^ 
        y_nr_in[31] ^ 
0; 



wire I6509c316d67bf9ff5e90f1e631beaf563265c11130e1bad2767b88ddb7de623a;
assign I6509c316d67bf9ff5e90f1e631beaf563265c11130e1bad2767b88ddb7de623a = 
        y_nr_in[35] ^ 
        y_nr_in[39] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[51] = 
Iaa7fcac337b655b01c8c08546d9e383ead46575b522ed4a4355628ba67ca4fb1 ^ 
I23c894d4e3c2edc79f5908165fc3b87646e64d996e0ae4798d87a1d86e8726bd ^ 
I6509c316d67bf9ff5e90f1e631beaf563265c11130e1bad2767b88ddb7de623a ^ 
0; 



wire Ifbe4a51ca6a0ff79d51706849ccac91d91013bf1d4c10860f9c09fec7d7acaf8;
assign Ifbe4a51ca6a0ff79d51706849ccac91d91013bf1d4c10860f9c09fec7d7acaf8 = 
        y_nr_in[1] ^ 
        y_nr_in[6] ^ 
        y_nr_in[12] ^ 
0; 



wire I63d4a749a2da42615978e61d57f01af3334adac002ceadfb9a4f834d56fbc4bc;
assign I63d4a749a2da42615978e61d57f01af3334adac002ceadfb9a4f834d56fbc4bc = 
        y_nr_in[16] ^ 
        y_nr_in[32] ^ 
        y_nr_in[41] ^ 
0; 



wire I065f1c1fa92148d8a8e97d6de75afae5ac42cfba572350bd15cf60b60294a55e;
assign I065f1c1fa92148d8a8e97d6de75afae5ac42cfba572350bd15cf60b60294a55e = 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[52] = 
Ifbe4a51ca6a0ff79d51706849ccac91d91013bf1d4c10860f9c09fec7d7acaf8 ^ 
I63d4a749a2da42615978e61d57f01af3334adac002ceadfb9a4f834d56fbc4bc ^ 
I065f1c1fa92148d8a8e97d6de75afae5ac42cfba572350bd15cf60b60294a55e ^ 
0; 



wire I85e3a5446ecf87fa69161582b8d2570fffbf6166b18f3e3fb7dab2b3934173c6;
assign I85e3a5446ecf87fa69161582b8d2570fffbf6166b18f3e3fb7dab2b3934173c6 = 
        y_nr_in[2] ^ 
        y_nr_in[7] ^ 
        y_nr_in[13] ^ 
0; 



wire I0cffe790d64c26837cbba6f717923aadc0327bb17cd72c189116df14c4b1fb7c;
assign I0cffe790d64c26837cbba6f717923aadc0327bb17cd72c189116df14c4b1fb7c = 
        y_nr_in[17] ^ 
        y_nr_in[33] ^ 
        y_nr_in[42] ^ 
0; 



wire Ide7d97a170efe804f9382f41dc808e00c035c07ccf99ecfa96dbeef17dce5b4a;
assign Ide7d97a170efe804f9382f41dc808e00c035c07ccf99ecfa96dbeef17dce5b4a = 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[53] = 
I85e3a5446ecf87fa69161582b8d2570fffbf6166b18f3e3fb7dab2b3934173c6 ^ 
I0cffe790d64c26837cbba6f717923aadc0327bb17cd72c189116df14c4b1fb7c ^ 
Ide7d97a170efe804f9382f41dc808e00c035c07ccf99ecfa96dbeef17dce5b4a ^ 
0; 



wire I3e60785d78abce1e17afa451061f2c16cf218fde5959c5b8c3773cdfefb00357;
assign I3e60785d78abce1e17afa451061f2c16cf218fde5959c5b8c3773cdfefb00357 = 
        y_nr_in[3] ^ 
        y_nr_in[4] ^ 
        y_nr_in[14] ^ 
0; 



wire Ic8cd56e758a6b346f6030dcfd7ec51cd1be5fe180e3c1eb97490ff1ad9437f70;
assign Ic8cd56e758a6b346f6030dcfd7ec51cd1be5fe180e3c1eb97490ff1ad9437f70 = 
        y_nr_in[18] ^ 
        y_nr_in[34] ^ 
        y_nr_in[43] ^ 
0; 



wire I4df28361fa0a7a8aa895f8db68419f0c9add226d1848577e3fbc5627a8c0ae7d;
assign I4df28361fa0a7a8aa895f8db68419f0c9add226d1848577e3fbc5627a8c0ae7d = 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[54] = 
I3e60785d78abce1e17afa451061f2c16cf218fde5959c5b8c3773cdfefb00357 ^ 
Ic8cd56e758a6b346f6030dcfd7ec51cd1be5fe180e3c1eb97490ff1ad9437f70 ^ 
I4df28361fa0a7a8aa895f8db68419f0c9add226d1848577e3fbc5627a8c0ae7d ^ 
0; 



wire Ib6f4d9266a6f14fc6caf20815aa51585d46b9bb64cbc3583614a9f47a04aedc5;
assign Ib6f4d9266a6f14fc6caf20815aa51585d46b9bb64cbc3583614a9f47a04aedc5 = 
        y_nr_in[0] ^ 
        y_nr_in[5] ^ 
        y_nr_in[15] ^ 
0; 



wire I09137be6f84d69fc679ceb6395d173bb214f2c3f73d489eb0f8c791768704bc6;
assign I09137be6f84d69fc679ceb6395d173bb214f2c3f73d489eb0f8c791768704bc6 = 
        y_nr_in[19] ^ 
        y_nr_in[35] ^ 
        y_nr_in[40] ^ 
0; 



wire I5fe33ad68de87bff766adbe2ae2f6fbbb5652577746d2087785d2e9330459691;
assign I5fe33ad68de87bff766adbe2ae2f6fbbb5652577746d2087785d2e9330459691 = 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[55] = 
Ib6f4d9266a6f14fc6caf20815aa51585d46b9bb64cbc3583614a9f47a04aedc5 ^ 
I09137be6f84d69fc679ceb6395d173bb214f2c3f73d489eb0f8c791768704bc6 ^ 
I5fe33ad68de87bff766adbe2ae2f6fbbb5652577746d2087785d2e9330459691 ^ 
0; 



wire Ia89469f2c045394fd67fc5894edf5a18e01cec8b06d2330030b2650a1ac75095;
assign Ia89469f2c045394fd67fc5894edf5a18e01cec8b06d2330030b2650a1ac75095 = 
        y_nr_in[3] ^ 
        y_nr_in[6] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[56] = 
Ia89469f2c045394fd67fc5894edf5a18e01cec8b06d2330030b2650a1ac75095 ^ 
0; 



wire I615148ffa13066e02286c8fe3cb5e02104938f716f63286ea03a31309b5ef87d;
assign I615148ffa13066e02286c8fe3cb5e02104938f716f63286ea03a31309b5ef87d = 
        y_nr_in[0] ^ 
        y_nr_in[7] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[57] = 
I615148ffa13066e02286c8fe3cb5e02104938f716f63286ea03a31309b5ef87d ^ 
0; 



wire Ie963a8840cb2771f615bd29bc69d572a2992b1ae6391979fff65625d8a31cc8f;
assign Ie963a8840cb2771f615bd29bc69d572a2992b1ae6391979fff65625d8a31cc8f = 
        y_nr_in[1] ^ 
        y_nr_in[4] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[58] = 
Ie963a8840cb2771f615bd29bc69d572a2992b1ae6391979fff65625d8a31cc8f ^ 
0; 



wire Ie77f954a2c57942bfa06d607d78ea178a615bf38c160431bff53683987a1fed5;
assign Ie77f954a2c57942bfa06d607d78ea178a615bf38c160431bff53683987a1fed5 = 
        y_nr_in[2] ^ 
        y_nr_in[5] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[59] = 
Ie77f954a2c57942bfa06d607d78ea178a615bf38c160431bff53683987a1fed5 ^ 
0; 



wire I57ae842a4001d14a9ead5fbdda7ed281087e3d9c6a838e9f23d583e7b9580d3e;
assign I57ae842a4001d14a9ead5fbdda7ed281087e3d9c6a838e9f23d583e7b9580d3e = 
        y_nr_in[3] ^ 
        y_nr_in[5] ^ 
        y_nr_in[22] ^ 
0; 



wire I2372eae8be20255d9196b8eaca424420614b1fcb506174c9dbaf33d47fcc0584;
assign I2372eae8be20255d9196b8eaca424420614b1fcb506174c9dbaf33d47fcc0584 = 
        y_nr_in[31] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[60] = 
I57ae842a4001d14a9ead5fbdda7ed281087e3d9c6a838e9f23d583e7b9580d3e ^ 
I2372eae8be20255d9196b8eaca424420614b1fcb506174c9dbaf33d47fcc0584 ^ 
0; 



wire I53fbf7ceacac2cb4382d381d1397bf17070108bbca2a2a7f6c5c74ea262c0efd;
assign I53fbf7ceacac2cb4382d381d1397bf17070108bbca2a2a7f6c5c74ea262c0efd = 
        y_nr_in[0] ^ 
        y_nr_in[6] ^ 
        y_nr_in[23] ^ 
0; 



wire Iee963cac29e88334eec5d027674ef03159de83d4deed1fde3debd840e986cdb2;
assign Iee963cac29e88334eec5d027674ef03159de83d4deed1fde3debd840e986cdb2 = 
        y_nr_in[28] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[61] = 
I53fbf7ceacac2cb4382d381d1397bf17070108bbca2a2a7f6c5c74ea262c0efd ^ 
Iee963cac29e88334eec5d027674ef03159de83d4deed1fde3debd840e986cdb2 ^ 
0; 



wire Icbbd64503e6a0d82ec8627bebd70e7b3d0781e378b46fe8deefc4aae0f552c1c;
assign Icbbd64503e6a0d82ec8627bebd70e7b3d0781e378b46fe8deefc4aae0f552c1c = 
        y_nr_in[1] ^ 
        y_nr_in[7] ^ 
        y_nr_in[20] ^ 
0; 



wire I286072f35d8290d6c8e9e3def951d8acd165dee25d8e779a61db19f19f669b1d;
assign I286072f35d8290d6c8e9e3def951d8acd165dee25d8e779a61db19f19f669b1d = 
        y_nr_in[29] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[62] = 
Icbbd64503e6a0d82ec8627bebd70e7b3d0781e378b46fe8deefc4aae0f552c1c ^ 
I286072f35d8290d6c8e9e3def951d8acd165dee25d8e779a61db19f19f669b1d ^ 
0; 



wire Ie80a6a85ea5a89ff4d07c8d0f73db32f967fae4ce8c4d7d08a0588ea9f1f8690;
assign Ie80a6a85ea5a89ff4d07c8d0f73db32f967fae4ce8c4d7d08a0588ea9f1f8690 = 
        y_nr_in[2] ^ 
        y_nr_in[4] ^ 
        y_nr_in[21] ^ 
0; 



wire I2ba5ef033b7b82351761dff13dfefd872c97b8685a5d1bc784b4bf02d6c87d39;
assign I2ba5ef033b7b82351761dff13dfefd872c97b8685a5d1bc784b4bf02d6c87d39 = 
        y_nr_in[30] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[63] = 
Ie80a6a85ea5a89ff4d07c8d0f73db32f967fae4ce8c4d7d08a0588ea9f1f8690 ^ 
I2ba5ef033b7b82351761dff13dfefd872c97b8685a5d1bc784b4bf02d6c87d39 ^ 
0; 



wire I36f163a586d548d9b2289c99f0ee152ce6af33124f04fdc15b7934eb27e80e57;
assign I36f163a586d548d9b2289c99f0ee152ce6af33124f04fdc15b7934eb27e80e57 = 
        y_nr_in[3] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
0; 



wire I808cb4ae6f2ba0af20803f85b5d1545aec5eb2df38c6ab5ffa8e35082b4a3c04;
assign I808cb4ae6f2ba0af20803f85b5d1545aec5eb2df38c6ab5ffa8e35082b4a3c04 = 
        y_nr_in[36] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[64] = 
I36f163a586d548d9b2289c99f0ee152ce6af33124f04fdc15b7934eb27e80e57 ^ 
I808cb4ae6f2ba0af20803f85b5d1545aec5eb2df38c6ab5ffa8e35082b4a3c04 ^ 
0; 



wire Ib8ca8cb082f23a8576f5be9d860e817e4b4b743a50e7acb71d670fd34eb3a757;
assign Ib8ca8cb082f23a8576f5be9d860e817e4b4b743a50e7acb71d670fd34eb3a757 = 
        y_nr_in[0] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
0; 



wire If6f14239e9773fee0a9e8a8774d66890cf2673d753a562014ff7410ff024ccc6;
assign If6f14239e9773fee0a9e8a8774d66890cf2673d753a562014ff7410ff024ccc6 = 
        y_nr_in[37] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[65] = 
Ib8ca8cb082f23a8576f5be9d860e817e4b4b743a50e7acb71d670fd34eb3a757 ^ 
If6f14239e9773fee0a9e8a8774d66890cf2673d753a562014ff7410ff024ccc6 ^ 
0; 



wire I596474d97feb75010bbe35074c3d27ab53abab03c5f847dde9ed7e12c18a06b3;
assign I596474d97feb75010bbe35074c3d27ab53abab03c5f847dde9ed7e12c18a06b3 = 
        y_nr_in[1] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
0; 



wire I79bb23a7cece0720233c04f1b17cf33245cb734060f09fb48d6d4b616aa1a18b;
assign I79bb23a7cece0720233c04f1b17cf33245cb734060f09fb48d6d4b616aa1a18b = 
        y_nr_in[38] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[66] = 
I596474d97feb75010bbe35074c3d27ab53abab03c5f847dde9ed7e12c18a06b3 ^ 
I79bb23a7cece0720233c04f1b17cf33245cb734060f09fb48d6d4b616aa1a18b ^ 
0; 



wire I1ab665c6065ef3648ba7c3f60490950063786ffa51ecfe072b7b742287e40e08;
assign I1ab665c6065ef3648ba7c3f60490950063786ffa51ecfe072b7b742287e40e08 = 
        y_nr_in[2] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
0; 



wire I10323882c29157f609df5db826348e4bae6940d64129ac87b330976a2fe64027;
assign I10323882c29157f609df5db826348e4bae6940d64129ac87b330976a2fe64027 = 
        y_nr_in[39] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[67] = 
I1ab665c6065ef3648ba7c3f60490950063786ffa51ecfe072b7b742287e40e08 ^ 
I10323882c29157f609df5db826348e4bae6940d64129ac87b330976a2fe64027 ^ 
0; 



wire I8af4fe02e31ae2c79e572080447a2006f2c54deee1e3f370e18aa76d8e6e8009;
assign I8af4fe02e31ae2c79e572080447a2006f2c54deee1e3f370e18aa76d8e6e8009 = 
        y_nr_in[5] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
0; 



wire I74216e9a73872e99794068c277f9a181d4e3c30967bbea6a32379cc3e5e42abb;
assign I74216e9a73872e99794068c277f9a181d4e3c30967bbea6a32379cc3e5e42abb = 
        y_nr_in[47] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[68] = 
I8af4fe02e31ae2c79e572080447a2006f2c54deee1e3f370e18aa76d8e6e8009 ^ 
I74216e9a73872e99794068c277f9a181d4e3c30967bbea6a32379cc3e5e42abb ^ 
0; 



wire I517f12ae677e7d31fe721b16e3d659791b88c96a49f102fc4f8f784fab4e16cf;
assign I517f12ae677e7d31fe721b16e3d659791b88c96a49f102fc4f8f784fab4e16cf = 
        y_nr_in[6] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
0; 



wire I02d93a628f7ce5d2282b00d757b1c927103ecef65317e72750294857c4712f50;
assign I02d93a628f7ce5d2282b00d757b1c927103ecef65317e72750294857c4712f50 = 
        y_nr_in[44] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[69] = 
I517f12ae677e7d31fe721b16e3d659791b88c96a49f102fc4f8f784fab4e16cf ^ 
I02d93a628f7ce5d2282b00d757b1c927103ecef65317e72750294857c4712f50 ^ 
0; 



wire I5080b7960640e21fb77dc33352d27bf9decc8acbed5287cfa78f7c86f5185b67;
assign I5080b7960640e21fb77dc33352d27bf9decc8acbed5287cfa78f7c86f5185b67 = 
        y_nr_in[7] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
0; 



wire Ie0404d66f0866b036473b06f02ef982272d9132860b51fa17968331a2e608d22;
assign Ie0404d66f0866b036473b06f02ef982272d9132860b51fa17968331a2e608d22 = 
        y_nr_in[45] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[70] = 
I5080b7960640e21fb77dc33352d27bf9decc8acbed5287cfa78f7c86f5185b67 ^ 
Ie0404d66f0866b036473b06f02ef982272d9132860b51fa17968331a2e608d22 ^ 
0; 



wire I49252a481f98d44f48d620df37f7d2d75e8a81d0cfab91bb4eb7916b02e723f1;
assign I49252a481f98d44f48d620df37f7d2d75e8a81d0cfab91bb4eb7916b02e723f1 = 
        y_nr_in[4] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
0; 



wire I7e1e23d5c281dd756a4f0c0c90de3eb67b3f7d9d6bdf7350565d3e3f07fb40e9;
assign I7e1e23d5c281dd756a4f0c0c90de3eb67b3f7d9d6bdf7350565d3e3f07fb40e9 = 
        y_nr_in[46] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[71] = 
I49252a481f98d44f48d620df37f7d2d75e8a81d0cfab91bb4eb7916b02e723f1 ^ 
I7e1e23d5c281dd756a4f0c0c90de3eb67b3f7d9d6bdf7350565d3e3f07fb40e9 ^ 
0; 



wire I73435e48db187904fd803883a02dbb1dd75475a4acafef77a92b97309c741547;
assign I73435e48db187904fd803883a02dbb1dd75475a4acafef77a92b97309c741547 = 
        y_nr_in[2] ^ 
        y_nr_in[6] ^ 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[72] = 
I73435e48db187904fd803883a02dbb1dd75475a4acafef77a92b97309c741547 ^ 
0; 



wire Id591d53cae95d78d56e6790d8d48fdb1fccd924a3d74702da7da5906959360e3;
assign Id591d53cae95d78d56e6790d8d48fdb1fccd924a3d74702da7da5906959360e3 = 
        y_nr_in[3] ^ 
        y_nr_in[7] ^ 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[73] = 
Id591d53cae95d78d56e6790d8d48fdb1fccd924a3d74702da7da5906959360e3 ^ 
0; 



wire I713925d1fb7388f25956294817f33209972f03f18c8aacec62e323d73ce4d899;
assign I713925d1fb7388f25956294817f33209972f03f18c8aacec62e323d73ce4d899 = 
        y_nr_in[0] ^ 
        y_nr_in[4] ^ 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[74] = 
I713925d1fb7388f25956294817f33209972f03f18c8aacec62e323d73ce4d899 ^ 
0; 



wire I53dc58bcb983b221b7a34972e449bc96837c8331da3c4766e2b8f7dadfbe1df5;
assign I53dc58bcb983b221b7a34972e449bc96837c8331da3c4766e2b8f7dadfbe1df5 = 
        y_nr_in[1] ^ 
        y_nr_in[5] ^ 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[75] = 
I53dc58bcb983b221b7a34972e449bc96837c8331da3c4766e2b8f7dadfbe1df5 ^ 
0; 



wire I749df42857ecb08093aee2c6644a8d7ae85aacfbdd2223f385356c9c6d9debf2;
assign I749df42857ecb08093aee2c6644a8d7ae85aacfbdd2223f385356c9c6d9debf2 = 
        y_nr_in[7] ^ 
        y_nr_in[33] ^ 
        y_nr_in[41] ^ 
0; 



wire I87bfbcced728304ba648e08318be4a27aafbcb58f304a43b2179eaab05fd1da7;
assign I87bfbcced728304ba648e08318be4a27aafbcb58f304a43b2179eaab05fd1da7 = 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[76] = 
I749df42857ecb08093aee2c6644a8d7ae85aacfbdd2223f385356c9c6d9debf2 ^ 
I87bfbcced728304ba648e08318be4a27aafbcb58f304a43b2179eaab05fd1da7 ^ 
0; 



wire I4c5fd7f7ce5884fa78166d52d40761ae321ea77b9af18883e25457e5b8669979;
assign I4c5fd7f7ce5884fa78166d52d40761ae321ea77b9af18883e25457e5b8669979 = 
        y_nr_in[4] ^ 
        y_nr_in[34] ^ 
        y_nr_in[42] ^ 
0; 



wire I88f4b0ab82a5eda15c8279f1ab38fbf080d8eb2683e4c902f21ae9aa87cbb0b4;
assign I88f4b0ab82a5eda15c8279f1ab38fbf080d8eb2683e4c902f21ae9aa87cbb0b4 = 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[77] = 
I4c5fd7f7ce5884fa78166d52d40761ae321ea77b9af18883e25457e5b8669979 ^ 
I88f4b0ab82a5eda15c8279f1ab38fbf080d8eb2683e4c902f21ae9aa87cbb0b4 ^ 
0; 



wire I6eb66d4ad80b754c798d8c65f508f306cb534e3e6f249c4b0fa2ee249edd48b4;
assign I6eb66d4ad80b754c798d8c65f508f306cb534e3e6f249c4b0fa2ee249edd48b4 = 
        y_nr_in[5] ^ 
        y_nr_in[35] ^ 
        y_nr_in[43] ^ 
0; 



wire Ief6c16e2213875ba07e9778af61e6aa712e9f090115e50b808aaf555a9d0faa3;
assign Ief6c16e2213875ba07e9778af61e6aa712e9f090115e50b808aaf555a9d0faa3 = 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[78] = 
I6eb66d4ad80b754c798d8c65f508f306cb534e3e6f249c4b0fa2ee249edd48b4 ^ 
Ief6c16e2213875ba07e9778af61e6aa712e9f090115e50b808aaf555a9d0faa3 ^ 
0; 



wire I34b0ed27c72aebdc29f3e3cc6a170d2b86346de7b312ffebc3590537e8c36dda;
assign I34b0ed27c72aebdc29f3e3cc6a170d2b86346de7b312ffebc3590537e8c36dda = 
        y_nr_in[6] ^ 
        y_nr_in[32] ^ 
        y_nr_in[40] ^ 
0; 



wire I2e8db43d753a8065090cee7e4c38937040521dad8913bcea1ee83ddb7c261263;
assign I2e8db43d753a8065090cee7e4c38937040521dad8913bcea1ee83ddb7c261263 = 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[79] = 
I34b0ed27c72aebdc29f3e3cc6a170d2b86346de7b312ffebc3590537e8c36dda ^ 
I2e8db43d753a8065090cee7e4c38937040521dad8913bcea1ee83ddb7c261263 ^ 
0; 



wire Ie24702beb392c5cd6079ed852052c54b3c86e2f10600e0dca3b8da0b62173a37;
assign Ie24702beb392c5cd6079ed852052c54b3c86e2f10600e0dca3b8da0b62173a37 = 
        y_nr_in[3] ^ 
        y_nr_in[5] ^ 
        y_nr_in[24] ^ 
0; 



wire I29a049af74c07786f814c55fd562d3ae21f89db660bfeeab49e8465d8d6adce2;
assign I29a049af74c07786f814c55fd562d3ae21f89db660bfeeab49e8465d8d6adce2 = 
        y_nr_in[29] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[80] = 
Ie24702beb392c5cd6079ed852052c54b3c86e2f10600e0dca3b8da0b62173a37 ^ 
I29a049af74c07786f814c55fd562d3ae21f89db660bfeeab49e8465d8d6adce2 ^ 
0; 



wire I3588f0f60c6328afd0bfe1581a303b8f31e2ae540c44f66b3d384abaa24adfa1;
assign I3588f0f60c6328afd0bfe1581a303b8f31e2ae540c44f66b3d384abaa24adfa1 = 
        y_nr_in[0] ^ 
        y_nr_in[6] ^ 
        y_nr_in[25] ^ 
0; 



wire I68dcb1be9f7ffb526fb93d6151542e5147a2e48aa913d24a278324b0239734e8;
assign I68dcb1be9f7ffb526fb93d6151542e5147a2e48aa913d24a278324b0239734e8 = 
        y_nr_in[30] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[81] = 
I3588f0f60c6328afd0bfe1581a303b8f31e2ae540c44f66b3d384abaa24adfa1 ^ 
I68dcb1be9f7ffb526fb93d6151542e5147a2e48aa913d24a278324b0239734e8 ^ 
0; 



wire I8508ddaab52430f316f9f16f378014ffc6a953fc4c4925dc22b3f01fab1e04ec;
assign I8508ddaab52430f316f9f16f378014ffc6a953fc4c4925dc22b3f01fab1e04ec = 
        y_nr_in[1] ^ 
        y_nr_in[7] ^ 
        y_nr_in[26] ^ 
0; 



wire I9547f6e0fbd79d0314d3c2eca2c1f156b8df82742647263e4a58b3576c52abb2;
assign I9547f6e0fbd79d0314d3c2eca2c1f156b8df82742647263e4a58b3576c52abb2 = 
        y_nr_in[31] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[82] = 
I8508ddaab52430f316f9f16f378014ffc6a953fc4c4925dc22b3f01fab1e04ec ^ 
I9547f6e0fbd79d0314d3c2eca2c1f156b8df82742647263e4a58b3576c52abb2 ^ 
0; 



wire Id67bcba60edfed75aaccd2da1f874ebc0f9f0724c9e4e6eb7de598640c2fd1ee;
assign Id67bcba60edfed75aaccd2da1f874ebc0f9f0724c9e4e6eb7de598640c2fd1ee = 
        y_nr_in[2] ^ 
        y_nr_in[4] ^ 
        y_nr_in[27] ^ 
0; 



wire Id5899e25d911565cccda3cf9d743585ebe31d67293c58da28d009521882ff970;
assign Id5899e25d911565cccda3cf9d743585ebe31d67293c58da28d009521882ff970 = 
        y_nr_in[28] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[83] = 
Id67bcba60edfed75aaccd2da1f874ebc0f9f0724c9e4e6eb7de598640c2fd1ee ^ 
Id5899e25d911565cccda3cf9d743585ebe31d67293c58da28d009521882ff970 ^ 
0; 



wire I47715d5589693a211add4325635d4f400f10ff3764c88053c43945b8987786a0;
assign I47715d5589693a211add4325635d4f400f10ff3764c88053c43945b8987786a0 = 
        y_nr_in[3] ^ 
        y_nr_in[28] ^ 
        y_nr_in[38] ^ 
0; 



wire I544b46255aeb64cb243890e282884a2bb6f6621d0b15da83d1011f70f575e7b4;
assign I544b46255aeb64cb243890e282884a2bb6f6621d0b15da83d1011f70f575e7b4 = 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[84] = 
I47715d5589693a211add4325635d4f400f10ff3764c88053c43945b8987786a0 ^ 
I544b46255aeb64cb243890e282884a2bb6f6621d0b15da83d1011f70f575e7b4 ^ 
0; 



wire Ie287803eacbc0f4a71a1a0ac982c3ee7fa386e67f8660465bb0753e8222a6eb0;
assign Ie287803eacbc0f4a71a1a0ac982c3ee7fa386e67f8660465bb0753e8222a6eb0 = 
        y_nr_in[0] ^ 
        y_nr_in[29] ^ 
        y_nr_in[39] ^ 
0; 



wire I465e4d2978d3ba72563a24d7a472e161978a4a0a32c68a7b743812921bf2b251;
assign I465e4d2978d3ba72563a24d7a472e161978a4a0a32c68a7b743812921bf2b251 = 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[85] = 
Ie287803eacbc0f4a71a1a0ac982c3ee7fa386e67f8660465bb0753e8222a6eb0 ^ 
I465e4d2978d3ba72563a24d7a472e161978a4a0a32c68a7b743812921bf2b251 ^ 
0; 



wire Iee6d3f0d039c72da19a800305f1b5ae80057a2366ab53fb37bcbbf6fe541da47;
assign Iee6d3f0d039c72da19a800305f1b5ae80057a2366ab53fb37bcbbf6fe541da47 = 
        y_nr_in[1] ^ 
        y_nr_in[30] ^ 
        y_nr_in[36] ^ 
0; 



wire I7ad296c1cd3e7cb14f68633c581941ca97ee647e3cee75abb2369c9ff502ce15;
assign I7ad296c1cd3e7cb14f68633c581941ca97ee647e3cee75abb2369c9ff502ce15 = 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[86] = 
Iee6d3f0d039c72da19a800305f1b5ae80057a2366ab53fb37bcbbf6fe541da47 ^ 
I7ad296c1cd3e7cb14f68633c581941ca97ee647e3cee75abb2369c9ff502ce15 ^ 
0; 



wire I3493fe8f496c669528edad1b2638d9849cd91fe9aaad26300f8fed57aa5af16b;
assign I3493fe8f496c669528edad1b2638d9849cd91fe9aaad26300f8fed57aa5af16b = 
        y_nr_in[2] ^ 
        y_nr_in[31] ^ 
        y_nr_in[37] ^ 
0; 



wire Id870b3bfde35f3c9874846f92d335fbec810153d4af2b08a7cb41adc5d8cf82b;
assign Id870b3bfde35f3c9874846f92d335fbec810153d4af2b08a7cb41adc5d8cf82b = 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[87] = 
I3493fe8f496c669528edad1b2638d9849cd91fe9aaad26300f8fed57aa5af16b ^ 
Id870b3bfde35f3c9874846f92d335fbec810153d4af2b08a7cb41adc5d8cf82b ^ 
0; 



wire Icd8eb0102066b27b8a486a88894c9df50f922063098ef993825f3ac1b4924686;
assign Icd8eb0102066b27b8a486a88894c9df50f922063098ef993825f3ac1b4924686 = 
        y_nr_in[7] ^ 
        y_nr_in[15] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[88] = 
Icd8eb0102066b27b8a486a88894c9df50f922063098ef993825f3ac1b4924686 ^ 
0; 



wire If40b9c212bd0e0de6f44f266a1bdc600f3aacc50aa5bde4a4d88f3edd1bf545c;
assign If40b9c212bd0e0de6f44f266a1bdc600f3aacc50aa5bde4a4d88f3edd1bf545c = 
        y_nr_in[4] ^ 
        y_nr_in[12] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[89] = 
If40b9c212bd0e0de6f44f266a1bdc600f3aacc50aa5bde4a4d88f3edd1bf545c ^ 
0; 



wire Ia864fdd01430b3da092a9470cf806a86a8c8a8af5ea75238dde57eb4dc0152dc;
assign Ia864fdd01430b3da092a9470cf806a86a8c8a8af5ea75238dde57eb4dc0152dc = 
        y_nr_in[5] ^ 
        y_nr_in[13] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[90] = 
Ia864fdd01430b3da092a9470cf806a86a8c8a8af5ea75238dde57eb4dc0152dc ^ 
0; 



wire Ib27dc99958ae9b7eb461d6d0c638490563f842df99914da2d3b080bdd6ca8cf4;
assign Ib27dc99958ae9b7eb461d6d0c638490563f842df99914da2d3b080bdd6ca8cf4 = 
        y_nr_in[6] ^ 
        y_nr_in[14] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[91] = 
Ib27dc99958ae9b7eb461d6d0c638490563f842df99914da2d3b080bdd6ca8cf4 ^ 
0; 



wire Ic3a6500f0db687d0d51af6fbdb08f18912f269e77726fdfa48dd416825b289f9;
assign Ic3a6500f0db687d0d51af6fbdb08f18912f269e77726fdfa48dd416825b289f9 = 
        y_nr_in[3] ^ 
        y_nr_in[6] ^ 
        y_nr_in[34] ^ 
0; 



wire I0a0bdc1f0ad53c82619129048bc4767c5943fa126303e1c2732a4011206368ce;
assign I0a0bdc1f0ad53c82619129048bc4767c5943fa126303e1c2732a4011206368ce = 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[92] = 
Ic3a6500f0db687d0d51af6fbdb08f18912f269e77726fdfa48dd416825b289f9 ^ 
I0a0bdc1f0ad53c82619129048bc4767c5943fa126303e1c2732a4011206368ce ^ 
0; 



wire I856ef2bb3dc89e261fcfd023d50ce1779036a51c8abccb8eff03feadeb2136c1;
assign I856ef2bb3dc89e261fcfd023d50ce1779036a51c8abccb8eff03feadeb2136c1 = 
        y_nr_in[0] ^ 
        y_nr_in[7] ^ 
        y_nr_in[35] ^ 
0; 



wire Ic19fde74f844e3c149ea45163c5a367e003533a9102eedf1d1c94a74c3fb736c;
assign Ic19fde74f844e3c149ea45163c5a367e003533a9102eedf1d1c94a74c3fb736c = 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[93] = 
I856ef2bb3dc89e261fcfd023d50ce1779036a51c8abccb8eff03feadeb2136c1 ^ 
Ic19fde74f844e3c149ea45163c5a367e003533a9102eedf1d1c94a74c3fb736c ^ 
0; 



wire I17884245955f22f700a4465acc6df8ea9a629629dbfa7317da5b1639d55d1328;
assign I17884245955f22f700a4465acc6df8ea9a629629dbfa7317da5b1639d55d1328 = 
        y_nr_in[1] ^ 
        y_nr_in[4] ^ 
        y_nr_in[32] ^ 
0; 



wire If8dbbb14e8187550ba2a78d2ca0ddffdb0652e4a4534e941814f24847a4ab1ab;
assign If8dbbb14e8187550ba2a78d2ca0ddffdb0652e4a4534e941814f24847a4ab1ab = 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[94] = 
I17884245955f22f700a4465acc6df8ea9a629629dbfa7317da5b1639d55d1328 ^ 
If8dbbb14e8187550ba2a78d2ca0ddffdb0652e4a4534e941814f24847a4ab1ab ^ 
0; 



wire Ie2b96c7554f57d93f81837f59c7f9a2c8f6cb907e2338b0c70294da7d0127afb;
assign Ie2b96c7554f57d93f81837f59c7f9a2c8f6cb907e2338b0c70294da7d0127afb = 
        y_nr_in[2] ^ 
        y_nr_in[5] ^ 
        y_nr_in[33] ^ 
0; 



wire Idafc600229f800e83c3212c1ebe290da56790a4899c881856b03c609c885f60c;
assign Idafc600229f800e83c3212c1ebe290da56790a4899c881856b03c609c885f60c = 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[95] = 
Ie2b96c7554f57d93f81837f59c7f9a2c8f6cb907e2338b0c70294da7d0127afb ^ 
Idafc600229f800e83c3212c1ebe290da56790a4899c881856b03c609c885f60c ^ 
0; 



wire I91641d702f8e03b4ac11a95d171c335003dc9432f89e8c5b2de0b1a15af20f83;
assign I91641d702f8e03b4ac11a95d171c335003dc9432f89e8c5b2de0b1a15af20f83 = 
        y_nr_in[7] ^ 
        y_nr_in[25] ^ 
        y_nr_in[47] ^ 
0; 



wire Ifc3aef378b28c216a4af8fb5f7dcdf89cf548b2e36f0bf0c77ad0b11d82eddce;
assign Ifc3aef378b28c216a4af8fb5f7dcdf89cf548b2e36f0bf0c77ad0b11d82eddce = 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[96] = 
I91641d702f8e03b4ac11a95d171c335003dc9432f89e8c5b2de0b1a15af20f83 ^ 
Ifc3aef378b28c216a4af8fb5f7dcdf89cf548b2e36f0bf0c77ad0b11d82eddce ^ 
0; 



wire I6e417d3a471a9e0d9f5d49dea659fcf95546c65bf8a89b4ff8236b99e60f164f;
assign I6e417d3a471a9e0d9f5d49dea659fcf95546c65bf8a89b4ff8236b99e60f164f = 
        y_nr_in[4] ^ 
        y_nr_in[26] ^ 
        y_nr_in[44] ^ 
0; 



wire I491c60a528bfdd4cb94bf33383eeef5c85a5278bac31ed0f7b506350ac7f36f9;
assign I491c60a528bfdd4cb94bf33383eeef5c85a5278bac31ed0f7b506350ac7f36f9 = 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[97] = 
I6e417d3a471a9e0d9f5d49dea659fcf95546c65bf8a89b4ff8236b99e60f164f ^ 
I491c60a528bfdd4cb94bf33383eeef5c85a5278bac31ed0f7b506350ac7f36f9 ^ 
0; 



wire I6a680c4155beebef7694e7ee0792fae3bda79332e666cf11255339a2c8d7058b;
assign I6a680c4155beebef7694e7ee0792fae3bda79332e666cf11255339a2c8d7058b = 
        y_nr_in[5] ^ 
        y_nr_in[27] ^ 
        y_nr_in[45] ^ 
0; 



wire Ib069571649c5c887e2cbd7a4d0338ab559f7c4dd886046a2d09167a46334c555;
assign Ib069571649c5c887e2cbd7a4d0338ab559f7c4dd886046a2d09167a46334c555 = 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[98] = 
I6a680c4155beebef7694e7ee0792fae3bda79332e666cf11255339a2c8d7058b ^ 
Ib069571649c5c887e2cbd7a4d0338ab559f7c4dd886046a2d09167a46334c555 ^ 
0; 



wire Ic815e6831394d6bd3233a3e4459d1bf98d212c4e76047397ea19d092b25e36df;
assign Ic815e6831394d6bd3233a3e4459d1bf98d212c4e76047397ea19d092b25e36df = 
        y_nr_in[6] ^ 
        y_nr_in[24] ^ 
        y_nr_in[46] ^ 
0; 



wire I187ae6c92c5db73f13c20c8c99a5d179a56b9cb61b478de1310032a0fd4ff666;
assign I187ae6c92c5db73f13c20c8c99a5d179a56b9cb61b478de1310032a0fd4ff666 = 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[99] = 
Ic815e6831394d6bd3233a3e4459d1bf98d212c4e76047397ea19d092b25e36df ^ 
I187ae6c92c5db73f13c20c8c99a5d179a56b9cb61b478de1310032a0fd4ff666 ^ 
0; 



wire Ice55a85f2415b4c7279ede14afed095c630a5bc515e04d114b4b0d51cd3799d6;
assign Ice55a85f2415b4c7279ede14afed095c630a5bc515e04d114b4b0d51cd3799d6 = 
        y_nr_in[3] ^ 
        y_nr_in[43] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[100] = 
Ice55a85f2415b4c7279ede14afed095c630a5bc515e04d114b4b0d51cd3799d6 ^ 
0; 



wire Ide2a61371c25d75c6fe8b6f961d9d61ffa5a571c624df6eca6606b9ec20d1bba;
assign Ide2a61371c25d75c6fe8b6f961d9d61ffa5a571c624df6eca6606b9ec20d1bba = 
        y_nr_in[0] ^ 
        y_nr_in[40] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[101] = 
Ide2a61371c25d75c6fe8b6f961d9d61ffa5a571c624df6eca6606b9ec20d1bba ^ 
0; 



wire I57c8dc6535a07e9500c1d69fb47ae667fe2f17d2582a74d8353a783a62c45a8a;
assign I57c8dc6535a07e9500c1d69fb47ae667fe2f17d2582a74d8353a783a62c45a8a = 
        y_nr_in[1] ^ 
        y_nr_in[41] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[102] = 
I57c8dc6535a07e9500c1d69fb47ae667fe2f17d2582a74d8353a783a62c45a8a ^ 
0; 



wire Ie0f8f4f7109da8084b2b8eca4bc4215906cfc7e6edd880b1aa29939559202701;
assign Ie0f8f4f7109da8084b2b8eca4bc4215906cfc7e6edd880b1aa29939559202701 = 
        y_nr_in[2] ^ 
        y_nr_in[42] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[103] = 
Ie0f8f4f7109da8084b2b8eca4bc4215906cfc7e6edd880b1aa29939559202701 ^ 
0; 



wire Ibc45c4ef0bbb3d113baea1e18c7f8d3f6f96e321f2ab4ebe81f846bf69777242;
assign Ibc45c4ef0bbb3d113baea1e18c7f8d3f6f96e321f2ab4ebe81f846bf69777242 = 
        y_nr_in[7] ^ 
        y_nr_in[38] ^ 
        y_nr_in[44] ^ 
0; 



wire I3f01361b7c4ce8ebd96c22ab1453db87d96e7f873603c7b30d56ca47f13b6714;
assign I3f01361b7c4ce8ebd96c22ab1453db87d96e7f873603c7b30d56ca47f13b6714 = 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[104] = 
Ibc45c4ef0bbb3d113baea1e18c7f8d3f6f96e321f2ab4ebe81f846bf69777242 ^ 
I3f01361b7c4ce8ebd96c22ab1453db87d96e7f873603c7b30d56ca47f13b6714 ^ 
0; 



wire Ibbe4b59beb321340409af03246b06a8e9a4d456aa02b0997ebc46f152fa802a8;
assign Ibbe4b59beb321340409af03246b06a8e9a4d456aa02b0997ebc46f152fa802a8 = 
        y_nr_in[4] ^ 
        y_nr_in[39] ^ 
        y_nr_in[45] ^ 
0; 



wire I162055d6ef485b5e4b0dbb94462101188b37208dabd17dc96a39c06f6b30a8e4;
assign I162055d6ef485b5e4b0dbb94462101188b37208dabd17dc96a39c06f6b30a8e4 = 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[105] = 
Ibbe4b59beb321340409af03246b06a8e9a4d456aa02b0997ebc46f152fa802a8 ^ 
I162055d6ef485b5e4b0dbb94462101188b37208dabd17dc96a39c06f6b30a8e4 ^ 
0; 



wire I9b1e08a0ca00dc7e8f7daf895fda5497cbe70eaa656ac4ff277551e97018fefb;
assign I9b1e08a0ca00dc7e8f7daf895fda5497cbe70eaa656ac4ff277551e97018fefb = 
        y_nr_in[5] ^ 
        y_nr_in[36] ^ 
        y_nr_in[46] ^ 
0; 



wire I587dfa066c058e19f7f8df7e189a414e9fe2272f17dcc1dbc23cfc32c5f368e4;
assign I587dfa066c058e19f7f8df7e189a414e9fe2272f17dcc1dbc23cfc32c5f368e4 = 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[106] = 
I9b1e08a0ca00dc7e8f7daf895fda5497cbe70eaa656ac4ff277551e97018fefb ^ 
I587dfa066c058e19f7f8df7e189a414e9fe2272f17dcc1dbc23cfc32c5f368e4 ^ 
0; 



wire I460fa50de867246cdbafbb2ed7c1ecd55ded8d3aedcfdb817d6ccf8db5871d23;
assign I460fa50de867246cdbafbb2ed7c1ecd55ded8d3aedcfdb817d6ccf8db5871d23 = 
        y_nr_in[6] ^ 
        y_nr_in[37] ^ 
        y_nr_in[47] ^ 
0; 



wire Ie72c6bbd4f0254c15d6fa7bea2c562a9c5ac7b7266b19ba472e7e90d53ac3cc9;
assign Ie72c6bbd4f0254c15d6fa7bea2c562a9c5ac7b7266b19ba472e7e90d53ac3cc9 = 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[107] = 
I460fa50de867246cdbafbb2ed7c1ecd55ded8d3aedcfdb817d6ccf8db5871d23 ^ 
Ie72c6bbd4f0254c15d6fa7bea2c562a9c5ac7b7266b19ba472e7e90d53ac3cc9 ^ 
0; 



wire Icdf9ac94d836cad93dfa839c9a62b7e868031f7668df7c94ef1697e802dcc877;
assign Icdf9ac94d836cad93dfa839c9a62b7e868031f7668df7c94ef1697e802dcc877 = 
        y_nr_in[6] ^ 
        y_nr_in[20] ^ 
        y_nr_in[46] ^ 
0; 



wire I61fd8679995a76dfae8612070cc2f5076c5f927d6a74c74e20594c0204e582a8;
assign I61fd8679995a76dfae8612070cc2f5076c5f927d6a74c74e20594c0204e582a8 = 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[108] = 
Icdf9ac94d836cad93dfa839c9a62b7e868031f7668df7c94ef1697e802dcc877 ^ 
I61fd8679995a76dfae8612070cc2f5076c5f927d6a74c74e20594c0204e582a8 ^ 
0; 



wire I0e482967ea7d57374d6f59e40de6353c393a3d4a2a00d2ba78e8771b2fc70c49;
assign I0e482967ea7d57374d6f59e40de6353c393a3d4a2a00d2ba78e8771b2fc70c49 = 
        y_nr_in[7] ^ 
        y_nr_in[21] ^ 
        y_nr_in[47] ^ 
0; 



wire I1d2c7f473b80536c78739cb61fe4b82f212f19bf96e30a8c767456f7395e5b57;
assign I1d2c7f473b80536c78739cb61fe4b82f212f19bf96e30a8c767456f7395e5b57 = 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[109] = 
I0e482967ea7d57374d6f59e40de6353c393a3d4a2a00d2ba78e8771b2fc70c49 ^ 
I1d2c7f473b80536c78739cb61fe4b82f212f19bf96e30a8c767456f7395e5b57 ^ 
0; 



wire I568ed6b5eb066fb08f700df101440b08ab685ae80d50bbe9001d0631786bb568;
assign I568ed6b5eb066fb08f700df101440b08ab685ae80d50bbe9001d0631786bb568 = 
        y_nr_in[4] ^ 
        y_nr_in[22] ^ 
        y_nr_in[44] ^ 
0; 



wire I6526732e56e3f5dcd1535b6ecb28529241fe7a4f5edfc8e98552d7809b71a2f3;
assign I6526732e56e3f5dcd1535b6ecb28529241fe7a4f5edfc8e98552d7809b71a2f3 = 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[110] = 
I568ed6b5eb066fb08f700df101440b08ab685ae80d50bbe9001d0631786bb568 ^ 
I6526732e56e3f5dcd1535b6ecb28529241fe7a4f5edfc8e98552d7809b71a2f3 ^ 
0; 



wire Idf28e7e65f6083f41b0e07b8e973799209c760d5847f4455789ca23d090e95a4;
assign Idf28e7e65f6083f41b0e07b8e973799209c760d5847f4455789ca23d090e95a4 = 
        y_nr_in[5] ^ 
        y_nr_in[23] ^ 
        y_nr_in[45] ^ 
0; 



wire If137b1c6ddff5cbc91b835e9e6a58bf730fe508bf743278acc77bcfc08055740;
assign If137b1c6ddff5cbc91b835e9e6a58bf730fe508bf743278acc77bcfc08055740 = 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[111] = 
Idf28e7e65f6083f41b0e07b8e973799209c760d5847f4455789ca23d090e95a4 ^ 
If137b1c6ddff5cbc91b835e9e6a58bf730fe508bf743278acc77bcfc08055740 ^ 
0; 



wire I11a3fb05b63d83c01200575b62acae3aadc314ce9aab3cfc712ad953e8c6be0d;
assign I11a3fb05b63d83c01200575b62acae3aadc314ce9aab3cfc712ad953e8c6be0d = 
        y_nr_in[0] ^ 
        y_nr_in[26] ^ 
        y_nr_in[30] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[112] = 
I11a3fb05b63d83c01200575b62acae3aadc314ce9aab3cfc712ad953e8c6be0d ^ 
0; 



wire If4b9e7140e7d54fc9a5edf7419466cc3b1ffafae193e57955ab6ba0126935612;
assign If4b9e7140e7d54fc9a5edf7419466cc3b1ffafae193e57955ab6ba0126935612 = 
        y_nr_in[1] ^ 
        y_nr_in[27] ^ 
        y_nr_in[31] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[113] = 
If4b9e7140e7d54fc9a5edf7419466cc3b1ffafae193e57955ab6ba0126935612 ^ 
0; 



wire I8270680f0bdef107e425e370941e7551c61b94445426e1d05ae82ebccd640a31;
assign I8270680f0bdef107e425e370941e7551c61b94445426e1d05ae82ebccd640a31 = 
        y_nr_in[2] ^ 
        y_nr_in[24] ^ 
        y_nr_in[28] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[114] = 
I8270680f0bdef107e425e370941e7551c61b94445426e1d05ae82ebccd640a31 ^ 
0; 



wire I0e74277dc013daff01c991b662f603636c49561ddcdcce2a615c6e436223375e;
assign I0e74277dc013daff01c991b662f603636c49561ddcdcce2a615c6e436223375e = 
        y_nr_in[3] ^ 
        y_nr_in[25] ^ 
        y_nr_in[29] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[115] = 
I0e74277dc013daff01c991b662f603636c49561ddcdcce2a615c6e436223375e ^ 
0; 



wire If9954bea361542b75caef106626c8c70a82af99e72e42bb3ef82bcdce6812c14;
assign If9954bea361542b75caef106626c8c70a82af99e72e42bb3ef82bcdce6812c14 = 
        y_nr_in[3] ^ 
        y_nr_in[4] ^ 
        y_nr_in[41] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[116] = 
If9954bea361542b75caef106626c8c70a82af99e72e42bb3ef82bcdce6812c14 ^ 
0; 



wire I828edcf234bef402fe2316bb47470ed601da0d7c8873c5a08924ed7d7b8acc13;
assign I828edcf234bef402fe2316bb47470ed601da0d7c8873c5a08924ed7d7b8acc13 = 
        y_nr_in[0] ^ 
        y_nr_in[5] ^ 
        y_nr_in[42] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[117] = 
I828edcf234bef402fe2316bb47470ed601da0d7c8873c5a08924ed7d7b8acc13 ^ 
0; 



wire I0016f92178cc6d08a0bf61e8ace71cb46a555e6d5691390e2e8d68f36cf884f1;
assign I0016f92178cc6d08a0bf61e8ace71cb46a555e6d5691390e2e8d68f36cf884f1 = 
        y_nr_in[1] ^ 
        y_nr_in[6] ^ 
        y_nr_in[43] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[118] = 
I0016f92178cc6d08a0bf61e8ace71cb46a555e6d5691390e2e8d68f36cf884f1 ^ 
0; 



wire I6f6357d36e2e7908a0040f12e0e72e8fbee173fa530262abf4fd5ca4d98f4668;
assign I6f6357d36e2e7908a0040f12e0e72e8fbee173fa530262abf4fd5ca4d98f4668 = 
        y_nr_in[2] ^ 
        y_nr_in[7] ^ 
        y_nr_in[40] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[119] = 
I6f6357d36e2e7908a0040f12e0e72e8fbee173fa530262abf4fd5ca4d98f4668 ^ 
0; 



wire I73018bcf124b97c0bc6e72cd6ea93dbfa91414b23010be5b621483f62f3a4578;
assign I73018bcf124b97c0bc6e72cd6ea93dbfa91414b23010be5b621483f62f3a4578 = 
        y_nr_in[6] ^ 
        y_nr_in[17] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[120] = 
I73018bcf124b97c0bc6e72cd6ea93dbfa91414b23010be5b621483f62f3a4578 ^ 
0; 



wire I198acfe9869520864d1e204df0f6f9c2de50b8e2d495153b89eed1618a9aa245;
assign I198acfe9869520864d1e204df0f6f9c2de50b8e2d495153b89eed1618a9aa245 = 
        y_nr_in[7] ^ 
        y_nr_in[18] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[121] = 
I198acfe9869520864d1e204df0f6f9c2de50b8e2d495153b89eed1618a9aa245 ^ 
0; 



wire Ie3eb10e9c58d1d3a6b6508f0e4e6f01474249cb13ffb479b1f5413308fb904d5;
assign Ie3eb10e9c58d1d3a6b6508f0e4e6f01474249cb13ffb479b1f5413308fb904d5 = 
        y_nr_in[4] ^ 
        y_nr_in[19] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[122] = 
Ie3eb10e9c58d1d3a6b6508f0e4e6f01474249cb13ffb479b1f5413308fb904d5 ^ 
0; 



wire I8a013efc26787c6ce8f85e42c73d78841020ba2c76844a4dae33aeece25c5357;
assign I8a013efc26787c6ce8f85e42c73d78841020ba2c76844a4dae33aeece25c5357 = 
        y_nr_in[5] ^ 
        y_nr_in[16] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[123] = 
I8a013efc26787c6ce8f85e42c73d78841020ba2c76844a4dae33aeece25c5357 ^ 
0; 



wire I09dd53def80e325c7ea5c3c8e2f064b02ebfe59c3b761e79a215a689b5e7cc40;
assign I09dd53def80e325c7ea5c3c8e2f064b02ebfe59c3b761e79a215a689b5e7cc40 = 
        y_nr_in[0] ^ 
        y_nr_in[34] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[124] = 
I09dd53def80e325c7ea5c3c8e2f064b02ebfe59c3b761e79a215a689b5e7cc40 ^ 
0; 



wire Icb2b0bd16431524939cdded20f245161f930c9c47942f8120e64560b9bc36d7b;
assign Icb2b0bd16431524939cdded20f245161f930c9c47942f8120e64560b9bc36d7b = 
        y_nr_in[1] ^ 
        y_nr_in[35] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[125] = 
Icb2b0bd16431524939cdded20f245161f930c9c47942f8120e64560b9bc36d7b ^ 
0; 



wire I6ae1ea820cf145f6e4643d41e39249c25380a19ccaa261f4cb5bc84ca04d1269;
assign I6ae1ea820cf145f6e4643d41e39249c25380a19ccaa261f4cb5bc84ca04d1269 = 
        y_nr_in[2] ^ 
        y_nr_in[32] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[126] = 
I6ae1ea820cf145f6e4643d41e39249c25380a19ccaa261f4cb5bc84ca04d1269 ^ 
0; 



wire I0e0ac64caea92a1d75ed5a9ff960681180e0d9a0b5a7e7522163cd406b908016;
assign I0e0ac64caea92a1d75ed5a9ff960681180e0d9a0b5a7e7522163cd406b908016 = 
        y_nr_in[3] ^ 
        y_nr_in[33] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[127] = 
I0e0ac64caea92a1d75ed5a9ff960681180e0d9a0b5a7e7522163cd406b908016 ^ 
0; 



wire I04e612eeeb21a866edeba1827f31fa3cfc5da5103261c5ff87c84c10b29e377d;
assign I04e612eeeb21a866edeba1827f31fa3cfc5da5103261c5ff87c84c10b29e377d = 
        y_nr_in[6] ^ 
        y_nr_in[11] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[128] = 
I04e612eeeb21a866edeba1827f31fa3cfc5da5103261c5ff87c84c10b29e377d ^ 
0; 



wire Iee83a9c6af510d609d531cafcc69628ca25af630d1b1c423885d4bbac737161f;
assign Iee83a9c6af510d609d531cafcc69628ca25af630d1b1c423885d4bbac737161f = 
        y_nr_in[7] ^ 
        y_nr_in[8] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[129] = 
Iee83a9c6af510d609d531cafcc69628ca25af630d1b1c423885d4bbac737161f ^ 
0; 



wire Ifdeff48f8f63ae1b707c6d44f01b027e2fb439655b8f09b37027edd781ee975e;
assign Ifdeff48f8f63ae1b707c6d44f01b027e2fb439655b8f09b37027edd781ee975e = 
        y_nr_in[4] ^ 
        y_nr_in[9] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[130] = 
Ifdeff48f8f63ae1b707c6d44f01b027e2fb439655b8f09b37027edd781ee975e ^ 
0; 



wire I54b1cfe31e5bd3dbbd4fa7c0e7800e1690c59de900c6dc0fe6045bff598d6972;
assign I54b1cfe31e5bd3dbbd4fa7c0e7800e1690c59de900c6dc0fe6045bff598d6972 = 
        y_nr_in[5] ^ 
        y_nr_in[10] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[131] = 
I54b1cfe31e5bd3dbbd4fa7c0e7800e1690c59de900c6dc0fe6045bff598d6972 ^ 
0; 



wire I0808f3f511663abe7288885dd511c482c1b6b7f8bff3b15b4a791e9004c78b75;
assign I0808f3f511663abe7288885dd511c482c1b6b7f8bff3b15b4a791e9004c78b75 = 
        y_nr_in[3] ^ 
        y_nr_in[15] ^ 
        y_nr_in[22] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[132] = 
I0808f3f511663abe7288885dd511c482c1b6b7f8bff3b15b4a791e9004c78b75 ^ 
0; 



wire I6b6989abe368b02139bf779aa6bd0ea63a67a493bf3a170d2fe37b0f62462b7b;
assign I6b6989abe368b02139bf779aa6bd0ea63a67a493bf3a170d2fe37b0f62462b7b = 
        y_nr_in[0] ^ 
        y_nr_in[12] ^ 
        y_nr_in[23] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[133] = 
I6b6989abe368b02139bf779aa6bd0ea63a67a493bf3a170d2fe37b0f62462b7b ^ 
0; 



wire I8723d833aaa6375f50399022729689f26a214a6d3386577cbe76e43bfaead2f9;
assign I8723d833aaa6375f50399022729689f26a214a6d3386577cbe76e43bfaead2f9 = 
        y_nr_in[1] ^ 
        y_nr_in[13] ^ 
        y_nr_in[20] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[134] = 
I8723d833aaa6375f50399022729689f26a214a6d3386577cbe76e43bfaead2f9 ^ 
0; 



wire I9036d79d85649603ba008bee293e9a61721de8dfb3ea0c780caf8befb8c59da2;
assign I9036d79d85649603ba008bee293e9a61721de8dfb3ea0c780caf8befb8c59da2 = 
        y_nr_in[2] ^ 
        y_nr_in[14] ^ 
        y_nr_in[21] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[135] = 
I9036d79d85649603ba008bee293e9a61721de8dfb3ea0c780caf8befb8c59da2 ^ 
0; 



wire I68abd03f6b7e831232b1811637b67182a1547f4b49ce74bf3c64be5d8c92a353;
assign I68abd03f6b7e831232b1811637b67182a1547f4b49ce74bf3c64be5d8c92a353 = 
        y_nr_in[6] ^ 
        y_nr_in[11] ^ 
        y_nr_in[36] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[136] = 
I68abd03f6b7e831232b1811637b67182a1547f4b49ce74bf3c64be5d8c92a353 ^ 
0; 



wire I5a2c723ed8fd3c3a348a0c101a5dc19af4119ed12bf2e21b4a99534a0f4c685b;
assign I5a2c723ed8fd3c3a348a0c101a5dc19af4119ed12bf2e21b4a99534a0f4c685b = 
        y_nr_in[7] ^ 
        y_nr_in[8] ^ 
        y_nr_in[37] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[137] = 
I5a2c723ed8fd3c3a348a0c101a5dc19af4119ed12bf2e21b4a99534a0f4c685b ^ 
0; 



wire Ia304d4a11073812e03c60d974ce8263b191a6a8e0e607016cb97e203e1ce574c;
assign Ia304d4a11073812e03c60d974ce8263b191a6a8e0e607016cb97e203e1ce574c = 
        y_nr_in[4] ^ 
        y_nr_in[9] ^ 
        y_nr_in[38] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[138] = 
Ia304d4a11073812e03c60d974ce8263b191a6a8e0e607016cb97e203e1ce574c ^ 
0; 



wire If0fdcc606689de54b4d5c073b32361cd4e2dd18918d442f8ba79f91104fdb8d1;
assign If0fdcc606689de54b4d5c073b32361cd4e2dd18918d442f8ba79f91104fdb8d1 = 
        y_nr_in[5] ^ 
        y_nr_in[10] ^ 
        y_nr_in[39] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[139] = 
If0fdcc606689de54b4d5c073b32361cd4e2dd18918d442f8ba79f91104fdb8d1 ^ 
0; 



wire Ib76ac2efd49415c33cd7fcdf86117582203844469bef6fb1aa6f18900ca60a5c;
assign Ib76ac2efd49415c33cd7fcdf86117582203844469bef6fb1aa6f18900ca60a5c = 
        y_nr_in[0] ^ 
        y_nr_in[20] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[140] = 
Ib76ac2efd49415c33cd7fcdf86117582203844469bef6fb1aa6f18900ca60a5c ^ 
0; 



wire I92b68e093194b90a895bbcb5099de8d29c6794a60a577d4eed46d76e9b32c771;
assign I92b68e093194b90a895bbcb5099de8d29c6794a60a577d4eed46d76e9b32c771 = 
        y_nr_in[1] ^ 
        y_nr_in[21] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[141] = 
I92b68e093194b90a895bbcb5099de8d29c6794a60a577d4eed46d76e9b32c771 ^ 
0; 



wire Ieffbeb4c9fb0242ffc90388bc5d16c0c78b4062ddbdfbb930493030a31fbc952;
assign Ieffbeb4c9fb0242ffc90388bc5d16c0c78b4062ddbdfbb930493030a31fbc952 = 
        y_nr_in[2] ^ 
        y_nr_in[22] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[142] = 
Ieffbeb4c9fb0242ffc90388bc5d16c0c78b4062ddbdfbb930493030a31fbc952 ^ 
0; 



wire Icd559c515beaeb5e638188f70e32299ef43943b0ce1d19e80f29eba0679bee12;
assign Icd559c515beaeb5e638188f70e32299ef43943b0ce1d19e80f29eba0679bee12 = 
        y_nr_in[3] ^ 
        y_nr_in[23] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[143] = 
Icd559c515beaeb5e638188f70e32299ef43943b0ce1d19e80f29eba0679bee12 ^ 
0; 



wire Ie2e2b08e080a117ff65e7040ffa15e72db6c1310243629d972c7139b0f5a3c05;
assign Ie2e2b08e080a117ff65e7040ffa15e72db6c1310243629d972c7139b0f5a3c05 = 
        y_nr_in[9] ^ 
        y_nr_in[31] ^ 
        y_nr_in[48] ^ 
0; 



wire I684fc51d495fedfd9bdafe94485a2cd8688ee121e5c2978bab87f9fd4e37d80b;
assign I684fc51d495fedfd9bdafe94485a2cd8688ee121e5c2978bab87f9fd4e37d80b = 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[144] = 
Ie2e2b08e080a117ff65e7040ffa15e72db6c1310243629d972c7139b0f5a3c05 ^ 
I684fc51d495fedfd9bdafe94485a2cd8688ee121e5c2978bab87f9fd4e37d80b ^ 
0; 



wire Ie32b6bd5e13ab6e0255cfa736314da54c7eb2ed64454f351be4fc653cc73ad3d;
assign Ie32b6bd5e13ab6e0255cfa736314da54c7eb2ed64454f351be4fc653cc73ad3d = 
        y_nr_in[10] ^ 
        y_nr_in[28] ^ 
        y_nr_in[49] ^ 
0; 



wire If4991a5d7d21efa79dc59a917034abd85e727ca8e4d68922a3ba80b6dafeed93;
assign If4991a5d7d21efa79dc59a917034abd85e727ca8e4d68922a3ba80b6dafeed93 = 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[145] = 
Ie32b6bd5e13ab6e0255cfa736314da54c7eb2ed64454f351be4fc653cc73ad3d ^ 
If4991a5d7d21efa79dc59a917034abd85e727ca8e4d68922a3ba80b6dafeed93 ^ 
0; 



wire I4537c147914b240750383c57700b9c4687a349f441c6fda2c8ab80aa93ec8272;
assign I4537c147914b240750383c57700b9c4687a349f441c6fda2c8ab80aa93ec8272 = 
        y_nr_in[11] ^ 
        y_nr_in[29] ^ 
        y_nr_in[50] ^ 
0; 



wire Ic358968cbf334449efb91fe3a98a6228903c5c0bef6f2e81cfca8cd8735984d0;
assign Ic358968cbf334449efb91fe3a98a6228903c5c0bef6f2e81cfca8cd8735984d0 = 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[146] = 
I4537c147914b240750383c57700b9c4687a349f441c6fda2c8ab80aa93ec8272 ^ 
Ic358968cbf334449efb91fe3a98a6228903c5c0bef6f2e81cfca8cd8735984d0 ^ 
0; 



wire Ic80cfcf328cef7e9932b182f78996b4571cd505fce91f1bc6e1558c98751dc19;
assign Ic80cfcf328cef7e9932b182f78996b4571cd505fce91f1bc6e1558c98751dc19 = 
        y_nr_in[8] ^ 
        y_nr_in[30] ^ 
        y_nr_in[51] ^ 
0; 



wire Ib32fbf2ce5ebae1700f9ed1264dc6ccec4d49d411a6d0333aea050ce8139b610;
assign Ib32fbf2ce5ebae1700f9ed1264dc6ccec4d49d411a6d0333aea050ce8139b610 = 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[147] = 
Ic80cfcf328cef7e9932b182f78996b4571cd505fce91f1bc6e1558c98751dc19 ^ 
Ib32fbf2ce5ebae1700f9ed1264dc6ccec4d49d411a6d0333aea050ce8139b610 ^ 
0; 



wire I1e29ad7126c9994135a12ef7507fa4d7988055cc266445a55effbf6de0a0bf1a;
assign I1e29ad7126c9994135a12ef7507fa4d7988055cc266445a55effbf6de0a0bf1a = 
        y_nr_in[0] ^ 
        y_nr_in[27] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[148] = 
I1e29ad7126c9994135a12ef7507fa4d7988055cc266445a55effbf6de0a0bf1a ^ 
0; 



wire Idc56dcfa439c82ce544cec043fbb3f4b4ff644879ce68c071c6247ea236e1071;
assign Idc56dcfa439c82ce544cec043fbb3f4b4ff644879ce68c071c6247ea236e1071 = 
        y_nr_in[1] ^ 
        y_nr_in[24] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[149] = 
Idc56dcfa439c82ce544cec043fbb3f4b4ff644879ce68c071c6247ea236e1071 ^ 
0; 



wire Ifa3c0791921cff838fa1d35eed6744fd64727fc362c31d54baa6fc3d8cff13d2;
assign Ifa3c0791921cff838fa1d35eed6744fd64727fc362c31d54baa6fc3d8cff13d2 = 
        y_nr_in[2] ^ 
        y_nr_in[25] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[150] = 
Ifa3c0791921cff838fa1d35eed6744fd64727fc362c31d54baa6fc3d8cff13d2 ^ 
0; 



wire Ica3e70c51fbbb23af567352e4d10f1931a92bbfe1e3ea9d9888a9fd29b207813;
assign Ica3e70c51fbbb23af567352e4d10f1931a92bbfe1e3ea9d9888a9fd29b207813 = 
        y_nr_in[3] ^ 
        y_nr_in[26] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[151] = 
Ica3e70c51fbbb23af567352e4d10f1931a92bbfe1e3ea9d9888a9fd29b207813 ^ 
0; 



wire Icec9f82ed5458da4eeaed077c58e91d3501f3067dda84ffba55bf76aee5404cd;
assign Icec9f82ed5458da4eeaed077c58e91d3501f3067dda84ffba55bf76aee5404cd = 
        y_nr_in[6] ^ 
        y_nr_in[9] ^ 
        y_nr_in[23] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[152] = 
Icec9f82ed5458da4eeaed077c58e91d3501f3067dda84ffba55bf76aee5404cd ^ 
0; 



wire I76ce9b3a35c82ecffdcbed87005640a6ffdf4cbb54e8d0280fe0fe1a47ec4153;
assign I76ce9b3a35c82ecffdcbed87005640a6ffdf4cbb54e8d0280fe0fe1a47ec4153 = 
        y_nr_in[7] ^ 
        y_nr_in[10] ^ 
        y_nr_in[20] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[153] = 
I76ce9b3a35c82ecffdcbed87005640a6ffdf4cbb54e8d0280fe0fe1a47ec4153 ^ 
0; 



wire I8c2a7cade24a98f62797ff246db0618e2031ec48015c9fbfdf2d6559c0536377;
assign I8c2a7cade24a98f62797ff246db0618e2031ec48015c9fbfdf2d6559c0536377 = 
        y_nr_in[4] ^ 
        y_nr_in[11] ^ 
        y_nr_in[21] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[154] = 
I8c2a7cade24a98f62797ff246db0618e2031ec48015c9fbfdf2d6559c0536377 ^ 
0; 



wire I39b9e146b624c47c64074bc132b83b1c4753edc20128f1b570ce586aa990a361;
assign I39b9e146b624c47c64074bc132b83b1c4753edc20128f1b570ce586aa990a361 = 
        y_nr_in[5] ^ 
        y_nr_in[8] ^ 
        y_nr_in[22] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[155] = 
I39b9e146b624c47c64074bc132b83b1c4753edc20128f1b570ce586aa990a361 ^ 
0; 



wire Ifc905cf9062222c11f5bd5d42856c5cd90aef46202ad17cac28de6a4c79188a0;
assign Ifc905cf9062222c11f5bd5d42856c5cd90aef46202ad17cac28de6a4c79188a0 = 
        y_nr_in[2] ^ 
        y_nr_in[16] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[156] = 
Ifc905cf9062222c11f5bd5d42856c5cd90aef46202ad17cac28de6a4c79188a0 ^ 
0; 



wire Ic0dedd09d29bc666a177c4f8f1aac7e081134411a025698ffe952de1a47cd4ea;
assign Ic0dedd09d29bc666a177c4f8f1aac7e081134411a025698ffe952de1a47cd4ea = 
        y_nr_in[3] ^ 
        y_nr_in[17] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[157] = 
Ic0dedd09d29bc666a177c4f8f1aac7e081134411a025698ffe952de1a47cd4ea ^ 
0; 



wire I6de6fe4c522d22a10ebba344a52da5f9938ab78ea1170471deda3bda1568dee4;
assign I6de6fe4c522d22a10ebba344a52da5f9938ab78ea1170471deda3bda1568dee4 = 
        y_nr_in[0] ^ 
        y_nr_in[18] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[158] = 
I6de6fe4c522d22a10ebba344a52da5f9938ab78ea1170471deda3bda1568dee4 ^ 
0; 



wire I9e6675aa0733abe263e12611ab91432a8c0c8845b2cc6470c0892e4bf592b952;
assign I9e6675aa0733abe263e12611ab91432a8c0c8845b2cc6470c0892e4bf592b952 = 
        y_nr_in[1] ^ 
        y_nr_in[19] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[159] = 
I9e6675aa0733abe263e12611ab91432a8c0c8845b2cc6470c0892e4bf592b952 ^ 
0; 



wire I98abd59ea45c34049379ee6f12c587b30a1da4de32d3070f7e69adc0f9fc4f4c;
assign I98abd59ea45c34049379ee6f12c587b30a1da4de32d3070f7e69adc0f9fc4f4c = 
        y_nr_in[11] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
0; 



wire I575f70d8cdf578436f1c4a28df7193c167c3afad67d511e7a50ea08ee201328e;
assign I575f70d8cdf578436f1c4a28df7193c167c3afad67d511e7a50ea08ee201328e = 
        y_nr_in[36] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[160] = 
I98abd59ea45c34049379ee6f12c587b30a1da4de32d3070f7e69adc0f9fc4f4c ^ 
I575f70d8cdf578436f1c4a28df7193c167c3afad67d511e7a50ea08ee201328e ^ 
0; 



wire Ib1b3643dc8b0921d548e81b347057dc6dd4d5ad184fc51c67819bfe36308f9c3;
assign Ib1b3643dc8b0921d548e81b347057dc6dd4d5ad184fc51c67819bfe36308f9c3 = 
        y_nr_in[8] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
0; 



wire I3f46b46cdea70163ead954ce7cddb9426ca8af6c4ba1cd67fb81b25318dd1a51;
assign I3f46b46cdea70163ead954ce7cddb9426ca8af6c4ba1cd67fb81b25318dd1a51 = 
        y_nr_in[37] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[161] = 
Ib1b3643dc8b0921d548e81b347057dc6dd4d5ad184fc51c67819bfe36308f9c3 ^ 
I3f46b46cdea70163ead954ce7cddb9426ca8af6c4ba1cd67fb81b25318dd1a51 ^ 
0; 



wire I85d19610152535540624bce37e88a0212ea10e49076fa932cf011349f6047bf0;
assign I85d19610152535540624bce37e88a0212ea10e49076fa932cf011349f6047bf0 = 
        y_nr_in[9] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
0; 



wire I64791be3ad9109e626afa75a98c8d0d792149c1d54016881809da5af04a0e384;
assign I64791be3ad9109e626afa75a98c8d0d792149c1d54016881809da5af04a0e384 = 
        y_nr_in[38] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[162] = 
I85d19610152535540624bce37e88a0212ea10e49076fa932cf011349f6047bf0 ^ 
I64791be3ad9109e626afa75a98c8d0d792149c1d54016881809da5af04a0e384 ^ 
0; 



wire I66114ebf49758b85fa88173cde89be4e76b7d35cadcea53c73018b32c968928e;
assign I66114ebf49758b85fa88173cde89be4e76b7d35cadcea53c73018b32c968928e = 
        y_nr_in[10] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
0; 



wire I09ab146dcfc299eb45c496708ef501ae7adaddb3366bc9346fe2d0787a2462ad;
assign I09ab146dcfc299eb45c496708ef501ae7adaddb3366bc9346fe2d0787a2462ad = 
        y_nr_in[39] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[163] = 
I66114ebf49758b85fa88173cde89be4e76b7d35cadcea53c73018b32c968928e ^ 
I09ab146dcfc299eb45c496708ef501ae7adaddb3366bc9346fe2d0787a2462ad ^ 
0; 



wire I2b7edf8e0a2ea23cfc68797e318e75ad0d62c5279dcdd15f1f16f72c4f231745;
assign I2b7edf8e0a2ea23cfc68797e318e75ad0d62c5279dcdd15f1f16f72c4f231745 = 
        y_nr_in[6] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[164] = 
I2b7edf8e0a2ea23cfc68797e318e75ad0d62c5279dcdd15f1f16f72c4f231745 ^ 
0; 



wire If1ee4ad64aeb58b31a2d63964b9e7d9ed3262b98d14da43b315d4fe70ed9f413;
assign If1ee4ad64aeb58b31a2d63964b9e7d9ed3262b98d14da43b315d4fe70ed9f413 = 
        y_nr_in[7] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[165] = 
If1ee4ad64aeb58b31a2d63964b9e7d9ed3262b98d14da43b315d4fe70ed9f413 ^ 
0; 



wire Iac791f5d19a7c542254f5d4b9b0fa6eef7eeb9b06f8a9916a3dc9da1bbda42ba;
assign Iac791f5d19a7c542254f5d4b9b0fa6eef7eeb9b06f8a9916a3dc9da1bbda42ba = 
        y_nr_in[4] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[166] = 
Iac791f5d19a7c542254f5d4b9b0fa6eef7eeb9b06f8a9916a3dc9da1bbda42ba ^ 
0; 



wire Ic03b2bba447638cf5ba15e511366289ff81c1b93d193a0538489ba2565296f0a;
assign Ic03b2bba447638cf5ba15e511366289ff81c1b93d193a0538489ba2565296f0a = 
        y_nr_in[5] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[167] = 
Ic03b2bba447638cf5ba15e511366289ff81c1b93d193a0538489ba2565296f0a ^ 
0; 



wire I21fa77e5a81f26a9e9f40d3f48bc2151c80fd24cbf574170f55573397644282d;
assign I21fa77e5a81f26a9e9f40d3f48bc2151c80fd24cbf574170f55573397644282d = 
        y_nr_in[2] ^ 
        y_nr_in[20] ^ 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[168] = 
I21fa77e5a81f26a9e9f40d3f48bc2151c80fd24cbf574170f55573397644282d ^ 
0; 



wire I449f4582a33cd58e5ccefc84e612ffd9c0633f3d01ad38ff1742c29bf0f7c25c;
assign I449f4582a33cd58e5ccefc84e612ffd9c0633f3d01ad38ff1742c29bf0f7c25c = 
        y_nr_in[3] ^ 
        y_nr_in[21] ^ 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[169] = 
I449f4582a33cd58e5ccefc84e612ffd9c0633f3d01ad38ff1742c29bf0f7c25c ^ 
0; 



wire Ib34a78bac7ebc1319b1cd7c2e0eeca290a8f43dd45e362c114d2abf34c96bd0a;
assign Ib34a78bac7ebc1319b1cd7c2e0eeca290a8f43dd45e362c114d2abf34c96bd0a = 
        y_nr_in[0] ^ 
        y_nr_in[22] ^ 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[170] = 
Ib34a78bac7ebc1319b1cd7c2e0eeca290a8f43dd45e362c114d2abf34c96bd0a ^ 
0; 



wire I90cc2339497d2123745cb7b6dafeee4bb82b658d8481848ed4c7fda1f9122847;
assign I90cc2339497d2123745cb7b6dafeee4bb82b658d8481848ed4c7fda1f9122847 = 
        y_nr_in[1] ^ 
        y_nr_in[23] ^ 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[171] = 
I90cc2339497d2123745cb7b6dafeee4bb82b658d8481848ed4c7fda1f9122847 ^ 
0; 



wire I2379c3cf6069c6a6c01dda309ba58d21db07f6ff7dfaa200d3a1171490be1f76;
assign I2379c3cf6069c6a6c01dda309ba58d21db07f6ff7dfaa200d3a1171490be1f76 = 
        y_nr_in[8] ^ 
        y_nr_in[28] ^ 
        y_nr_in[43] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[172] = 
I2379c3cf6069c6a6c01dda309ba58d21db07f6ff7dfaa200d3a1171490be1f76 ^ 
0; 



wire I01b54b2ba6f28e27f96a5789970db20747b171ec0f11942feb617aadb3158684;
assign I01b54b2ba6f28e27f96a5789970db20747b171ec0f11942feb617aadb3158684 = 
        y_nr_in[9] ^ 
        y_nr_in[29] ^ 
        y_nr_in[40] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[173] = 
I01b54b2ba6f28e27f96a5789970db20747b171ec0f11942feb617aadb3158684 ^ 
0; 



wire I73fef83985557bd1f985a3c72580cda280a34adfd5f4e457873105e3b67407af;
assign I73fef83985557bd1f985a3c72580cda280a34adfd5f4e457873105e3b67407af = 
        y_nr_in[10] ^ 
        y_nr_in[30] ^ 
        y_nr_in[41] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[174] = 
I73fef83985557bd1f985a3c72580cda280a34adfd5f4e457873105e3b67407af ^ 
0; 



wire I5ee7865d0d96d5a82c66f4e984e1f4a7cd7a81b695858843426fda2644271ad8;
assign I5ee7865d0d96d5a82c66f4e984e1f4a7cd7a81b695858843426fda2644271ad8 = 
        y_nr_in[11] ^ 
        y_nr_in[31] ^ 
        y_nr_in[42] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[175] = 
I5ee7865d0d96d5a82c66f4e984e1f4a7cd7a81b695858843426fda2644271ad8 ^ 
0; 



wire Iacfa6ee6cded64a7d31cd730732d3b456a57ed38b75501b687177eee4d719361;
assign Iacfa6ee6cded64a7d31cd730732d3b456a57ed38b75501b687177eee4d719361 = 
        y_nr_in[3] ^ 
        y_nr_in[49] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[176] = 
Iacfa6ee6cded64a7d31cd730732d3b456a57ed38b75501b687177eee4d719361 ^ 
0; 



wire I8600b085ca062f8f1f4ab56c916b9c72f7d0dd0d38b6358770f5d5ae0a1b6e40;
assign I8600b085ca062f8f1f4ab56c916b9c72f7d0dd0d38b6358770f5d5ae0a1b6e40 = 
        y_nr_in[0] ^ 
        y_nr_in[50] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[177] = 
I8600b085ca062f8f1f4ab56c916b9c72f7d0dd0d38b6358770f5d5ae0a1b6e40 ^ 
0; 



wire I609aa0a411c7d48c715eb8b67e3158773ad6e05beff6af2341bf5593f39cfa35;
assign I609aa0a411c7d48c715eb8b67e3158773ad6e05beff6af2341bf5593f39cfa35 = 
        y_nr_in[1] ^ 
        y_nr_in[51] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[178] = 
I609aa0a411c7d48c715eb8b67e3158773ad6e05beff6af2341bf5593f39cfa35 ^ 
0; 



wire Ia53e276cf2bc4394c0d60d008d8a2fdb115a6add3435fca9b741f1287db3771a;
assign Ia53e276cf2bc4394c0d60d008d8a2fdb115a6add3435fca9b741f1287db3771a = 
        y_nr_in[2] ^ 
        y_nr_in[48] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[179] = 
Ia53e276cf2bc4394c0d60d008d8a2fdb115a6add3435fca9b741f1287db3771a ^ 
0; 



wire Iaa91736b40c1da6fee66919f1ba7ebd9692d8f699aab5a9a09a7e531a8036fd7;
assign Iaa91736b40c1da6fee66919f1ba7ebd9692d8f699aab5a9a09a7e531a8036fd7 = 
        y_nr_in[5] ^ 
        y_nr_in[20] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[180] = 
Iaa91736b40c1da6fee66919f1ba7ebd9692d8f699aab5a9a09a7e531a8036fd7 ^ 
0; 



wire I8b760098076aa5efa7b2060215d72a18b64e940d44fb83a6d6e81fe514a96138;
assign I8b760098076aa5efa7b2060215d72a18b64e940d44fb83a6d6e81fe514a96138 = 
        y_nr_in[6] ^ 
        y_nr_in[21] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[181] = 
I8b760098076aa5efa7b2060215d72a18b64e940d44fb83a6d6e81fe514a96138 ^ 
0; 



wire I529ac8530c23147d2c629faa71227f6ab5cc03fc95fe5196ca4a2b105604c17c;
assign I529ac8530c23147d2c629faa71227f6ab5cc03fc95fe5196ca4a2b105604c17c = 
        y_nr_in[7] ^ 
        y_nr_in[22] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[182] = 
I529ac8530c23147d2c629faa71227f6ab5cc03fc95fe5196ca4a2b105604c17c ^ 
0; 



wire I888faef0c69f1ae9066f60c4a99e2998d4760949ff15485b10c3f36f973538fe;
assign I888faef0c69f1ae9066f60c4a99e2998d4760949ff15485b10c3f36f973538fe = 
        y_nr_in[4] ^ 
        y_nr_in[23] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[183] = 
I888faef0c69f1ae9066f60c4a99e2998d4760949ff15485b10c3f36f973538fe ^ 
0; 



wire I96199897315f2ca22ddb787dccffe917debdd3106222739bc8618e519540db1a;
assign I96199897315f2ca22ddb787dccffe917debdd3106222739bc8618e519540db1a = 
        y_nr_in[0] ^ 
        y_nr_in[10] ^ 
        y_nr_in[30] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[184] = 
I96199897315f2ca22ddb787dccffe917debdd3106222739bc8618e519540db1a ^ 
0; 



wire I3744dd6c478ebb3849b9b4e44a9acc8bea99a04cb6395c9e9ec022c94e6035d9;
assign I3744dd6c478ebb3849b9b4e44a9acc8bea99a04cb6395c9e9ec022c94e6035d9 = 
        y_nr_in[1] ^ 
        y_nr_in[11] ^ 
        y_nr_in[31] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[185] = 
I3744dd6c478ebb3849b9b4e44a9acc8bea99a04cb6395c9e9ec022c94e6035d9 ^ 
0; 



wire I6c042cef2bea157867bd9478e29443e036be26676910a02f2a6f6069dc5b45d1;
assign I6c042cef2bea157867bd9478e29443e036be26676910a02f2a6f6069dc5b45d1 = 
        y_nr_in[2] ^ 
        y_nr_in[8] ^ 
        y_nr_in[28] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[186] = 
I6c042cef2bea157867bd9478e29443e036be26676910a02f2a6f6069dc5b45d1 ^ 
0; 



wire Ib57055a68b1ea83edb5b34f75f5aaf9cb01466b28a1c09336d95aa815cadc521;
assign Ib57055a68b1ea83edb5b34f75f5aaf9cb01466b28a1c09336d95aa815cadc521 = 
        y_nr_in[3] ^ 
        y_nr_in[9] ^ 
        y_nr_in[29] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[187] = 
Ib57055a68b1ea83edb5b34f75f5aaf9cb01466b28a1c09336d95aa815cadc521 ^ 
0; 



wire Ibc0ceb87b8f0f1b8525525066f9b9cbd62e9c9c1099097b9e2fdefa04f4acbdc;
assign Ibc0ceb87b8f0f1b8525525066f9b9cbd62e9c9c1099097b9e2fdefa04f4acbdc = 
        y_nr_in[43] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[188] = 
Ibc0ceb87b8f0f1b8525525066f9b9cbd62e9c9c1099097b9e2fdefa04f4acbdc ^ 
0; 



wire Ic573c5aa926eac7cbd92972e9b5e6d2adcbcf1e7f205b6c3eab7266fee29723c;
assign Ic573c5aa926eac7cbd92972e9b5e6d2adcbcf1e7f205b6c3eab7266fee29723c = 
        y_nr_in[40] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[189] = 
Ic573c5aa926eac7cbd92972e9b5e6d2adcbcf1e7f205b6c3eab7266fee29723c ^ 
0; 



wire I1a16b74aaafc24f89442aaa83ebd6bcd0adb09b1cf759d3575e8092371153c8e;
assign I1a16b74aaafc24f89442aaa83ebd6bcd0adb09b1cf759d3575e8092371153c8e = 
        y_nr_in[41] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[190] = 
I1a16b74aaafc24f89442aaa83ebd6bcd0adb09b1cf759d3575e8092371153c8e ^ 
0; 



wire I69b75da9c7aebb51cd9d89fcd50d2404b3bcf738a926b2b01b6b6e0eddb9c405;
assign I69b75da9c7aebb51cd9d89fcd50d2404b3bcf738a926b2b01b6b6e0eddb9c405 = 
        y_nr_in[42] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[191] = 
I69b75da9c7aebb51cd9d89fcd50d2404b3bcf738a926b2b01b6b6e0eddb9c405 ^ 
0; 



wire Ib05d1701654f94cd661984dcac05add1c2981f5e90eeb05d0076094133a9ddc1;
assign Ib05d1701654f94cd661984dcac05add1c2981f5e90eeb05d0076094133a9ddc1 = 
        y_nr_in[7] ^ 
        y_nr_in[22] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[192] = 
Ib05d1701654f94cd661984dcac05add1c2981f5e90eeb05d0076094133a9ddc1 ^ 
0; 



wire If0dcab30c4290bb717e6d21c9329f7c40dddd600cc75b99c19a2c5ba5bb51a2a;
assign If0dcab30c4290bb717e6d21c9329f7c40dddd600cc75b99c19a2c5ba5bb51a2a = 
        y_nr_in[4] ^ 
        y_nr_in[23] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[193] = 
If0dcab30c4290bb717e6d21c9329f7c40dddd600cc75b99c19a2c5ba5bb51a2a ^ 
0; 



wire Ifa0479777741a438c934ea6aba5a37467646d68607af06c6d3bfc042ca1ed59a;
assign Ifa0479777741a438c934ea6aba5a37467646d68607af06c6d3bfc042ca1ed59a = 
        y_nr_in[5] ^ 
        y_nr_in[20] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[194] = 
Ifa0479777741a438c934ea6aba5a37467646d68607af06c6d3bfc042ca1ed59a ^ 
0; 



wire I8ccfe8bb3c0c31595051ddd6db64786a133ce480d501551b0f0c8a5b99dbf534;
assign I8ccfe8bb3c0c31595051ddd6db64786a133ce480d501551b0f0c8a5b99dbf534 = 
        y_nr_in[6] ^ 
        y_nr_in[21] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[195] = 
I8ccfe8bb3c0c31595051ddd6db64786a133ce480d501551b0f0c8a5b99dbf534 ^ 
0; 



wire Ia2545bbc6069b89225a087e83b6e706050d5fbbff16714460c8ee1e817856761;
assign Ia2545bbc6069b89225a087e83b6e706050d5fbbff16714460c8ee1e817856761 = 
        y_nr_in[3] ^ 
        y_nr_in[28] ^ 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[196] = 
Ia2545bbc6069b89225a087e83b6e706050d5fbbff16714460c8ee1e817856761 ^ 
0; 



wire I2d96c8f7c509d18560c55c41ae060aa3e042e1754ba886a5faf6815965dfbda3;
assign I2d96c8f7c509d18560c55c41ae060aa3e042e1754ba886a5faf6815965dfbda3 = 
        y_nr_in[0] ^ 
        y_nr_in[29] ^ 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[197] = 
I2d96c8f7c509d18560c55c41ae060aa3e042e1754ba886a5faf6815965dfbda3 ^ 
0; 



wire Idd111f41418abd6a786f907799544dbb55017bb42762dc8eb4cf6c165f9cb1b8;
assign Idd111f41418abd6a786f907799544dbb55017bb42762dc8eb4cf6c165f9cb1b8 = 
        y_nr_in[1] ^ 
        y_nr_in[30] ^ 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[198] = 
Idd111f41418abd6a786f907799544dbb55017bb42762dc8eb4cf6c165f9cb1b8 ^ 
0; 



wire Iaa6a9b2ddd88712a8261c2c79a566c78ab5b20e94f14c23c3e2989c55f33fd06;
assign Iaa6a9b2ddd88712a8261c2c79a566c78ab5b20e94f14c23c3e2989c55f33fd06 = 
        y_nr_in[2] ^ 
        y_nr_in[31] ^ 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[199] = 
Iaa6a9b2ddd88712a8261c2c79a566c78ab5b20e94f14c23c3e2989c55f33fd06 ^ 
0; 



wire I1c5586335326244e76a57c47a5ca57234bd1676901680aa4ab663ef9b7d0ea07;
assign I1c5586335326244e76a57c47a5ca57234bd1676901680aa4ab663ef9b7d0ea07 = 
        y_nr_in[8] ^ 
        y_nr_in[43] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[200] = 
I1c5586335326244e76a57c47a5ca57234bd1676901680aa4ab663ef9b7d0ea07 ^ 
0; 



wire I7fca90a1faddef8c5ba25cdd400149c765653bc4879735d29a155ffb74d2dc81;
assign I7fca90a1faddef8c5ba25cdd400149c765653bc4879735d29a155ffb74d2dc81 = 
        y_nr_in[9] ^ 
        y_nr_in[40] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[201] = 
I7fca90a1faddef8c5ba25cdd400149c765653bc4879735d29a155ffb74d2dc81 ^ 
0; 



wire Ib06281301a6f6e22076bbe24e642ac2435d593d04c77b75a5279cdc08fcf5fb5;
assign Ib06281301a6f6e22076bbe24e642ac2435d593d04c77b75a5279cdc08fcf5fb5 = 
        y_nr_in[10] ^ 
        y_nr_in[41] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[202] = 
Ib06281301a6f6e22076bbe24e642ac2435d593d04c77b75a5279cdc08fcf5fb5 ^ 
0; 



wire I7e3cd64b48229d2a2907ce88797145214f38d739f5f9a26227956ae9f489f15c;
assign I7e3cd64b48229d2a2907ce88797145214f38d739f5f9a26227956ae9f489f15c = 
        y_nr_in[11] ^ 
        y_nr_in[42] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[203] = 
I7e3cd64b48229d2a2907ce88797145214f38d739f5f9a26227956ae9f489f15c ^ 
0; 



wire I7c482c810c03a89f5abb373a710f4ec89e78b6a3ce6640867f7dc32afa8534ba;
assign I7c482c810c03a89f5abb373a710f4ec89e78b6a3ce6640867f7dc32afa8534ba = 
        y_nr_in[5] ^ 
        y_nr_in[21] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[204] = 
I7c482c810c03a89f5abb373a710f4ec89e78b6a3ce6640867f7dc32afa8534ba ^ 
0; 



wire I7f1ed42839bf4c9b361d4835dcd68bac43b61e2431bee34001bf6fb1c9d73f7f;
assign I7f1ed42839bf4c9b361d4835dcd68bac43b61e2431bee34001bf6fb1c9d73f7f = 
        y_nr_in[6] ^ 
        y_nr_in[22] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[205] = 
I7f1ed42839bf4c9b361d4835dcd68bac43b61e2431bee34001bf6fb1c9d73f7f ^ 
0; 



wire If4b9077bfa6665f80a0231cebab9a278dcb6e096508eb45465040b02beb8be14;
assign If4b9077bfa6665f80a0231cebab9a278dcb6e096508eb45465040b02beb8be14 = 
        y_nr_in[7] ^ 
        y_nr_in[23] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[206] = 
If4b9077bfa6665f80a0231cebab9a278dcb6e096508eb45465040b02beb8be14 ^ 
0; 



wire Id71a1b83f9cab8086700743fd1fe698a4c35a45b452e457545c9ca0d24caa1c4;
assign Id71a1b83f9cab8086700743fd1fe698a4c35a45b452e457545c9ca0d24caa1c4 = 
        y_nr_in[4] ^ 
        y_nr_in[20] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[207] = 
Id71a1b83f9cab8086700743fd1fe698a4c35a45b452e457545c9ca0d24caa1c4 ^ 
0; 



assign y_nr[n_int-1:n_int-m_int] = Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[n_int-1:n_int-m_int];
assign y_nr[n_int-m_int-1:0] = y_nr_in[n_int-m_int-1:0];
