 reg  ['h7:0] [$clog2('h7000+1)-1:0] I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c ;
