//`include "GF2_LDPC_fgallag_0x0000a_assign_inc.sv"
//always_comb begin
              I45c1a80dd59b47025bbf3f233589964b['h00000] = 
          (!fgallag_sel['h0000a]) ? 
                       If9057226a42b596a6dd2c84a37efff79['h00000] : //%
                       If9057226a42b596a6dd2c84a37efff79['h00001] ;
//end
//always_comb begin
              I45c1a80dd59b47025bbf3f233589964b['h00001] = 
          (!fgallag_sel['h0000a]) ? 
                       If9057226a42b596a6dd2c84a37efff79['h00002] : //%
                       If9057226a42b596a6dd2c84a37efff79['h00003] ;
//end
//always_comb begin
              I45c1a80dd59b47025bbf3f233589964b['h00002] = 
          (!fgallag_sel['h0000a]) ? 
                       If9057226a42b596a6dd2c84a37efff79['h00004] : //%
                       If9057226a42b596a6dd2c84a37efff79['h00005] ;
//end
//always_comb begin
              I45c1a80dd59b47025bbf3f233589964b['h00003] = 
          (!fgallag_sel['h0000a]) ? 
                       If9057226a42b596a6dd2c84a37efff79['h00006] : //%
                       If9057226a42b596a6dd2c84a37efff79['h00007] ;
//end
//always_comb begin
              I45c1a80dd59b47025bbf3f233589964b['h00004] = 
          (!fgallag_sel['h0000a]) ? 
                       If9057226a42b596a6dd2c84a37efff79['h00008] : //%
                       If9057226a42b596a6dd2c84a37efff79['h00009] ;
//end
//always_comb begin
              I45c1a80dd59b47025bbf3f233589964b['h00005] = 
          (!fgallag_sel['h0000a]) ? 
                       If9057226a42b596a6dd2c84a37efff79['h0000a] : //%
                       If9057226a42b596a6dd2c84a37efff79['h0000b] ;
//end
//always_comb begin
              I45c1a80dd59b47025bbf3f233589964b['h00006] = 
          (!fgallag_sel['h0000a]) ? 
                       If9057226a42b596a6dd2c84a37efff79['h0000c] : //%
                       If9057226a42b596a6dd2c84a37efff79['h0000d] ;
//end
//always_comb begin
              I45c1a80dd59b47025bbf3f233589964b['h00007] = 
          (!fgallag_sel['h0000a]) ? 
                       If9057226a42b596a6dd2c84a37efff79['h0000e] : //%
                       If9057226a42b596a6dd2c84a37efff79['h0000f] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00008] =  If9057226a42b596a6dd2c84a37efff79['h00010] ;
//end
//always_comb begin
              I45c1a80dd59b47025bbf3f233589964b['h00009] = 
          (!fgallag_sel['h0000a]) ? 
                       If9057226a42b596a6dd2c84a37efff79['h00012] : //%
                       If9057226a42b596a6dd2c84a37efff79['h00013] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0000a] =  If9057226a42b596a6dd2c84a37efff79['h00014] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0000b] =  If9057226a42b596a6dd2c84a37efff79['h00016] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0000c] =  If9057226a42b596a6dd2c84a37efff79['h00018] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0000d] =  If9057226a42b596a6dd2c84a37efff79['h0001a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0000e] =  If9057226a42b596a6dd2c84a37efff79['h0001c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0000f] =  If9057226a42b596a6dd2c84a37efff79['h0001e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00010] =  If9057226a42b596a6dd2c84a37efff79['h00020] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00011] =  If9057226a42b596a6dd2c84a37efff79['h00022] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00012] =  If9057226a42b596a6dd2c84a37efff79['h00024] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00013] =  If9057226a42b596a6dd2c84a37efff79['h00026] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00014] =  If9057226a42b596a6dd2c84a37efff79['h00028] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00015] =  If9057226a42b596a6dd2c84a37efff79['h0002a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00016] =  If9057226a42b596a6dd2c84a37efff79['h0002c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00017] =  If9057226a42b596a6dd2c84a37efff79['h0002e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00018] =  If9057226a42b596a6dd2c84a37efff79['h00030] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00019] =  If9057226a42b596a6dd2c84a37efff79['h00032] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0001a] =  If9057226a42b596a6dd2c84a37efff79['h00034] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0001b] =  If9057226a42b596a6dd2c84a37efff79['h00036] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0001c] =  If9057226a42b596a6dd2c84a37efff79['h00038] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0001d] =  If9057226a42b596a6dd2c84a37efff79['h0003a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0001e] =  If9057226a42b596a6dd2c84a37efff79['h0003c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0001f] =  If9057226a42b596a6dd2c84a37efff79['h0003e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00020] =  If9057226a42b596a6dd2c84a37efff79['h00040] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00021] =  If9057226a42b596a6dd2c84a37efff79['h00042] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00022] =  If9057226a42b596a6dd2c84a37efff79['h00044] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00023] =  If9057226a42b596a6dd2c84a37efff79['h00046] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00024] =  If9057226a42b596a6dd2c84a37efff79['h00048] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00025] =  If9057226a42b596a6dd2c84a37efff79['h0004a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00026] =  If9057226a42b596a6dd2c84a37efff79['h0004c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00027] =  If9057226a42b596a6dd2c84a37efff79['h0004e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00028] =  If9057226a42b596a6dd2c84a37efff79['h00050] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00029] =  If9057226a42b596a6dd2c84a37efff79['h00052] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0002a] =  If9057226a42b596a6dd2c84a37efff79['h00054] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0002b] =  If9057226a42b596a6dd2c84a37efff79['h00056] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0002c] =  If9057226a42b596a6dd2c84a37efff79['h00058] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0002d] =  If9057226a42b596a6dd2c84a37efff79['h0005a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0002e] =  If9057226a42b596a6dd2c84a37efff79['h0005c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0002f] =  If9057226a42b596a6dd2c84a37efff79['h0005e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00030] =  If9057226a42b596a6dd2c84a37efff79['h00060] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00031] =  If9057226a42b596a6dd2c84a37efff79['h00062] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00032] =  If9057226a42b596a6dd2c84a37efff79['h00064] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00033] =  If9057226a42b596a6dd2c84a37efff79['h00066] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00034] =  If9057226a42b596a6dd2c84a37efff79['h00068] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00035] =  If9057226a42b596a6dd2c84a37efff79['h0006a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00036] =  If9057226a42b596a6dd2c84a37efff79['h0006c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00037] =  If9057226a42b596a6dd2c84a37efff79['h0006e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00038] =  If9057226a42b596a6dd2c84a37efff79['h00070] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00039] =  If9057226a42b596a6dd2c84a37efff79['h00072] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0003a] =  If9057226a42b596a6dd2c84a37efff79['h00074] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0003b] =  If9057226a42b596a6dd2c84a37efff79['h00076] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0003c] =  If9057226a42b596a6dd2c84a37efff79['h00078] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0003d] =  If9057226a42b596a6dd2c84a37efff79['h0007a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0003e] =  If9057226a42b596a6dd2c84a37efff79['h0007c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0003f] =  If9057226a42b596a6dd2c84a37efff79['h0007e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00040] =  If9057226a42b596a6dd2c84a37efff79['h00080] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00041] =  If9057226a42b596a6dd2c84a37efff79['h00082] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00042] =  If9057226a42b596a6dd2c84a37efff79['h00084] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00043] =  If9057226a42b596a6dd2c84a37efff79['h00086] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00044] =  If9057226a42b596a6dd2c84a37efff79['h00088] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00045] =  If9057226a42b596a6dd2c84a37efff79['h0008a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00046] =  If9057226a42b596a6dd2c84a37efff79['h0008c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00047] =  If9057226a42b596a6dd2c84a37efff79['h0008e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00048] =  If9057226a42b596a6dd2c84a37efff79['h00090] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00049] =  If9057226a42b596a6dd2c84a37efff79['h00092] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0004a] =  If9057226a42b596a6dd2c84a37efff79['h00094] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0004b] =  If9057226a42b596a6dd2c84a37efff79['h00096] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0004c] =  If9057226a42b596a6dd2c84a37efff79['h00098] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0004d] =  If9057226a42b596a6dd2c84a37efff79['h0009a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0004e] =  If9057226a42b596a6dd2c84a37efff79['h0009c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0004f] =  If9057226a42b596a6dd2c84a37efff79['h0009e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00050] =  If9057226a42b596a6dd2c84a37efff79['h000a0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00051] =  If9057226a42b596a6dd2c84a37efff79['h000a2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00052] =  If9057226a42b596a6dd2c84a37efff79['h000a4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00053] =  If9057226a42b596a6dd2c84a37efff79['h000a6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00054] =  If9057226a42b596a6dd2c84a37efff79['h000a8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00055] =  If9057226a42b596a6dd2c84a37efff79['h000aa] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00056] =  If9057226a42b596a6dd2c84a37efff79['h000ac] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00057] =  If9057226a42b596a6dd2c84a37efff79['h000ae] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00058] =  If9057226a42b596a6dd2c84a37efff79['h000b0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00059] =  If9057226a42b596a6dd2c84a37efff79['h000b2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0005a] =  If9057226a42b596a6dd2c84a37efff79['h000b4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0005b] =  If9057226a42b596a6dd2c84a37efff79['h000b6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0005c] =  If9057226a42b596a6dd2c84a37efff79['h000b8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0005d] =  If9057226a42b596a6dd2c84a37efff79['h000ba] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0005e] =  If9057226a42b596a6dd2c84a37efff79['h000bc] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0005f] =  If9057226a42b596a6dd2c84a37efff79['h000be] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00060] =  If9057226a42b596a6dd2c84a37efff79['h000c0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00061] =  If9057226a42b596a6dd2c84a37efff79['h000c2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00062] =  If9057226a42b596a6dd2c84a37efff79['h000c4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00063] =  If9057226a42b596a6dd2c84a37efff79['h000c6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00064] =  If9057226a42b596a6dd2c84a37efff79['h000c8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00065] =  If9057226a42b596a6dd2c84a37efff79['h000ca] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00066] =  If9057226a42b596a6dd2c84a37efff79['h000cc] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00067] =  If9057226a42b596a6dd2c84a37efff79['h000ce] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00068] =  If9057226a42b596a6dd2c84a37efff79['h000d0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00069] =  If9057226a42b596a6dd2c84a37efff79['h000d2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0006a] =  If9057226a42b596a6dd2c84a37efff79['h000d4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0006b] =  If9057226a42b596a6dd2c84a37efff79['h000d6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0006c] =  If9057226a42b596a6dd2c84a37efff79['h000d8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0006d] =  If9057226a42b596a6dd2c84a37efff79['h000da] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0006e] =  If9057226a42b596a6dd2c84a37efff79['h000dc] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0006f] =  If9057226a42b596a6dd2c84a37efff79['h000de] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00070] =  If9057226a42b596a6dd2c84a37efff79['h000e0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00071] =  If9057226a42b596a6dd2c84a37efff79['h000e2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00072] =  If9057226a42b596a6dd2c84a37efff79['h000e4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00073] =  If9057226a42b596a6dd2c84a37efff79['h000e6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00074] =  If9057226a42b596a6dd2c84a37efff79['h000e8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00075] =  If9057226a42b596a6dd2c84a37efff79['h000ea] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00076] =  If9057226a42b596a6dd2c84a37efff79['h000ec] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00077] =  If9057226a42b596a6dd2c84a37efff79['h000ee] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00078] =  If9057226a42b596a6dd2c84a37efff79['h000f0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00079] =  If9057226a42b596a6dd2c84a37efff79['h000f2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0007a] =  If9057226a42b596a6dd2c84a37efff79['h000f4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0007b] =  If9057226a42b596a6dd2c84a37efff79['h000f6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0007c] =  If9057226a42b596a6dd2c84a37efff79['h000f8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0007d] =  If9057226a42b596a6dd2c84a37efff79['h000fa] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0007e] =  If9057226a42b596a6dd2c84a37efff79['h000fc] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0007f] =  If9057226a42b596a6dd2c84a37efff79['h000fe] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00080] =  If9057226a42b596a6dd2c84a37efff79['h00100] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00081] =  If9057226a42b596a6dd2c84a37efff79['h00102] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00082] =  If9057226a42b596a6dd2c84a37efff79['h00104] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00083] =  If9057226a42b596a6dd2c84a37efff79['h00106] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00084] =  If9057226a42b596a6dd2c84a37efff79['h00108] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00085] =  If9057226a42b596a6dd2c84a37efff79['h0010a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00086] =  If9057226a42b596a6dd2c84a37efff79['h0010c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00087] =  If9057226a42b596a6dd2c84a37efff79['h0010e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00088] =  If9057226a42b596a6dd2c84a37efff79['h00110] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00089] =  If9057226a42b596a6dd2c84a37efff79['h00112] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0008a] =  If9057226a42b596a6dd2c84a37efff79['h00114] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0008b] =  If9057226a42b596a6dd2c84a37efff79['h00116] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0008c] =  If9057226a42b596a6dd2c84a37efff79['h00118] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0008d] =  If9057226a42b596a6dd2c84a37efff79['h0011a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0008e] =  If9057226a42b596a6dd2c84a37efff79['h0011c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0008f] =  If9057226a42b596a6dd2c84a37efff79['h0011e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00090] =  If9057226a42b596a6dd2c84a37efff79['h00120] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00091] =  If9057226a42b596a6dd2c84a37efff79['h00122] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00092] =  If9057226a42b596a6dd2c84a37efff79['h00124] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00093] =  If9057226a42b596a6dd2c84a37efff79['h00126] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00094] =  If9057226a42b596a6dd2c84a37efff79['h00128] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00095] =  If9057226a42b596a6dd2c84a37efff79['h0012a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00096] =  If9057226a42b596a6dd2c84a37efff79['h0012c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00097] =  If9057226a42b596a6dd2c84a37efff79['h0012e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00098] =  If9057226a42b596a6dd2c84a37efff79['h00130] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h00099] =  If9057226a42b596a6dd2c84a37efff79['h00132] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0009a] =  If9057226a42b596a6dd2c84a37efff79['h00134] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0009b] =  If9057226a42b596a6dd2c84a37efff79['h00136] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0009c] =  If9057226a42b596a6dd2c84a37efff79['h00138] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0009d] =  If9057226a42b596a6dd2c84a37efff79['h0013a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0009e] =  If9057226a42b596a6dd2c84a37efff79['h0013c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h0009f] =  If9057226a42b596a6dd2c84a37efff79['h0013e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000a0] =  If9057226a42b596a6dd2c84a37efff79['h00140] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000a1] =  If9057226a42b596a6dd2c84a37efff79['h00142] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000a2] =  If9057226a42b596a6dd2c84a37efff79['h00144] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000a3] =  If9057226a42b596a6dd2c84a37efff79['h00146] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000a4] =  If9057226a42b596a6dd2c84a37efff79['h00148] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000a5] =  If9057226a42b596a6dd2c84a37efff79['h0014a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000a6] =  If9057226a42b596a6dd2c84a37efff79['h0014c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000a7] =  If9057226a42b596a6dd2c84a37efff79['h0014e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000a8] =  If9057226a42b596a6dd2c84a37efff79['h00150] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000a9] =  If9057226a42b596a6dd2c84a37efff79['h00152] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000aa] =  If9057226a42b596a6dd2c84a37efff79['h00154] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ab] =  If9057226a42b596a6dd2c84a37efff79['h00156] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ac] =  If9057226a42b596a6dd2c84a37efff79['h00158] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ad] =  If9057226a42b596a6dd2c84a37efff79['h0015a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ae] =  If9057226a42b596a6dd2c84a37efff79['h0015c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000af] =  If9057226a42b596a6dd2c84a37efff79['h0015e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000b0] =  If9057226a42b596a6dd2c84a37efff79['h00160] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000b1] =  If9057226a42b596a6dd2c84a37efff79['h00162] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000b2] =  If9057226a42b596a6dd2c84a37efff79['h00164] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000b3] =  If9057226a42b596a6dd2c84a37efff79['h00166] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000b4] =  If9057226a42b596a6dd2c84a37efff79['h00168] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000b5] =  If9057226a42b596a6dd2c84a37efff79['h0016a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000b6] =  If9057226a42b596a6dd2c84a37efff79['h0016c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000b7] =  If9057226a42b596a6dd2c84a37efff79['h0016e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000b8] =  If9057226a42b596a6dd2c84a37efff79['h00170] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000b9] =  If9057226a42b596a6dd2c84a37efff79['h00172] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ba] =  If9057226a42b596a6dd2c84a37efff79['h00174] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000bb] =  If9057226a42b596a6dd2c84a37efff79['h00176] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000bc] =  If9057226a42b596a6dd2c84a37efff79['h00178] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000bd] =  If9057226a42b596a6dd2c84a37efff79['h0017a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000be] =  If9057226a42b596a6dd2c84a37efff79['h0017c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000bf] =  If9057226a42b596a6dd2c84a37efff79['h0017e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000c0] =  If9057226a42b596a6dd2c84a37efff79['h00180] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000c1] =  If9057226a42b596a6dd2c84a37efff79['h00182] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000c2] =  If9057226a42b596a6dd2c84a37efff79['h00184] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000c3] =  If9057226a42b596a6dd2c84a37efff79['h00186] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000c4] =  If9057226a42b596a6dd2c84a37efff79['h00188] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000c5] =  If9057226a42b596a6dd2c84a37efff79['h0018a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000c6] =  If9057226a42b596a6dd2c84a37efff79['h0018c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000c7] =  If9057226a42b596a6dd2c84a37efff79['h0018e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000c8] =  If9057226a42b596a6dd2c84a37efff79['h00190] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000c9] =  If9057226a42b596a6dd2c84a37efff79['h00192] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ca] =  If9057226a42b596a6dd2c84a37efff79['h00194] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000cb] =  If9057226a42b596a6dd2c84a37efff79['h00196] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000cc] =  If9057226a42b596a6dd2c84a37efff79['h00198] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000cd] =  If9057226a42b596a6dd2c84a37efff79['h0019a] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ce] =  If9057226a42b596a6dd2c84a37efff79['h0019c] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000cf] =  If9057226a42b596a6dd2c84a37efff79['h0019e] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000d0] =  If9057226a42b596a6dd2c84a37efff79['h001a0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000d1] =  If9057226a42b596a6dd2c84a37efff79['h001a2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000d2] =  If9057226a42b596a6dd2c84a37efff79['h001a4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000d3] =  If9057226a42b596a6dd2c84a37efff79['h001a6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000d4] =  If9057226a42b596a6dd2c84a37efff79['h001a8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000d5] =  If9057226a42b596a6dd2c84a37efff79['h001aa] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000d6] =  If9057226a42b596a6dd2c84a37efff79['h001ac] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000d7] =  If9057226a42b596a6dd2c84a37efff79['h001ae] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000d8] =  If9057226a42b596a6dd2c84a37efff79['h001b0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000d9] =  If9057226a42b596a6dd2c84a37efff79['h001b2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000da] =  If9057226a42b596a6dd2c84a37efff79['h001b4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000db] =  If9057226a42b596a6dd2c84a37efff79['h001b6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000dc] =  If9057226a42b596a6dd2c84a37efff79['h001b8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000dd] =  If9057226a42b596a6dd2c84a37efff79['h001ba] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000de] =  If9057226a42b596a6dd2c84a37efff79['h001bc] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000df] =  If9057226a42b596a6dd2c84a37efff79['h001be] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000e0] =  If9057226a42b596a6dd2c84a37efff79['h001c0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000e1] =  If9057226a42b596a6dd2c84a37efff79['h001c2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000e2] =  If9057226a42b596a6dd2c84a37efff79['h001c4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000e3] =  If9057226a42b596a6dd2c84a37efff79['h001c6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000e4] =  If9057226a42b596a6dd2c84a37efff79['h001c8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000e5] =  If9057226a42b596a6dd2c84a37efff79['h001ca] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000e6] =  If9057226a42b596a6dd2c84a37efff79['h001cc] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000e7] =  If9057226a42b596a6dd2c84a37efff79['h001ce] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000e8] =  If9057226a42b596a6dd2c84a37efff79['h001d0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000e9] =  If9057226a42b596a6dd2c84a37efff79['h001d2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ea] =  If9057226a42b596a6dd2c84a37efff79['h001d4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000eb] =  If9057226a42b596a6dd2c84a37efff79['h001d6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ec] =  If9057226a42b596a6dd2c84a37efff79['h001d8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ed] =  If9057226a42b596a6dd2c84a37efff79['h001da] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ee] =  If9057226a42b596a6dd2c84a37efff79['h001dc] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ef] =  If9057226a42b596a6dd2c84a37efff79['h001de] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000f0] =  If9057226a42b596a6dd2c84a37efff79['h001e0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000f1] =  If9057226a42b596a6dd2c84a37efff79['h001e2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000f2] =  If9057226a42b596a6dd2c84a37efff79['h001e4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000f3] =  If9057226a42b596a6dd2c84a37efff79['h001e6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000f4] =  If9057226a42b596a6dd2c84a37efff79['h001e8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000f5] =  If9057226a42b596a6dd2c84a37efff79['h001ea] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000f6] =  If9057226a42b596a6dd2c84a37efff79['h001ec] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000f7] =  If9057226a42b596a6dd2c84a37efff79['h001ee] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000f8] =  If9057226a42b596a6dd2c84a37efff79['h001f0] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000f9] =  If9057226a42b596a6dd2c84a37efff79['h001f2] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000fa] =  If9057226a42b596a6dd2c84a37efff79['h001f4] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000fb] =  If9057226a42b596a6dd2c84a37efff79['h001f6] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000fc] =  If9057226a42b596a6dd2c84a37efff79['h001f8] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000fd] =  If9057226a42b596a6dd2c84a37efff79['h001fa] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000fe] =  If9057226a42b596a6dd2c84a37efff79['h001fc] ;
//end
//always_comb begin // 
               I45c1a80dd59b47025bbf3f233589964b['h000ff] =  If9057226a42b596a6dd2c84a37efff79['h001fe] ;
//end
