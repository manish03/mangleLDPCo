 reg  ['h1f:0] [$clog2('h7000+1)-1:0] Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478 ;
