 reg  ['h7f:0] [$clog2('h7000+1)-1:0] Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96 ;
