 reg  ['hf:0] [$clog2('h7000+1)-1:0] I9d96959b6b7fd9b9e978d3f23959e9e1 ;
