 reg  ['h1ff:0] [$clog2('h7000+1)-1:0] Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd ;
