 reg  ['h1ff:0] [$clog2('h7000+1)-1:0] If9057226a42b596a6dd2c84a37efff79 ;
