//`include "GF2_LDPC_fgallag_0x00008_assign_inc.sv"
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00000] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00000] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00001] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00001] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00002] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00003] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00002] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00004] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00005] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00003] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00006] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00007] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00004] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00008] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00009] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00005] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000a] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000b] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00006] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000c] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000d] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00007] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000e] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000f] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00008] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00010] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00011] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00009] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00012] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00013] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0000a] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00014] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00015] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0000b] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00016] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00017] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0000c] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00018] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00019] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0000d] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001a] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001b] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0000e] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001c] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001d] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0000f] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001e] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001f] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00010] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00020] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00021] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00011] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00022] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00023] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00012] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00024] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00025] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00013] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00026] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00027] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00014] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00028] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00029] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00015] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002a] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002b] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00016] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002c] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002d] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00017] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002e] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002f] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00018] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00030] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00031] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00019] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00032] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00033] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0001a] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00034] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00035] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0001b] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00036] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00037] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0001c] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00038] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00039] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0001d] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003a] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003b] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0001e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003c] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h0001f] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003e] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003f] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00020] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00040] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00021] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00042] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00022] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00044] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00023] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00046] ;
//end
//always_comb begin
              Icff8af1f5c3ae89ef95ed8451273154b['h00024] = 
          (!fgallag_sel['h00008]) ? 
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00048] : //%
                       Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00049] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00025] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0004a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00026] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0004c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00027] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0004e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00028] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00050] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00029] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00052] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0002a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00054] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0002b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00056] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0002c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00058] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0002d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0005a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0002e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0005c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0002f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0005e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00030] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00060] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00031] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00062] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00032] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00064] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00033] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00066] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00034] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00068] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00035] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0006a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00036] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0006c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00037] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0006e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00038] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00070] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00039] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00072] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0003a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00074] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0003b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00076] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0003c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00078] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0003d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0007a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0003e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0007c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0003f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0007e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00040] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00080] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00041] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00082] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00042] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00084] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00043] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00086] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00044] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00088] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00045] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0008a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00046] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0008c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00047] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0008e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00048] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00090] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00049] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00092] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0004a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00094] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0004b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00096] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0004c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00098] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0004d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0009a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0004e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0009c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0004f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0009e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00050] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00051] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00052] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00053] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00054] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00055] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000aa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00056] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ac] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00057] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ae] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00058] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00059] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0005a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0005b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0005c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0005d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ba] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0005e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000bc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0005f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000be] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00060] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00061] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00062] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00063] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00064] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00065] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ca] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00066] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000cc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00067] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ce] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00068] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00069] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0006a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0006b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0006c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0006d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000da] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0006e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000dc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0006f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000de] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00070] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00071] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00072] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00073] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00074] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00075] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ea] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00076] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ec] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00077] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ee] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00078] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00079] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0007a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0007b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0007c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0007d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000fa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0007e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000fc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0007f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000fe] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00080] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00100] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00081] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00102] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00082] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00104] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00083] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00106] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00084] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00108] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00085] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0010a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00086] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0010c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00087] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0010e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00088] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00110] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00089] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00112] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0008a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00114] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0008b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00116] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0008c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00118] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0008d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0011a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0008e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0011c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0008f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0011e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00090] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00120] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00091] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00122] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00092] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00124] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00093] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00126] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00094] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00128] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00095] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0012a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00096] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0012c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00097] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0012e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00098] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00130] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00099] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00132] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0009a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00134] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0009b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00136] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0009c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00138] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0009d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0013a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0009e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0013c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0009f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0013e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000a0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00140] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000a1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00142] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000a2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00144] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000a3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00146] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000a4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00148] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000a5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0014a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000a6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0014c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000a7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0014e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000a8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00150] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000a9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00152] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000aa] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00154] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ab] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00156] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ac] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00158] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ad] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0015a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ae] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0015c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000af] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0015e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000b0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00160] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000b1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00162] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000b2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00164] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000b3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00166] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000b4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00168] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000b5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0016a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000b6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0016c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000b7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0016e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000b8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00170] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000b9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00172] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ba] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00174] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000bb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00176] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000bc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00178] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000bd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0017a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000be] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0017c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000bf] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0017e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000c0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00180] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000c1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00182] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000c2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00184] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000c3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00186] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000c4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00188] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000c5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0018a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000c6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0018c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000c7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0018e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000c8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00190] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000c9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00192] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ca] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00194] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000cb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00196] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000cc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00198] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000cd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0019a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ce] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0019c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000cf] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0019e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000d0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000d1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000d2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000d3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000d4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000d5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001aa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000d6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ac] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000d7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ae] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000d8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000d9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000da] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000db] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000dc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000dd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ba] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000de] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001bc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000df] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001be] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000e0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000e1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000e2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000e3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000e4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000e5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ca] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000e6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001cc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000e7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ce] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000e8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000e9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ea] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000eb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ec] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ed] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001da] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ee] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001dc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ef] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001de] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000f0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000f1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000f2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000f3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000f4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000f5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ea] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000f6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ec] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000f7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ee] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000f8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000f9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000fa] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000fb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000fc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000fd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001fa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000fe] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001fc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h000ff] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001fe] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00100] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00200] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00101] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00202] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00102] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00204] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00103] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00206] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00104] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00208] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00105] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0020a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00106] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0020c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00107] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0020e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00108] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00210] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00109] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00212] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0010a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00214] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0010b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00216] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0010c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00218] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0010d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0021a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0010e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0021c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0010f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0021e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00110] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00220] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00111] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00222] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00112] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00224] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00113] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00226] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00114] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00228] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00115] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0022a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00116] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0022c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00117] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0022e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00118] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00230] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00119] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00232] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0011a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00234] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0011b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00236] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0011c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00238] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0011d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0023a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0011e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0023c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0011f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0023e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00120] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00240] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00121] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00242] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00122] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00244] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00123] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00246] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00124] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00248] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00125] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0024a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00126] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0024c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00127] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0024e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00128] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00250] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00129] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00252] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0012a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00254] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0012b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00256] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0012c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00258] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0012d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0025a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0012e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0025c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0012f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0025e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00130] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00260] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00131] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00262] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00132] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00264] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00133] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00266] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00134] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00268] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00135] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0026a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00136] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0026c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00137] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0026e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00138] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00270] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00139] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00272] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0013a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00274] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0013b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00276] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0013c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00278] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0013d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0027a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0013e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0027c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0013f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0027e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00140] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00280] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00141] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00282] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00142] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00284] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00143] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00286] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00144] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00288] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00145] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0028a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00146] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0028c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00147] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0028e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00148] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00290] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00149] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00292] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0014a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00294] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0014b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00296] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0014c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00298] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0014d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0029a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0014e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0029c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0014f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0029e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00150] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00151] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00152] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00153] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00154] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00155] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002aa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00156] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ac] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00157] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ae] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00158] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00159] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0015a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0015b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0015c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0015d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ba] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0015e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002bc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0015f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002be] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00160] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00161] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00162] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00163] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00164] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00165] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ca] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00166] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002cc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00167] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ce] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00168] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00169] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0016a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0016b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0016c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0016d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002da] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0016e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002dc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0016f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002de] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00170] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00171] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00172] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00173] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00174] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00175] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ea] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00176] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ec] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00177] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ee] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00178] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00179] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0017a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0017b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0017c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0017d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002fa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0017e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002fc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0017f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002fe] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00180] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00300] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00181] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00302] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00182] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00304] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00183] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00306] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00184] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00308] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00185] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0030a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00186] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0030c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00187] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0030e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00188] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00310] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00189] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00312] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0018a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00314] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0018b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00316] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0018c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00318] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0018d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0031a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0018e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0031c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0018f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0031e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00190] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00320] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00191] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00322] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00192] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00324] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00193] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00326] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00194] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00328] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00195] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0032a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00196] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0032c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00197] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0032e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00198] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00330] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00199] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00332] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0019a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00334] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0019b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00336] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0019c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00338] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0019d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0033a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0019e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0033c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0019f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0033e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001a0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00340] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001a1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00342] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001a2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00344] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001a3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00346] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001a4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00348] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001a5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0034a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001a6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0034c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001a7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0034e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001a8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00350] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001a9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00352] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001aa] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00354] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ab] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00356] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ac] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00358] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ad] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0035a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ae] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0035c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001af] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0035e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001b0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00360] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001b1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00362] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001b2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00364] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001b3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00366] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001b4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00368] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001b5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0036a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001b6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0036c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001b7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0036e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001b8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00370] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001b9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00372] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ba] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00374] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001bb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00376] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001bc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00378] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001bd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0037a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001be] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0037c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001bf] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0037e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001c0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00380] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001c1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00382] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001c2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00384] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001c3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00386] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001c4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00388] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001c5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0038a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001c6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0038c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001c7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0038e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001c8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00390] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001c9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00392] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ca] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00394] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001cb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00396] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001cc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00398] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001cd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0039a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ce] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0039c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001cf] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0039e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001d0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001d1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001d2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001d3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001d4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001d5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003aa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001d6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ac] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001d7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ae] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001d8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001d9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001da] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001db] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001dc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001dd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ba] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001de] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003bc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001df] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003be] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001e0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001e1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001e2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001e3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001e4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001e5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ca] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001e6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003cc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001e7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ce] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001e8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001e9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ea] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001eb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ec] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ed] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003da] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ee] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003dc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ef] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003de] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001f0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001f1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001f2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001f3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001f4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001f5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ea] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001f6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ec] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001f7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ee] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001f8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001f9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001fa] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001fb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001fc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001fd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003fa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001fe] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003fc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h001ff] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003fe] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00200] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00400] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00201] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00402] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00202] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00404] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00203] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00406] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00204] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00408] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00205] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0040a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00206] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0040c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00207] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0040e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00208] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00410] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00209] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00412] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0020a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00414] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0020b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00416] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0020c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00418] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0020d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0041a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0020e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0041c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0020f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0041e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00210] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00420] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00211] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00422] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00212] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00424] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00213] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00426] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00214] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00428] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00215] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0042a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00216] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0042c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00217] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0042e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00218] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00430] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00219] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00432] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0021a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00434] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0021b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00436] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0021c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00438] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0021d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0043a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0021e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0043c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0021f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0043e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00220] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00440] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00221] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00442] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00222] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00444] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00223] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00446] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00224] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00448] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00225] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0044a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00226] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0044c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00227] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0044e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00228] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00450] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00229] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00452] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0022a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00454] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0022b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00456] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0022c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00458] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0022d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0045a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0022e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0045c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0022f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0045e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00230] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00460] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00231] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00462] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00232] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00464] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00233] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00466] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00234] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00468] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00235] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0046a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00236] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0046c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00237] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0046e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00238] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00470] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00239] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00472] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0023a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00474] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0023b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00476] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0023c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00478] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0023d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0047a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0023e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0047c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0023f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0047e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00240] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00480] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00241] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00482] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00242] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00484] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00243] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00486] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00244] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00488] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00245] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0048a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00246] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0048c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00247] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0048e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00248] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00490] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00249] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00492] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0024a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00494] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0024b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00496] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0024c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00498] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0024d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0049a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0024e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0049c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0024f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0049e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00250] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00251] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00252] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00253] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00254] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00255] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004aa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00256] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ac] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00257] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ae] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00258] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00259] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0025a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0025b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0025c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0025d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ba] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0025e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004bc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0025f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004be] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00260] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00261] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00262] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00263] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00264] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00265] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ca] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00266] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004cc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00267] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ce] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00268] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00269] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0026a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0026b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0026c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0026d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004da] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0026e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004dc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0026f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004de] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00270] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00271] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00272] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00273] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00274] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00275] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ea] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00276] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ec] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00277] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ee] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00278] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00279] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0027a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0027b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0027c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0027d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004fa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0027e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004fc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0027f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004fe] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00280] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00500] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00281] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00502] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00282] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00504] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00283] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00506] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00284] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00508] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00285] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0050a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00286] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0050c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00287] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0050e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00288] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00510] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00289] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00512] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0028a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00514] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0028b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00516] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0028c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00518] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0028d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0051a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0028e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0051c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0028f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0051e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00290] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00520] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00291] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00522] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00292] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00524] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00293] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00526] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00294] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00528] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00295] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0052a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00296] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0052c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00297] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0052e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00298] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00530] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00299] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00532] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0029a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00534] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0029b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00536] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0029c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00538] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0029d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0053a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0029e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0053c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0029f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0053e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002a0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00540] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002a1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00542] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002a2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00544] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002a3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00546] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002a4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00548] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002a5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0054a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002a6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0054c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002a7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0054e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002a8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00550] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002a9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00552] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002aa] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00554] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ab] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00556] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ac] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00558] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ad] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0055a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ae] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0055c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002af] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0055e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002b0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00560] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002b1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00562] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002b2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00564] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002b3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00566] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002b4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00568] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002b5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0056a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002b6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0056c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002b7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0056e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002b8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00570] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002b9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00572] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ba] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00574] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002bb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00576] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002bc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00578] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002bd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0057a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002be] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0057c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002bf] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0057e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002c0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00580] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002c1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00582] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002c2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00584] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002c3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00586] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002c4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00588] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002c5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0058a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002c6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0058c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002c7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0058e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002c8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00590] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002c9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00592] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ca] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00594] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002cb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00596] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002cc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00598] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002cd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0059a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ce] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0059c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002cf] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0059e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002d0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002d1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002d2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002d3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002d4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002d5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005aa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002d6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ac] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002d7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ae] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002d8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002d9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002da] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002db] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002dc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002dd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ba] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002de] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005bc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002df] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005be] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002e0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002e1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002e2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002e3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002e4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002e5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ca] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002e6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005cc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002e7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ce] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002e8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002e9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ea] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002eb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ec] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ed] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005da] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ee] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005dc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ef] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005de] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002f0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002f1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002f2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002f3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002f4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002f5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ea] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002f6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ec] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002f7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ee] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002f8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002f9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002fa] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002fb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002fc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002fd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005fa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002fe] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005fc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h002ff] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005fe] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00300] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00600] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00301] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00602] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00302] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00604] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00303] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00606] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00304] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00608] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00305] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0060a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00306] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0060c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00307] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0060e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00308] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00610] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00309] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00612] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0030a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00614] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0030b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00616] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0030c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00618] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0030d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0061a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0030e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0061c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0030f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0061e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00310] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00620] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00311] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00622] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00312] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00624] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00313] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00626] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00314] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00628] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00315] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0062a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00316] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0062c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00317] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0062e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00318] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00630] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00319] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00632] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0031a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00634] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0031b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00636] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0031c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00638] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0031d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0063a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0031e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0063c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0031f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0063e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00320] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00640] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00321] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00642] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00322] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00644] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00323] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00646] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00324] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00648] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00325] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0064a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00326] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0064c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00327] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0064e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00328] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00650] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00329] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00652] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0032a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00654] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0032b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00656] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0032c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00658] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0032d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0065a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0032e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0065c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0032f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0065e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00330] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00660] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00331] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00662] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00332] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00664] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00333] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00666] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00334] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00668] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00335] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0066a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00336] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0066c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00337] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0066e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00338] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00670] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00339] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00672] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0033a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00674] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0033b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00676] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0033c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00678] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0033d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0067a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0033e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0067c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0033f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0067e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00340] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00680] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00341] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00682] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00342] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00684] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00343] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00686] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00344] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00688] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00345] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0068a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00346] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0068c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00347] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0068e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00348] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00690] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00349] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00692] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0034a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00694] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0034b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00696] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0034c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00698] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0034d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0069a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0034e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0069c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0034f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0069e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00350] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00351] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00352] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00353] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00354] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00355] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006aa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00356] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ac] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00357] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ae] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00358] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00359] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0035a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0035b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0035c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0035d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ba] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0035e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006bc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0035f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006be] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00360] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00361] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00362] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00363] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00364] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00365] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ca] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00366] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006cc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00367] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ce] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00368] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00369] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0036a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0036b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0036c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0036d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006da] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0036e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006dc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0036f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006de] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00370] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00371] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00372] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00373] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00374] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00375] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ea] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00376] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ec] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00377] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ee] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00378] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00379] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0037a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0037b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0037c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0037d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006fa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0037e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006fc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0037f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006fe] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00380] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00700] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00381] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00702] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00382] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00704] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00383] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00706] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00384] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00708] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00385] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0070a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00386] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0070c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00387] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0070e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00388] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00710] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00389] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00712] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0038a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00714] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0038b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00716] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0038c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00718] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0038d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0071a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0038e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0071c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0038f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0071e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00390] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00720] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00391] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00722] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00392] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00724] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00393] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00726] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00394] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00728] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00395] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0072a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00396] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0072c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00397] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0072e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00398] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00730] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h00399] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00732] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0039a] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00734] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0039b] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00736] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0039c] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00738] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0039d] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0073a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0039e] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0073c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h0039f] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0073e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003a0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00740] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003a1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00742] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003a2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00744] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003a3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00746] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003a4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00748] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003a5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0074a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003a6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0074c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003a7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0074e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003a8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00750] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003a9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00752] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003aa] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00754] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ab] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00756] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ac] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00758] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ad] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0075a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ae] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0075c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003af] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0075e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003b0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00760] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003b1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00762] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003b2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00764] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003b3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00766] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003b4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00768] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003b5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0076a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003b6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0076c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003b7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0076e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003b8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00770] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003b9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00772] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ba] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00774] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003bb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00776] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003bc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00778] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003bd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0077a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003be] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0077c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003bf] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0077e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003c0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00780] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003c1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00782] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003c2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00784] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003c3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00786] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003c4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00788] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003c5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0078a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003c6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0078c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003c7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0078e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003c8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00790] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003c9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00792] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ca] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00794] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003cb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00796] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003cc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00798] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003cd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0079a] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ce] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0079c] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003cf] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0079e] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003d0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003d1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003d2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003d3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003d4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003d5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007aa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003d6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ac] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003d7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ae] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003d8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003d9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003da] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003db] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003dc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003dd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ba] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003de] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007bc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003df] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007be] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003e0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003e1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003e2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003e3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003e4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003e5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ca] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003e6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007cc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003e7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ce] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003e8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003e9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ea] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003eb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ec] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ed] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007da] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ee] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007dc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ef] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007de] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003f0] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003f1] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003f2] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003f3] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003f4] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003f5] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ea] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003f6] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ec] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003f7] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ee] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003f8] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f0] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003f9] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f2] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003fa] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f4] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003fb] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f6] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003fc] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f8] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003fd] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007fa] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003fe] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007fc] ;
//end
//always_comb begin // 
               Icff8af1f5c3ae89ef95ed8451273154b['h003ff] =  Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007fe] ;
//end
