reg [flogtanh_WDTH -1:0] flogtanh0x00001_0, flogtanh0x00001_0_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_1, flogtanh0x00001_1_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_2, flogtanh0x00001_2_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_3, flogtanh0x00001_3_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_4, flogtanh0x00001_4_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_5, flogtanh0x00001_5_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_6, flogtanh0x00001_6_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_7, flogtanh0x00001_7_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_8, flogtanh0x00001_8_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_9, flogtanh0x00001_9_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_10, flogtanh0x00001_10_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_11, flogtanh0x00001_11_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_12, flogtanh0x00001_12_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_13, flogtanh0x00001_13_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_14, flogtanh0x00001_14_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_15, flogtanh0x00001_15_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_16, flogtanh0x00001_16_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_17, flogtanh0x00001_17_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_18, flogtanh0x00001_18_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_19, flogtanh0x00001_19_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_20, flogtanh0x00001_20_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_21, flogtanh0x00001_21_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_22, flogtanh0x00001_22_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_23, flogtanh0x00001_23_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_24, flogtanh0x00001_24_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_25, flogtanh0x00001_25_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_26, flogtanh0x00001_26_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_27, flogtanh0x00001_27_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_28, flogtanh0x00001_28_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_29, flogtanh0x00001_29_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_30, flogtanh0x00001_30_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_31, flogtanh0x00001_31_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_32, flogtanh0x00001_32_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_33, flogtanh0x00001_33_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_34, flogtanh0x00001_34_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_35, flogtanh0x00001_35_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_36, flogtanh0x00001_36_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_37, flogtanh0x00001_37_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_38, flogtanh0x00001_38_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_39, flogtanh0x00001_39_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_40, flogtanh0x00001_40_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_41, flogtanh0x00001_41_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_42, flogtanh0x00001_42_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_43, flogtanh0x00001_43_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_44, flogtanh0x00001_44_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_45, flogtanh0x00001_45_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_46, flogtanh0x00001_46_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_47, flogtanh0x00001_47_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_48, flogtanh0x00001_48_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_49, flogtanh0x00001_49_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_50, flogtanh0x00001_50_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_51, flogtanh0x00001_51_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_52, flogtanh0x00001_52_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_53, flogtanh0x00001_53_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_54, flogtanh0x00001_54_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_55, flogtanh0x00001_55_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_56, flogtanh0x00001_56_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_57, flogtanh0x00001_57_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_58, flogtanh0x00001_58_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_59, flogtanh0x00001_59_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_60, flogtanh0x00001_60_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_61, flogtanh0x00001_61_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_62, flogtanh0x00001_62_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_63, flogtanh0x00001_63_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_64, flogtanh0x00001_64_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_65, flogtanh0x00001_65_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_66, flogtanh0x00001_66_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_67, flogtanh0x00001_67_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_68, flogtanh0x00001_68_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_69, flogtanh0x00001_69_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_70, flogtanh0x00001_70_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_71, flogtanh0x00001_71_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_72, flogtanh0x00001_72_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_73, flogtanh0x00001_73_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_74, flogtanh0x00001_74_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_75, flogtanh0x00001_75_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_76, flogtanh0x00001_76_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_77, flogtanh0x00001_77_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_78, flogtanh0x00001_78_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_79, flogtanh0x00001_79_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_80, flogtanh0x00001_80_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_81, flogtanh0x00001_81_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_82, flogtanh0x00001_82_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_83, flogtanh0x00001_83_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_84, flogtanh0x00001_84_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_85, flogtanh0x00001_85_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_86, flogtanh0x00001_86_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_87, flogtanh0x00001_87_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_88, flogtanh0x00001_88_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_89, flogtanh0x00001_89_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_90, flogtanh0x00001_90_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_91, flogtanh0x00001_91_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_92, flogtanh0x00001_92_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_93, flogtanh0x00001_93_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_94, flogtanh0x00001_94_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_95, flogtanh0x00001_95_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_96, flogtanh0x00001_96_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_97, flogtanh0x00001_97_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_98, flogtanh0x00001_98_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_99, flogtanh0x00001_99_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_100, flogtanh0x00001_100_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_101, flogtanh0x00001_101_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_102, flogtanh0x00001_102_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_103, flogtanh0x00001_103_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_104, flogtanh0x00001_104_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_105, flogtanh0x00001_105_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_106, flogtanh0x00001_106_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_107, flogtanh0x00001_107_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_108, flogtanh0x00001_108_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_109, flogtanh0x00001_109_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_110, flogtanh0x00001_110_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_111, flogtanh0x00001_111_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_112, flogtanh0x00001_112_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_113, flogtanh0x00001_113_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_114, flogtanh0x00001_114_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_115, flogtanh0x00001_115_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_116, flogtanh0x00001_116_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_117, flogtanh0x00001_117_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_118, flogtanh0x00001_118_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_119, flogtanh0x00001_119_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_120, flogtanh0x00001_120_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_121, flogtanh0x00001_121_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_122, flogtanh0x00001_122_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_123, flogtanh0x00001_123_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_124, flogtanh0x00001_124_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_125, flogtanh0x00001_125_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_126, flogtanh0x00001_126_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_127, flogtanh0x00001_127_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_128, flogtanh0x00001_128_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_129, flogtanh0x00001_129_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_130, flogtanh0x00001_130_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_131, flogtanh0x00001_131_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_132, flogtanh0x00001_132_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_133, flogtanh0x00001_133_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_134, flogtanh0x00001_134_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_135, flogtanh0x00001_135_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_136, flogtanh0x00001_136_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_137, flogtanh0x00001_137_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_138, flogtanh0x00001_138_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_139, flogtanh0x00001_139_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_140, flogtanh0x00001_140_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_141, flogtanh0x00001_141_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_142, flogtanh0x00001_142_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_143, flogtanh0x00001_143_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_144, flogtanh0x00001_144_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_145, flogtanh0x00001_145_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_146, flogtanh0x00001_146_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_147, flogtanh0x00001_147_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_148, flogtanh0x00001_148_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_149, flogtanh0x00001_149_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_150, flogtanh0x00001_150_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_151, flogtanh0x00001_151_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_152, flogtanh0x00001_152_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_153, flogtanh0x00001_153_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_154, flogtanh0x00001_154_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_155, flogtanh0x00001_155_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_156, flogtanh0x00001_156_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_157, flogtanh0x00001_157_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_158, flogtanh0x00001_158_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_159, flogtanh0x00001_159_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_160, flogtanh0x00001_160_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_161, flogtanh0x00001_161_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_162, flogtanh0x00001_162_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_163, flogtanh0x00001_163_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_164, flogtanh0x00001_164_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_165, flogtanh0x00001_165_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_166, flogtanh0x00001_166_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_167, flogtanh0x00001_167_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_168, flogtanh0x00001_168_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_169, flogtanh0x00001_169_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_170, flogtanh0x00001_170_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_171, flogtanh0x00001_171_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_172, flogtanh0x00001_172_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_173, flogtanh0x00001_173_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_174, flogtanh0x00001_174_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_175, flogtanh0x00001_175_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_176, flogtanh0x00001_176_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00001_177, flogtanh0x00001_177_q;
reg start_d_flogtanh0x00001_q ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 flogtanh0x00001_0_q <= 'h0;
 flogtanh0x00001_1_q <= 'h0;
 flogtanh0x00001_2_q <= 'h0;
 flogtanh0x00001_3_q <= 'h0;
 flogtanh0x00001_4_q <= 'h0;
 flogtanh0x00001_5_q <= 'h0;
 flogtanh0x00001_6_q <= 'h0;
 flogtanh0x00001_7_q <= 'h0;
 flogtanh0x00001_8_q <= 'h0;
 flogtanh0x00001_9_q <= 'h0;
 flogtanh0x00001_10_q <= 'h0;
 flogtanh0x00001_11_q <= 'h0;
 flogtanh0x00001_12_q <= 'h0;
 flogtanh0x00001_13_q <= 'h0;
 flogtanh0x00001_14_q <= 'h0;
 flogtanh0x00001_15_q <= 'h0;
 flogtanh0x00001_16_q <= 'h0;
 flogtanh0x00001_17_q <= 'h0;
 flogtanh0x00001_18_q <= 'h0;
 flogtanh0x00001_19_q <= 'h0;
 flogtanh0x00001_20_q <= 'h0;
 flogtanh0x00001_21_q <= 'h0;
 flogtanh0x00001_22_q <= 'h0;
 flogtanh0x00001_23_q <= 'h0;
 flogtanh0x00001_24_q <= 'h0;
 flogtanh0x00001_25_q <= 'h0;
 flogtanh0x00001_26_q <= 'h0;
 flogtanh0x00001_27_q <= 'h0;
 flogtanh0x00001_28_q <= 'h0;
 flogtanh0x00001_29_q <= 'h0;
 flogtanh0x00001_30_q <= 'h0;
 flogtanh0x00001_31_q <= 'h0;
 flogtanh0x00001_32_q <= 'h0;
 flogtanh0x00001_33_q <= 'h0;
 flogtanh0x00001_34_q <= 'h0;
 flogtanh0x00001_35_q <= 'h0;
 flogtanh0x00001_36_q <= 'h0;
 flogtanh0x00001_37_q <= 'h0;
 flogtanh0x00001_38_q <= 'h0;
 flogtanh0x00001_39_q <= 'h0;
 flogtanh0x00001_40_q <= 'h0;
 flogtanh0x00001_41_q <= 'h0;
 flogtanh0x00001_42_q <= 'h0;
 flogtanh0x00001_43_q <= 'h0;
 flogtanh0x00001_44_q <= 'h0;
 flogtanh0x00001_45_q <= 'h0;
 flogtanh0x00001_46_q <= 'h0;
 flogtanh0x00001_47_q <= 'h0;
 flogtanh0x00001_48_q <= 'h0;
 flogtanh0x00001_49_q <= 'h0;
 flogtanh0x00001_50_q <= 'h0;
 flogtanh0x00001_51_q <= 'h0;
 flogtanh0x00001_52_q <= 'h0;
 flogtanh0x00001_53_q <= 'h0;
 flogtanh0x00001_54_q <= 'h0;
 flogtanh0x00001_55_q <= 'h0;
 flogtanh0x00001_56_q <= 'h0;
 flogtanh0x00001_57_q <= 'h0;
 flogtanh0x00001_58_q <= 'h0;
 flogtanh0x00001_59_q <= 'h0;
 flogtanh0x00001_60_q <= 'h0;
 flogtanh0x00001_61_q <= 'h0;
 flogtanh0x00001_62_q <= 'h0;
 flogtanh0x00001_63_q <= 'h0;
 flogtanh0x00001_64_q <= 'h0;
 flogtanh0x00001_65_q <= 'h0;
 flogtanh0x00001_66_q <= 'h0;
 flogtanh0x00001_67_q <= 'h0;
 flogtanh0x00001_68_q <= 'h0;
 flogtanh0x00001_69_q <= 'h0;
 flogtanh0x00001_70_q <= 'h0;
 flogtanh0x00001_71_q <= 'h0;
 flogtanh0x00001_72_q <= 'h0;
 flogtanh0x00001_73_q <= 'h0;
 flogtanh0x00001_74_q <= 'h0;
 flogtanh0x00001_75_q <= 'h0;
 flogtanh0x00001_76_q <= 'h0;
 flogtanh0x00001_77_q <= 'h0;
 flogtanh0x00001_78_q <= 'h0;
 flogtanh0x00001_79_q <= 'h0;
 flogtanh0x00001_80_q <= 'h0;
 flogtanh0x00001_81_q <= 'h0;
 flogtanh0x00001_82_q <= 'h0;
 flogtanh0x00001_83_q <= 'h0;
 flogtanh0x00001_84_q <= 'h0;
 flogtanh0x00001_85_q <= 'h0;
 flogtanh0x00001_86_q <= 'h0;
 flogtanh0x00001_87_q <= 'h0;
 flogtanh0x00001_88_q <= 'h0;
 flogtanh0x00001_89_q <= 'h0;
 flogtanh0x00001_90_q <= 'h0;
 flogtanh0x00001_91_q <= 'h0;
 flogtanh0x00001_92_q <= 'h0;
 flogtanh0x00001_93_q <= 'h0;
 flogtanh0x00001_94_q <= 'h0;
 flogtanh0x00001_95_q <= 'h0;
 flogtanh0x00001_96_q <= 'h0;
 flogtanh0x00001_97_q <= 'h0;
 flogtanh0x00001_98_q <= 'h0;
 flogtanh0x00001_99_q <= 'h0;
 flogtanh0x00001_100_q <= 'h0;
 flogtanh0x00001_101_q <= 'h0;
 flogtanh0x00001_102_q <= 'h0;
 flogtanh0x00001_103_q <= 'h0;
 flogtanh0x00001_104_q <= 'h0;
 flogtanh0x00001_105_q <= 'h0;
 flogtanh0x00001_106_q <= 'h0;
 flogtanh0x00001_107_q <= 'h0;
 flogtanh0x00001_108_q <= 'h0;
 flogtanh0x00001_109_q <= 'h0;
 flogtanh0x00001_110_q <= 'h0;
 flogtanh0x00001_111_q <= 'h0;
 flogtanh0x00001_112_q <= 'h0;
 flogtanh0x00001_113_q <= 'h0;
 flogtanh0x00001_114_q <= 'h0;
 flogtanh0x00001_115_q <= 'h0;
 flogtanh0x00001_116_q <= 'h0;
 flogtanh0x00001_117_q <= 'h0;
 flogtanh0x00001_118_q <= 'h0;
 flogtanh0x00001_119_q <= 'h0;
 flogtanh0x00001_120_q <= 'h0;
 flogtanh0x00001_121_q <= 'h0;
 flogtanh0x00001_122_q <= 'h0;
 flogtanh0x00001_123_q <= 'h0;
 flogtanh0x00001_124_q <= 'h0;
 flogtanh0x00001_125_q <= 'h0;
 flogtanh0x00001_126_q <= 'h0;
 flogtanh0x00001_127_q <= 'h0;
 flogtanh0x00001_128_q <= 'h0;
 flogtanh0x00001_129_q <= 'h0;
 flogtanh0x00001_130_q <= 'h0;
 flogtanh0x00001_131_q <= 'h0;
 flogtanh0x00001_132_q <= 'h0;
 flogtanh0x00001_133_q <= 'h0;
 flogtanh0x00001_134_q <= 'h0;
 flogtanh0x00001_135_q <= 'h0;
 flogtanh0x00001_136_q <= 'h0;
 flogtanh0x00001_137_q <= 'h0;
 flogtanh0x00001_138_q <= 'h0;
 flogtanh0x00001_139_q <= 'h0;
 flogtanh0x00001_140_q <= 'h0;
 flogtanh0x00001_141_q <= 'h0;
 flogtanh0x00001_142_q <= 'h0;
 flogtanh0x00001_143_q <= 'h0;
 flogtanh0x00001_144_q <= 'h0;
 flogtanh0x00001_145_q <= 'h0;
 flogtanh0x00001_146_q <= 'h0;
 flogtanh0x00001_147_q <= 'h0;
 flogtanh0x00001_148_q <= 'h0;
 flogtanh0x00001_149_q <= 'h0;
 flogtanh0x00001_150_q <= 'h0;
 flogtanh0x00001_151_q <= 'h0;
 flogtanh0x00001_152_q <= 'h0;
 flogtanh0x00001_153_q <= 'h0;
 flogtanh0x00001_154_q <= 'h0;
 flogtanh0x00001_155_q <= 'h0;
 flogtanh0x00001_156_q <= 'h0;
 flogtanh0x00001_157_q <= 'h0;
 flogtanh0x00001_158_q <= 'h0;
 flogtanh0x00001_159_q <= 'h0;
 flogtanh0x00001_160_q <= 'h0;
 flogtanh0x00001_161_q <= 'h0;
 flogtanh0x00001_162_q <= 'h0;
 flogtanh0x00001_163_q <= 'h0;
 flogtanh0x00001_164_q <= 'h0;
 flogtanh0x00001_165_q <= 'h0;
 flogtanh0x00001_166_q <= 'h0;
 flogtanh0x00001_167_q <= 'h0;
 flogtanh0x00001_168_q <= 'h0;
 flogtanh0x00001_169_q <= 'h0;
 flogtanh0x00001_170_q <= 'h0;
 flogtanh0x00001_171_q <= 'h0;
 flogtanh0x00001_172_q <= 'h0;
 flogtanh0x00001_173_q <= 'h0;
 flogtanh0x00001_174_q <= 'h0;
 flogtanh0x00001_175_q <= 'h0;
 flogtanh0x00001_176_q <= 'h0;
 flogtanh0x00001_177_q <= 'h0;
 start_d_flogtanh0x00001_q <= 'h0;
end
else
begin
 flogtanh0x00001_0_q <=  flogtanh0x00001_0;
 flogtanh0x00001_1_q <=  flogtanh0x00001_1;
 flogtanh0x00001_2_q <=  flogtanh0x00001_2;
 flogtanh0x00001_3_q <=  flogtanh0x00001_3;
 flogtanh0x00001_4_q <=  flogtanh0x00001_4;
 flogtanh0x00001_5_q <=  flogtanh0x00001_5;
 flogtanh0x00001_6_q <=  flogtanh0x00001_6;
 flogtanh0x00001_7_q <=  flogtanh0x00001_7;
 flogtanh0x00001_8_q <=  flogtanh0x00001_8;
 flogtanh0x00001_9_q <=  flogtanh0x00001_9;
 flogtanh0x00001_10_q <=  flogtanh0x00001_10;
 flogtanh0x00001_11_q <=  flogtanh0x00001_11;
 flogtanh0x00001_12_q <=  flogtanh0x00001_12;
 flogtanh0x00001_13_q <=  flogtanh0x00001_13;
 flogtanh0x00001_14_q <=  flogtanh0x00001_14;
 flogtanh0x00001_15_q <=  flogtanh0x00001_15;
 flogtanh0x00001_16_q <=  flogtanh0x00001_16;
 flogtanh0x00001_17_q <=  flogtanh0x00001_17;
 flogtanh0x00001_18_q <=  flogtanh0x00001_18;
 flogtanh0x00001_19_q <=  flogtanh0x00001_19;
 flogtanh0x00001_20_q <=  flogtanh0x00001_20;
 flogtanh0x00001_21_q <=  flogtanh0x00001_21;
 flogtanh0x00001_22_q <=  flogtanh0x00001_22;
 flogtanh0x00001_23_q <=  flogtanh0x00001_23;
 flogtanh0x00001_24_q <=  flogtanh0x00001_24;
 flogtanh0x00001_25_q <=  flogtanh0x00001_25;
 flogtanh0x00001_26_q <=  flogtanh0x00001_26;
 flogtanh0x00001_27_q <=  flogtanh0x00001_27;
 flogtanh0x00001_28_q <=  flogtanh0x00001_28;
 flogtanh0x00001_29_q <=  flogtanh0x00001_29;
 flogtanh0x00001_30_q <=  flogtanh0x00001_30;
 flogtanh0x00001_31_q <=  flogtanh0x00001_31;
 flogtanh0x00001_32_q <=  flogtanh0x00001_32;
 flogtanh0x00001_33_q <=  flogtanh0x00001_33;
 flogtanh0x00001_34_q <=  flogtanh0x00001_34;
 flogtanh0x00001_35_q <=  flogtanh0x00001_35;
 flogtanh0x00001_36_q <=  flogtanh0x00001_36;
 flogtanh0x00001_37_q <=  flogtanh0x00001_37;
 flogtanh0x00001_38_q <=  flogtanh0x00001_38;
 flogtanh0x00001_39_q <=  flogtanh0x00001_39;
 flogtanh0x00001_40_q <=  flogtanh0x00001_40;
 flogtanh0x00001_41_q <=  flogtanh0x00001_41;
 flogtanh0x00001_42_q <=  flogtanh0x00001_42;
 flogtanh0x00001_43_q <=  flogtanh0x00001_43;
 flogtanh0x00001_44_q <=  flogtanh0x00001_44;
 flogtanh0x00001_45_q <=  flogtanh0x00001_45;
 flogtanh0x00001_46_q <=  flogtanh0x00001_46;
 flogtanh0x00001_47_q <=  flogtanh0x00001_47;
 flogtanh0x00001_48_q <=  flogtanh0x00001_48;
 flogtanh0x00001_49_q <=  flogtanh0x00001_49;
 flogtanh0x00001_50_q <=  flogtanh0x00001_50;
 flogtanh0x00001_51_q <=  flogtanh0x00001_51;
 flogtanh0x00001_52_q <=  flogtanh0x00001_52;
 flogtanh0x00001_53_q <=  flogtanh0x00001_53;
 flogtanh0x00001_54_q <=  flogtanh0x00001_54;
 flogtanh0x00001_55_q <=  flogtanh0x00001_55;
 flogtanh0x00001_56_q <=  flogtanh0x00001_56;
 flogtanh0x00001_57_q <=  flogtanh0x00001_57;
 flogtanh0x00001_58_q <=  flogtanh0x00001_58;
 flogtanh0x00001_59_q <=  flogtanh0x00001_59;
 flogtanh0x00001_60_q <=  flogtanh0x00001_60;
 flogtanh0x00001_61_q <=  flogtanh0x00001_61;
 flogtanh0x00001_62_q <=  flogtanh0x00001_62;
 flogtanh0x00001_63_q <=  flogtanh0x00001_63;
 flogtanh0x00001_64_q <=  flogtanh0x00001_64;
 flogtanh0x00001_65_q <=  flogtanh0x00001_65;
 flogtanh0x00001_66_q <=  flogtanh0x00001_66;
 flogtanh0x00001_67_q <=  flogtanh0x00001_67;
 flogtanh0x00001_68_q <=  flogtanh0x00001_68;
 flogtanh0x00001_69_q <=  flogtanh0x00001_69;
 flogtanh0x00001_70_q <=  flogtanh0x00001_70;
 flogtanh0x00001_71_q <=  flogtanh0x00001_71;
 flogtanh0x00001_72_q <=  flogtanh0x00001_72;
 flogtanh0x00001_73_q <=  flogtanh0x00001_73;
 flogtanh0x00001_74_q <=  flogtanh0x00001_74;
 flogtanh0x00001_75_q <=  flogtanh0x00001_75;
 flogtanh0x00001_76_q <=  flogtanh0x00001_76;
 flogtanh0x00001_77_q <=  flogtanh0x00001_77;
 flogtanh0x00001_78_q <=  flogtanh0x00001_78;
 flogtanh0x00001_79_q <=  flogtanh0x00001_79;
 flogtanh0x00001_80_q <=  flogtanh0x00001_80;
 flogtanh0x00001_81_q <=  flogtanh0x00001_81;
 flogtanh0x00001_82_q <=  flogtanh0x00001_82;
 flogtanh0x00001_83_q <=  flogtanh0x00001_83;
 flogtanh0x00001_84_q <=  flogtanh0x00001_84;
 flogtanh0x00001_85_q <=  flogtanh0x00001_85;
 flogtanh0x00001_86_q <=  flogtanh0x00001_86;
 flogtanh0x00001_87_q <=  flogtanh0x00001_87;
 flogtanh0x00001_88_q <=  flogtanh0x00001_88;
 flogtanh0x00001_89_q <=  flogtanh0x00001_89;
 flogtanh0x00001_90_q <=  flogtanh0x00001_90;
 flogtanh0x00001_91_q <=  flogtanh0x00001_91;
 flogtanh0x00001_92_q <=  flogtanh0x00001_92;
 flogtanh0x00001_93_q <=  flogtanh0x00001_93;
 flogtanh0x00001_94_q <=  flogtanh0x00001_94;
 flogtanh0x00001_95_q <=  flogtanh0x00001_95;
 flogtanh0x00001_96_q <=  flogtanh0x00001_96;
 flogtanh0x00001_97_q <=  flogtanh0x00001_97;
 flogtanh0x00001_98_q <=  flogtanh0x00001_98;
 flogtanh0x00001_99_q <=  flogtanh0x00001_99;
 flogtanh0x00001_100_q <=  flogtanh0x00001_100;
 flogtanh0x00001_101_q <=  flogtanh0x00001_101;
 flogtanh0x00001_102_q <=  flogtanh0x00001_102;
 flogtanh0x00001_103_q <=  flogtanh0x00001_103;
 flogtanh0x00001_104_q <=  flogtanh0x00001_104;
 flogtanh0x00001_105_q <=  flogtanh0x00001_105;
 flogtanh0x00001_106_q <=  flogtanh0x00001_106;
 flogtanh0x00001_107_q <=  flogtanh0x00001_107;
 flogtanh0x00001_108_q <=  flogtanh0x00001_108;
 flogtanh0x00001_109_q <=  flogtanh0x00001_109;
 flogtanh0x00001_110_q <=  flogtanh0x00001_110;
 flogtanh0x00001_111_q <=  flogtanh0x00001_111;
 flogtanh0x00001_112_q <=  flogtanh0x00001_112;
 flogtanh0x00001_113_q <=  flogtanh0x00001_113;
 flogtanh0x00001_114_q <=  flogtanh0x00001_114;
 flogtanh0x00001_115_q <=  flogtanh0x00001_115;
 flogtanh0x00001_116_q <=  flogtanh0x00001_116;
 flogtanh0x00001_117_q <=  flogtanh0x00001_117;
 flogtanh0x00001_118_q <=  flogtanh0x00001_118;
 flogtanh0x00001_119_q <=  flogtanh0x00001_119;
 flogtanh0x00001_120_q <=  flogtanh0x00001_120;
 flogtanh0x00001_121_q <=  flogtanh0x00001_121;
 flogtanh0x00001_122_q <=  flogtanh0x00001_122;
 flogtanh0x00001_123_q <=  flogtanh0x00001_123;
 flogtanh0x00001_124_q <=  flogtanh0x00001_124;
 flogtanh0x00001_125_q <=  flogtanh0x00001_125;
 flogtanh0x00001_126_q <=  flogtanh0x00001_126;
 flogtanh0x00001_127_q <=  flogtanh0x00001_127;
 flogtanh0x00001_128_q <=  flogtanh0x00001_128;
 flogtanh0x00001_129_q <=  flogtanh0x00001_129;
 flogtanh0x00001_130_q <=  flogtanh0x00001_130;
 flogtanh0x00001_131_q <=  flogtanh0x00001_131;
 flogtanh0x00001_132_q <=  flogtanh0x00001_132;
 flogtanh0x00001_133_q <=  flogtanh0x00001_133;
 flogtanh0x00001_134_q <=  flogtanh0x00001_134;
 flogtanh0x00001_135_q <=  flogtanh0x00001_135;
 flogtanh0x00001_136_q <=  flogtanh0x00001_136;
 flogtanh0x00001_137_q <=  flogtanh0x00001_137;
 flogtanh0x00001_138_q <=  flogtanh0x00001_138;
 flogtanh0x00001_139_q <=  flogtanh0x00001_139;
 flogtanh0x00001_140_q <=  flogtanh0x00001_140;
 flogtanh0x00001_141_q <=  flogtanh0x00001_141;
 flogtanh0x00001_142_q <=  flogtanh0x00001_142;
 flogtanh0x00001_143_q <=  flogtanh0x00001_143;
 flogtanh0x00001_144_q <=  flogtanh0x00001_144;
 flogtanh0x00001_145_q <=  flogtanh0x00001_145;
 flogtanh0x00001_146_q <=  flogtanh0x00001_146;
 flogtanh0x00001_147_q <=  flogtanh0x00001_147;
 flogtanh0x00001_148_q <=  flogtanh0x00001_148;
 flogtanh0x00001_149_q <=  flogtanh0x00001_149;
 flogtanh0x00001_150_q <=  flogtanh0x00001_150;
 flogtanh0x00001_151_q <=  flogtanh0x00001_151;
 flogtanh0x00001_152_q <=  flogtanh0x00001_152;
 flogtanh0x00001_153_q <=  flogtanh0x00001_153;
 flogtanh0x00001_154_q <=  flogtanh0x00001_154;
 flogtanh0x00001_155_q <=  flogtanh0x00001_155;
 flogtanh0x00001_156_q <=  flogtanh0x00001_156;
 flogtanh0x00001_157_q <=  flogtanh0x00001_157;
 flogtanh0x00001_158_q <=  flogtanh0x00001_158;
 flogtanh0x00001_159_q <=  flogtanh0x00001_159;
 flogtanh0x00001_160_q <=  flogtanh0x00001_160;
 flogtanh0x00001_161_q <=  flogtanh0x00001_161;
 flogtanh0x00001_162_q <=  flogtanh0x00001_162;
 flogtanh0x00001_163_q <=  flogtanh0x00001_163;
 flogtanh0x00001_164_q <=  flogtanh0x00001_164;
 flogtanh0x00001_165_q <=  flogtanh0x00001_165;
 flogtanh0x00001_166_q <=  flogtanh0x00001_166;
 flogtanh0x00001_167_q <=  flogtanh0x00001_167;
 flogtanh0x00001_168_q <=  flogtanh0x00001_168;
 flogtanh0x00001_169_q <=  flogtanh0x00001_169;
 flogtanh0x00001_170_q <=  flogtanh0x00001_170;
 flogtanh0x00001_171_q <=  flogtanh0x00001_171;
 flogtanh0x00001_172_q <=  flogtanh0x00001_172;
 flogtanh0x00001_173_q <=  flogtanh0x00001_173;
 flogtanh0x00001_174_q <=  flogtanh0x00001_174;
 flogtanh0x00001_175_q <=  flogtanh0x00001_175;
 flogtanh0x00001_176_q <=  flogtanh0x00001_176;
 flogtanh0x00001_177_q <=  flogtanh0x00001_177;
 start_d_flogtanh0x00001_q <=  start_d_flogtanh0x00000_q;
end
