//`include "GF2_LDPC_flogtanh_0x0000d_assign_inc.sv"
//always_comb begin
              If72de6675c42172560d5d150642f3da8['h00000] = 
          (!flogtanh_sel['h0000d]) ? 
                       Ie4acdb20b1de9050267f708a13a337e0['h00000] : //%
                       Ie4acdb20b1de9050267f708a13a337e0['h00001] ;
//end
//always_comb begin
              If72de6675c42172560d5d150642f3da8['h00001] = 
          (!flogtanh_sel['h0000d]) ? 
                       Ie4acdb20b1de9050267f708a13a337e0['h00002] : //%
                       Ie4acdb20b1de9050267f708a13a337e0['h00003] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00002] =  Ie4acdb20b1de9050267f708a13a337e0['h00004] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00003] =  Ie4acdb20b1de9050267f708a13a337e0['h00006] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00004] =  Ie4acdb20b1de9050267f708a13a337e0['h00008] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00005] =  Ie4acdb20b1de9050267f708a13a337e0['h0000a] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00006] =  Ie4acdb20b1de9050267f708a13a337e0['h0000c] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00007] =  Ie4acdb20b1de9050267f708a13a337e0['h0000e] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00008] =  Ie4acdb20b1de9050267f708a13a337e0['h00010] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00009] =  Ie4acdb20b1de9050267f708a13a337e0['h00012] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0000a] =  Ie4acdb20b1de9050267f708a13a337e0['h00014] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0000b] =  Ie4acdb20b1de9050267f708a13a337e0['h00016] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0000c] =  Ie4acdb20b1de9050267f708a13a337e0['h00018] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0000d] =  Ie4acdb20b1de9050267f708a13a337e0['h0001a] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0000e] =  Ie4acdb20b1de9050267f708a13a337e0['h0001c] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0000f] =  Ie4acdb20b1de9050267f708a13a337e0['h0001e] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00010] =  Ie4acdb20b1de9050267f708a13a337e0['h00020] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00011] =  Ie4acdb20b1de9050267f708a13a337e0['h00022] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00012] =  Ie4acdb20b1de9050267f708a13a337e0['h00024] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00013] =  Ie4acdb20b1de9050267f708a13a337e0['h00026] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00014] =  Ie4acdb20b1de9050267f708a13a337e0['h00028] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00015] =  Ie4acdb20b1de9050267f708a13a337e0['h0002a] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00016] =  Ie4acdb20b1de9050267f708a13a337e0['h0002c] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00017] =  Ie4acdb20b1de9050267f708a13a337e0['h0002e] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00018] =  Ie4acdb20b1de9050267f708a13a337e0['h00030] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h00019] =  Ie4acdb20b1de9050267f708a13a337e0['h00032] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0001a] =  Ie4acdb20b1de9050267f708a13a337e0['h00034] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0001b] =  Ie4acdb20b1de9050267f708a13a337e0['h00036] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0001c] =  Ie4acdb20b1de9050267f708a13a337e0['h00038] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0001d] =  Ie4acdb20b1de9050267f708a13a337e0['h0003a] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0001e] =  Ie4acdb20b1de9050267f708a13a337e0['h0003c] ;
//end
//always_comb begin // 
               If72de6675c42172560d5d150642f3da8['h0001f] =  Ie4acdb20b1de9050267f708a13a337e0['h0003e] ;
//end
