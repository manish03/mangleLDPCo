              I85e2d7a9e28f224cac9188370cccc37b = 
          (!flogtanh_sel[1]) ? 
                       I6ceb8a53497c625c878b1bd0b10147d1: 
                       Iebd6f893703430ccce739c17a091180a;
              I17540db3c63ade2b53e82ca752a6cd99 = 
          (!flogtanh_sel[1]) ? 
                       I87206f7a8f80c6791355b9e35fa789d4: 
                       Ibeedd439ada9e1204f23f8b4c59d160e;
              I43b24a45247c83d2a986a6e352e7a38a = 
          (!flogtanh_sel[1]) ? 
                       I722b96e8bbdedcbbf709b7ff75a343f2: 
                       Id82ca4ddd6bd7bd3eba9321f61fc83b1;
              I92680f7db736ef5df4e81244ffcff59b = 
          (!flogtanh_sel[1]) ? 
                       I2cf927aba0ba024e37641e82687e3134: 
                       I0495eb40055242fe8d9886724a00437b;
              I39764779466097d56a3a65718704d030 = 
          (!flogtanh_sel[1]) ? 
                       Iaabf9a9cb8e18da9c94d145c54613499: 
                       I9de00fb5f405754b7af66ab5206ee12c;
              I1e7b702101a2cb5064b151835830a57d = 
          (!flogtanh_sel[1]) ? 
                       I8f63c4af862af47948080677b089cc32: 
                       Iec915d0edfe90c0a3889228715277570;
              I57b599739f81aba00c5a7aa795ea08c8 = 
          (!flogtanh_sel[1]) ? 
                       I79f6ccccd78a7701f6302aab4293286c: 
                       I90fe152dd5144845dd3b473f4cafb74e;
              Ied56219095ff64722213c69d58e6b74f = 
          (!flogtanh_sel[1]) ? 
                       I0bab994e09bb74cd97afe36943a98690: 
                       Ic806ded37e428ee89a5725a3f0c69632;
              I5fbce88eb0e5add5adc151439b070eff = 
          (!flogtanh_sel[1]) ? 
                       I1bb8a779c4c359bfc508d95a8d99c676: 
                       Ic7037aee76219d7437fb16a34cd0575b;
              Ibaf106dee88a6d70caa3ca247be96938 = 
          (!flogtanh_sel[1]) ? 
                       I31653f719f0514a1e8b4dc749fa89eab: 
                       Iee53e3dc893e03efc0d4f8b9e165a5df;
              I47decd52e0f93d6281011a92a9a7081e = 
          (!flogtanh_sel[1]) ? 
                       I12f3e3785de1cf141ea2c3efa11b6323: 
                       I415f363f69a1088c765e22738019ec87;
              I4b74e2c1db97dcec11a65b57b1035acf = 
          (!flogtanh_sel[1]) ? 
                       I3e72d56a69d40deafd501605f0257ac0: 
                       I6529b2ba884c7977f550cf3410db444d;
              Ib8190cccfd6f5afb2b6cef33e5376d19 = 
          (!flogtanh_sel[1]) ? 
                       If14fba2b2f70d2602b88ff0e739e113e: 
                       I0685af82b58f41fa65efe1125fdaabeb;
              Icbc0f6167d607f74c80c23a3257cd2e1 = 
          (!flogtanh_sel[1]) ? 
                       I1ad44f9d9abb2121b183a93dd1af4fa5: 
                       I0f9dbc9aa169f7d63cc5789cb75c3a2d;
              Ieac93250ec9be2ef318d48baf88b1ef5 = 
          (!flogtanh_sel[1]) ? 
                       I5e458356e7698884ee785b2d5f1c368a: 
                       I9b0f07f47267e3b0e0c545f44f5dd9f9;
              I5db1844e769af7943f93da66b475d99e = 
          (!flogtanh_sel[1]) ? 
                       I3a4dd73e8b3f48746a991573531315dd: 
                       If727e9507d63727b0d597e9a5fee202a;
              I8f242f17610cae369dbfb2aaa0453b79 = 
          (!flogtanh_sel[1]) ? 
                       I9253bbcea2dc3a74433955d5f5aff705: 
                       Ibbabd657d00fc10d293b680d89593ca7;
              I5bebf7ec46791bfa6d1dad7eceeea034 = 
          (!flogtanh_sel[1]) ? 
                       I79b7daae3f9f65acd3f79d579d2af25a: 
                       I74a4a1e449670380db8fbedbcf2aec04;
              Ife8a533289756df000f25a54a51bcfe3 = 
          (!flogtanh_sel[1]) ? 
                       I9f7da2708edf4c941682b24f3999b159: 
                       Id5d585b0c590354af34d02ba320f80d9;
              I5de464a27ad96e1c636efd974f129cfe = 
          (!flogtanh_sel[1]) ? 
                       Idab5b4bb4ed70dfe122f645eaf32852c: 
                       Ic1793b6e075a12f6c1dda7e9fddc8b6e;
              I5f1b79389154a01c7d846f5f8774dfa7 = 
          (!flogtanh_sel[1]) ? 
                       I168c51768b35b16f0033808f0b915e8c: 
                       Ia7fa2fefde3f2ad6a0bee771a131219b;
              If3d70b7c1e8f802b887c01e068428a4e = 
          (!flogtanh_sel[1]) ? 
                       I22d2ffb044bf579a2cccd3fcc70dae45: 
                       Ib4b3cd8d5376f6ddb653c8cf72dceabf;
              Ic10bc44ab0b4ca1d588d768859f1bb35 = 
          (!flogtanh_sel[1]) ? 
                       I2c0b6e7a1fbcd97b6b78e65bf6d61213: 
                       Ifabbe9c31875e40eb81a87f0b19134e5;
              Ie3cd02462472a4430da14641cda50452 = 
          (!flogtanh_sel[1]) ? 
                       Ic20259ce7eabae2029ca2ce312c6bfed: 
                       Icaf0213b02a3cad251718b9ff86c108b;
              I3071dd54b8e3e01163a9d17df901a502 = 
          (!flogtanh_sel[1]) ? 
                       If71ff543c013f0111318a06039267570: 
                       I7871649505392bea882ad24b821c953c;
              I7fa902c92592761b9689aec509e9e68f = 
          (!flogtanh_sel[1]) ? 
                       I5c4bcb5584cd15cbbec2709f29e15f36: 
                       I73b98efd2185919a61b91a641fd6bdd7;
              I13ac2bb6eb27b06cc93e19bec590ac44 = 
          (!flogtanh_sel[1]) ? 
                       Ic2519d8c4e9b2c6f2126407a7a39fefe: 
                       Ia806cdd7fbd6b44a8256aee7250ddd8b;
              Ied47c387d2e31433fbd752243e5e0aac = 
          (!flogtanh_sel[1]) ? 
                       I9badff60aa84397c6a408b846feceb91: 
                       I885c54956c3ff7dfcd971f9d7ddf2db1;
              I470d7fc38fd4e1b015a43ce4f898f2bd = 
          (!flogtanh_sel[1]) ? 
                       Ie3ae98a6abd28a3c39863a981e88e63f: 
                       Ia1fed14f941d2ef3e78c490f81a5bd04;
              If1f7c2655f45c9148824e4151ab448b6 = 
          (!flogtanh_sel[1]) ? 
                       I714c5a8ac1480b08aa2859680ae40660: 
                       I11d5e654536cd6b6e9b91487d76facb6;
              If120a179bc9b785016b64084d6e4d056 = 
          (!flogtanh_sel[1]) ? 
                       I32f53cb8d864ff40c8d0ef95e9bdde54: 
                       I0c3874311a119530873f475b01006dd4;
              I7fc7f688e30263828dfdaf9ec8ec2f7a = 
          (!flogtanh_sel[1]) ? 
                       I585684cf3ba45f359e0f0752e9e88819: 
                       I998f8a35c7ec923067dc75c76c9df713;
               Ia8804339708717f01d9a9069c72f0fbb =  I4e8f27bdc42f1e3f4024b020d5821dff ;
               I5079e19864882aa577c73731fcee0a31 =  I9ae8e176f8f34220d2cac97abe1fd32a ;
               Ia0dceddb9355f13a3a622f279c244f06 =  Ic9bc7816fcb1f128d833fde39ad8cf1d ;
               I75a27f997d71f89b8beb0484ec0402d5 =  I3479e7931017ab45aa4e99ca34b8b5cb ;
              I6557d5a7415612889373a46ee77437c5 = 
          (!flogtanh_sel[1]) ? 
                       I32769b7f105065785745633dfef8a4c5: 
                       I47e2d27cbd69c85106a4aa3ac2784eb0;
              Ieef6c1b5a0ec168747b3dedc3f88e803 = 
          (!flogtanh_sel[1]) ? 
                       Ibd0efa281371fa3b94eed5e021c73642: 
                       I82aaeb65a83948cd75521499d2719001;
              I892de6b0f85b4aea7ff9113d713552e2 = 
          (!flogtanh_sel[1]) ? 
                       If9854de536b8ba1392ba0328ef7cebba: 
                       I731416642a03748ca4698a73e094c500;
               Ie8c260c1c1a61ba194c563e25325b435 =  I23c90590a514d430c9828af570ebf16a ;
              Ic34456cc9dc2004ffb6ac0974c98e0e4 = 
          (!flogtanh_sel[1]) ? 
                       I89fc8a2a491dcc20f2556e7042d22384: 
                       I0f76a71ea70551bbf89f01a689811954;
              I59e956b7f374eed213b25d05b702aa7b = 
          (!flogtanh_sel[1]) ? 
                       I0b6ce8e59afb2e48df79fefd5450971e: 
                       I35a8c09862db36ffde26d27b74baa8ba;
               I3f03c8fa63d838b3d42c3f047e70fbf5 =  I920593851f5860485fd105f8d4c1b8c9 ;
              I3d899ecab223931d4c0e12833417e32b = 
          (!flogtanh_sel[1]) ? 
                       I79489994f40f88e0b5a8a8be6322f3ec: 
                       I6503341e5d6ced0d71bd29bbc622020b;
               I1c56ccfd13ce759046362280dce3ef9c =  I178d103fabf53395ce88cdbfc14917ce ;
              Icc0a9c979d7e154edb892315a4ca9cfd = 
          (!flogtanh_sel[1]) ? 
                       I4602a0caf02e37e360e5cf9de1003cd2: 
                       I245a6df9f9d730338cd52169a3f466d3;
               Ieac7270ea1f936fea6df9fa9233a78a1 =  Ia7a8ebe681523a490c83dcb84ac82a2a ;
              Id9a98abcca5f5bf46e2dce45066d2dd6 = 
          (!flogtanh_sel[1]) ? 
                       I401eb53331986f8474c861acb2b2a445: 
                       If3e4f18a03ca4b7b1d89ef842c68e96d;
               I240fa7efcb0d0196b865a47048e9f5e2 =  I0d6bc03eddef33a7d70ac2cc27049107 ;
               I83a9fc44b887c9b860d07ba9d9a90083 =  I6138bf9b2a35f3b08f216eeaf3c0ebee ;
              Ic20207f1d7c0f19dba8676141ca07549 = 
          (!flogtanh_sel[1]) ? 
                       I26faa75fc5dd15baf23481311b220832: 
                       I373328eb3cc59c5d3d7a5102535c5410;
               Ic4c14384ec86a331d36974bb41903efa =  I1bb3c77cdfd0b229bbdf7b33fd4a613c ;
               I87fab4038ff6c1bc1bcc170f9a202769 =  Ib911176056f3c0378dfa8a77e0c5b69a ;
              I47e00ea6506dbd4a360baf94cf63dc2a = 
          (!flogtanh_sel[1]) ? 
                       I6bb576223350a8373e430d185efe7fd9: 
                       Id7008a8f0d70f1e23a073745ed4a57c0;
               Ia2683d4666dbf6b9f8befa2d6bdbbfcb =  I87e0bcba46bcc28ad02b7e0af773d82a ;
               I1ed7dd07abe9aee415671c6222bdc16c =  Iea2bbf25e38901d15434dfc83d65ada4 ;
               I5ea7cfba8e7720077757862cf36ceaa2 =  Ibcc6c8744ee9a2ad9766c0f9fa196036 ;
              Ifb1ba203c0ec3fc5e1081393bf492c20 = 
          (!flogtanh_sel[1]) ? 
                       I78ba7a5627868f3c0b75555131470aa4: 
                       I3b5bd630c8d2bdb455b6f75a6a8a4a53;
               Id0417686b69b456644d09aaa861f26d4 =  I4274a587dd459b29ecee1ff1554a12f7 ;
               I4c3cbe58c98f3e0fdf9c89b7143e50a3 =  If77d0921ff0a38d2b3fcd28c5be4a131 ;
               I0915e1427b7e3267e7ffe79d0cc782f3 =  I6fbdabe9ecefa8648c4ca4ec51e251a4 ;
               Id5a895fa3677c1f973675aebec6b41f2 =  Ib68b82bab62a694692b3fd2191b5f29c ;
               I023b610b050357cc816939b6508bedb9 =  Id5c5e697446d9974b383880138f73778 ;
               Ia7f89e3fc13d2589f1a2a025830a8b9e =  Ic117c98ae21f7640aa5a68539ec03821 ;
               I51c00546226c98d468b69a85d8613b4d =  Idc31f916f132a0c203eb03a7d1de62bb ;
               Ie5f68f657e8123b2e971d4f3e5a675df =  I5e4276800e079f48c3953f01869bcfa0 ;
               Ia9194d615d26094f0c3e0399ab2e3da3 =  I5955344e0f04e1ddf15eecf2eede2346 ;
               I9f1ef03445a07c36defabb3abd5df4c4 =  I83df9b9b4dc9b0eeaf05f25e513d1603 ;
               I8f90fcb8534f00216e0f6c4a3dbad2f6 =  I5b3e2ec3e81cfbb4cff4a55faf1779ce ;
               I30166adbb988446bdb36723a2e4cd7c1 =  Iecc3e2589b1a21ad89360386cbc59203 ;
               Ief50b2820a6d32e602d4963c13b3f630 =  Ibce5b55e9f3477e8cac134660f3e056d ;
              If51760e69ff89f244fdb9cdb0b93bda4 = 
          (!flogtanh_sel[1]) ? 
                       Ic95be5fcb699a68e0e796dc0408fd5f3: 
                       I01c4e6856aaa370540e370d30223a3e9;
               Idf43504868969d00511ef6e8d809db66 =  I693343088a46766b65b21833e8c93424 ;
               Icfc6c999050d945d3a381ba869dd6e76 =  Ibcd20a65390727b99272e778f6b5cd48 ;
               Iec57a1e76f07f3c328f74bfe5b1da785 =  Iee99e323224f79b59ff094ca4e0b730f ;
               Ice973d37ca9816e4e5b7221463d76636 =  Icf2d8147505a677d965332527efd32e5 ;
               I87c9f04f74686c1dee6305deb51b9007 =  I7af4f3f04f52198149fab343b09a7c33 ;
               I9350b76d99dd94589a9997500354f19d =  I8d3688317aaf1a973e53e7d82c07aff5 ;
               Idd0acb6b0bc3d9e3a12715d4f6614149 =  I2145db99a9f07a8dcca7bb21537c3c6b ;
               Idab3e6bf2379a457d67cce07ca31ba57 =  Ia36d890f9c568613260b96683ad1442e ;
               Ie2f28a6c2445f5178eecc13507b72323 =  I83e8203369eabb1165454d054fc6368a ;
               I5d3b6f0d046829b096807ab4a49bcc25 =  I2cf7c8df11a71a3952a5c11fce1ab746 ;
               I0b3c995b0a12a14265de007d90300cec =  I964950b31cf4117e79e46a2282faf273 ;
               I31b53846b721e11cddea32c4b046a7fa =  I754ed93d8e7f3ed1b9bbf1aa0a780631 ;
               I1b40caccc7bf0db9618dd54d2959ee2a =  I0be6033ae52cefc976cf28e9c6972b2c ;
               I832959dc65f560a892c99dc05dfb19ff =  I332be99f2c509a0ad9ce2003f3894900 ;
               I515dd393df02b089c3afa5ef912c945a =  Ic98c3c04426af7540b59e85693f8c85e ;
               I55b2317ed99a99a1afd11aff3c296683 =  Ie34547c669ac94c6b215f01c235086e4 ;
              I8122943006aece7452a503e8c20375b4 = 
          (!flogtanh_sel[1]) ? 
                       I27def56001fb56e6a85c9c61ba8d55bd: 
                       I6540e74c5f9178782a17fe7460aaf4ee;
               Ida9814058169631dca9f83ee34741a75 =  0;
