 reg  ['hffff:0] [$clog2('h7000+1)-1:0] Idce7a2deb0c98f08daec6108083a2c7f ;
