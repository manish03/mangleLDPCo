//`include "GF2_LDPC_fgallag_0x00004_assign_inc.sv"
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00000] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00000] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00001] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00001] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00002] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00003] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00002] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00004] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00005] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00003] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00006] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00007] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00004] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00008] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00009] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00005] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0000a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0000b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00006] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0000c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0000d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00007] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0000e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0000f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00008] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00010] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00011] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00009] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00012] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00013] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0000a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00014] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00015] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0000b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00016] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00017] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0000c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00018] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00019] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0000d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0001a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0001b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0000e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0001c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0001d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0000f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0001e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0001f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00010] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00020] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00021] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00011] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00022] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00023] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00012] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00024] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00025] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00013] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00026] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00027] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00014] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00028] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00029] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00015] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0002a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0002b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00016] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0002c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0002d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00017] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0002e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0002f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00018] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00030] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00031] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00019] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00032] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00033] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0001a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00034] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00035] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0001b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00036] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00037] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0001c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00038] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00039] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0001d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0003a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0003b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0001e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0003c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0003d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0001f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0003e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0003f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00020] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00040] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00041] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00021] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00042] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00043] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00022] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00044] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00045] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00023] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00046] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00047] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00024] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00048] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00049] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00025] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0004a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0004b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00026] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0004c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0004d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00027] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0004e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0004f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00028] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00050] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00051] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00029] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00052] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00053] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0002a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00054] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00055] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0002b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00056] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00057] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0002c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00058] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00059] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0002d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0005a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0005b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0002e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0005c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0005d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0002f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0005e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0005f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00030] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00060] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00061] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00031] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00062] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00063] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00032] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00064] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00065] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00033] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00066] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00067] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00034] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00068] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00069] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00035] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0006a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0006b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00036] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0006c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0006d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00037] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0006e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0006f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00038] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00070] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00071] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00039] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00072] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00073] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0003a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00074] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00075] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0003b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00076] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00077] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0003c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00078] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00079] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0003d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0007a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0007b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0003e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0007c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0007d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0003f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0007e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0007f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00040] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00080] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00081] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00041] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00082] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00083] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00042] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00084] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00085] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00043] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00086] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00087] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00044] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00088] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00089] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00045] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0008a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0008b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00046] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0008c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0008d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00047] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0008e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0008f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00048] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00090] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00091] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00049] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00092] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00093] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0004a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00094] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00095] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0004b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00096] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00097] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0004c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00098] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00099] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0004d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0009a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0009b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0004e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0009c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0009d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0004f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0009e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0009f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00050] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000a0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000a1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00051] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000a2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000a3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00052] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000a4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000a5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00053] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000a6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000a7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00054] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000a8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000a9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00055] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000aa] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ab] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00056] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ac] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ad] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00057] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ae] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000af] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00058] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000b0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000b1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00059] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000b2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000b3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0005a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000b4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000b5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0005b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000b6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000b7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0005c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000b8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000b9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0005d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ba] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000bb] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0005e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000bc] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000bd] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0005f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000be] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000bf] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00060] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000c0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000c1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00061] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000c2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000c3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00062] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000c4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000c5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00063] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000c6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000c7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00064] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000c8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000c9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00065] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ca] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000cb] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00066] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000cc] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000cd] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00067] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ce] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000cf] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00068] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000d0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000d1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00069] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000d2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000d3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0006a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000d4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000d5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0006b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000d6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000d7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0006c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000d8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000d9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0006d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000da] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000db] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0006e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000dc] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000dd] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0006f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000de] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000df] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00070] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000e0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000e1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00071] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000e2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000e3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00072] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000e4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000e5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00073] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000e6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000e7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00074] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000e8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000e9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00075] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ea] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000eb] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00076] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ec] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ed] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00077] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ee] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ef] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00078] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000f0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000f1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00079] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000f2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000f3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0007a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000f4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000f5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0007b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000f6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000f7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0007c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000f8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000f9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0007d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000fa] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000fb] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0007e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000fc] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000fd] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0007f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000fe] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h000ff] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00080] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00100] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00101] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00081] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00102] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00103] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00082] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00104] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00105] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00083] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00106] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00107] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00084] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00108] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00109] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00085] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0010a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0010b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00086] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0010c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0010d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00087] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0010e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0010f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00088] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00110] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00111] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00089] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00112] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00113] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0008a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00114] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00115] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0008b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00116] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00117] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0008c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00118] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00119] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0008d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0011a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0011b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0008e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0011c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0011d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0008f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0011e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0011f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00090] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00120] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00121] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00091] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00122] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00123] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00092] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00124] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00125] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00093] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00126] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00127] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00094] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00128] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00129] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00095] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0012a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0012b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00096] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0012c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0012d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00097] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0012e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0012f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00098] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00130] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00131] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00099] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00132] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00133] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0009a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00134] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00135] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0009b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00136] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00137] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0009c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00138] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00139] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0009d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0013a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0013b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0009e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0013c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0013d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0009f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0013e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0013f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000a0] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00140] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00141] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000a1] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00142] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00143] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000a2] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00144] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00145] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000a3] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00146] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00147] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000a4] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00148] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00149] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000a5] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0014a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0014b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000a6] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0014c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0014d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000a7] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0014e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0014f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000a8] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00150] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00151] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000a9] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00152] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00153] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000aa] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00154] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00155] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ab] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00156] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00157] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ac] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00158] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00159] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ad] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0015a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0015b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ae] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0015c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0015d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000af] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0015e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0015f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000b0] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00160] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00161] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000b1] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00162] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00163] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000b2] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00164] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00165] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000b3] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00166] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00167] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000b4] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00168] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00169] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000b5] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0016a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0016b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000b6] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0016c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0016d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000b7] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0016e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0016f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000b8] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00170] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00171] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000b9] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00172] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00173] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ba] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00174] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00175] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000bb] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00176] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00177] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000bc] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00178] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00179] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000bd] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0017a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0017b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000be] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0017c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0017d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000bf] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0017e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0017f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000c0] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00180] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00181] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000c1] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00182] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00183] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000c2] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00184] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00185] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000c3] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00186] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00187] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000c4] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00188] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00189] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000c5] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0018a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0018b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000c6] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0018c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0018d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000c7] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0018e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0018f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000c8] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00190] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00191] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000c9] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00192] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00193] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ca] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00194] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00195] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000cb] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00196] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00197] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000cc] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00198] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00199] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000cd] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0019a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0019b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ce] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0019c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0019d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000cf] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0019e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0019f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000d0] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001a0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001a1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000d1] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001a2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001a3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000d2] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001a4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001a5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000d3] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001a6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001a7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000d4] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001a8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001a9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000d5] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001aa] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ab] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000d6] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ac] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ad] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000d7] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ae] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001af] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000d8] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001b0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001b1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000d9] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001b2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001b3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000da] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001b4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001b5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000db] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001b6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001b7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000dc] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001b8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001b9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000dd] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ba] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001bb] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000de] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001bc] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001bd] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000df] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001be] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001bf] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000e0] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001c0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001c1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000e1] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001c2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001c3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000e2] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001c4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001c5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000e3] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001c6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001c7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000e4] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001c8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001c9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000e5] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ca] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001cb] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000e6] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001cc] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001cd] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000e7] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ce] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001cf] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000e8] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001d0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001d1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000e9] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001d2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001d3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ea] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001d4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001d5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000eb] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001d6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001d7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ec] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001d8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001d9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ed] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001da] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001db] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ee] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001dc] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001dd] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ef] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001de] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001df] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000f0] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001e0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001e1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000f1] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001e2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001e3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000f2] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001e4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001e5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000f3] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001e6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001e7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000f4] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001e8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001e9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000f5] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ea] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001eb] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000f6] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ec] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ed] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000f7] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ee] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ef] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000f8] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001f0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001f1] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000f9] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001f2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001f3] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000fa] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001f4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001f5] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000fb] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001f6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001f7] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000fc] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001f8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001f9] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000fd] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001fa] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001fb] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000fe] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001fc] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001fd] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h000ff] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001fe] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h001ff] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00100] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00200] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00201] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00101] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00202] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00203] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00102] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00204] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00205] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00103] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00206] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00207] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00104] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00208] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00209] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00105] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0020a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0020b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00106] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0020c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0020d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00107] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0020e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0020f] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00108] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00210] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00211] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00109] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00212] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00213] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0010a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00214] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00215] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0010b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00216] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00217] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0010c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00218] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00219] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0010d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0021a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0021b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0010e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0021c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0021d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0010f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0021e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0021f] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00110] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00220] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00111] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00222] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00223] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00112] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00224] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00225] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00113] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00226] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00227] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00114] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00228] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00229] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00115] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0022a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0022b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00116] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0022c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0022d] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00117] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0022e] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00118] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00230] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00231] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00119] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00232] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00233] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0011a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00234] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00235] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0011b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00236] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00237] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0011c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00238] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0011d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0023a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0023b] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0011e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0023c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0023d] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0011f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0023e] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00120] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00240] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00241] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00121] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00242] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00243] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00122] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00244] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00245] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00123] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00246] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00124] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00248] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00249] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00125] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0024a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0024b] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00126] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0024c] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00127] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0024e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0024f] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00128] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00250] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00129] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00252] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00253] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0012a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00254] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00255] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0012b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00256] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0012c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00258] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00259] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0012d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0025a] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0012e] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0025c] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0025d] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0012f] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0025e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0025f] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00130] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00260] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00131] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00262] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00263] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00132] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00264] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00133] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00266] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00267] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00134] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00268] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00135] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0026a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0026b] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00136] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0026c] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00137] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0026e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0026f] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00138] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00270] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00139] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00272] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00273] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0013a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00274] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0013b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00276] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00277] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0013c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00278] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0013d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0027a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0027b] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0013e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0027c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0013f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0027e] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00140] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00280] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00281] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00141] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00282] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00142] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00284] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00285] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00143] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00286] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00144] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00288] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00145] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0028a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0028b] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00146] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0028c] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00147] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0028e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0028f] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00148] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00290] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00149] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00292] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0014a] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00294] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00295] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0014b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00296] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0014c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00298] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0014d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0029a] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0029b] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0014e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0029c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0014f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0029e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00150] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00151] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00152] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002a4] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00153] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002a6] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002a7] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00154] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00155] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002aa] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00156] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002ac] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002ad] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00157] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00158] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002b0] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00159] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002b2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002b3] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0015a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0015b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0015c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002b8] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0015d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002ba] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002bb] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0015e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0015f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002be] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00160] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002c0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002c1] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00161] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00162] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00163] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002c6] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00164] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002c8] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002c9] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00165] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00166] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00167] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00168] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002d0] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00169] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002d2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002d3] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0016a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0016b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0016c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002d8] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0016d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002da] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002db] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0016e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0016f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00170] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00171] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002e2] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00172] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002e4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002e5] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00173] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00174] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00175] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00176] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00177] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002ee] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00178] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002f0] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002f1] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00179] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0017a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0017b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0017c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002f8] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0017d] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002fa] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h002fb] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0017e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0017f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h002fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00180] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00300] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00181] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00302] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00182] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00304] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00183] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00306] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00184] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00308] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00309] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00185] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0030a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00186] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0030c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00187] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0030e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00188] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00310] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00189] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00312] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0018a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00314] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0018b] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00316] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00317] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0018c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00318] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0018d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0031a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0018e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0031c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0018f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0031e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00190] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00320] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00191] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00322] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00192] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00324] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00193] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00326] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00327] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00194] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00328] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00195] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0032a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00196] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0032c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00197] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0032e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00198] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00330] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00199] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00332] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0019a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00334] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0019b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00336] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h0019c] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00338] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00339] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0019d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0033a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0019e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0033c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0019f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0033e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00340] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00342] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00344] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00346] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00348] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0034a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0034c] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h001a7] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0034e] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h0034f] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00350] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00352] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00354] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00356] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00358] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0035a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0035c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0035e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00360] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00362] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00364] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00366] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h001b4] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00368] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00369] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0036a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0036c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0036e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00370] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00372] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00374] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00376] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00378] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0037a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0037c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0037e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00380] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00382] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00384] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00386] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h001c4] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00388] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00389] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0038a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0038c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0038e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00390] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00392] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00394] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00396] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00398] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0039a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0039c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0039e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003b0] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h001d9] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h003b2] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h003b3] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003f2] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h001fa] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h003f4] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h003f5] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h001ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h003fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00200] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00400] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00201] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00402] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00202] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00404] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00203] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00406] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00204] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00408] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00205] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0040a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00206] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0040c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00207] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0040e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00208] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00410] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00209] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00412] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0020a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00414] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0020b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00416] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0020c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00418] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0020d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0041a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0020e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0041c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0020f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0041e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00210] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00420] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00211] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00422] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00212] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00424] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00213] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00426] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00214] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00428] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00215] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0042a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00216] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0042c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00217] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0042e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00218] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00430] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00219] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00432] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0021a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00434] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0021b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00436] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0021c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00438] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0021d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0043a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0021e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0043c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0021f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0043e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00220] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00440] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00221] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00442] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00222] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00444] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00223] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00446] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00224] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00448] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00225] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0044a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00226] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0044c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00227] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0044e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00228] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00450] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00229] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00452] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0022a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00454] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0022b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00456] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0022c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00458] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0022d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0045a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0022e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0045c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0022f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0045e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00230] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00460] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00231] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00462] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00232] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00464] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00233] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00466] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00234] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00468] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00235] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0046a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00236] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0046c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00237] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0046e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00238] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00470] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00239] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00472] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0023a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00474] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0023b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00476] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0023c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00478] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0023d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0047a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0023e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0047c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0023f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0047e] ;
//end
//always_comb begin
              Ifd35529b44c957737bf422127283c08e['h00240] = 
          (!fgallag_sel['h00004]) ? 
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00480] : //%
                       I6eb3a3e04397efbe48cc2f5809bfcb98['h00481] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00241] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00482] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00242] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00484] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00243] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00486] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00244] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00488] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00245] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0048a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00246] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0048c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00247] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0048e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00248] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00490] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00249] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00492] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0024a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00494] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0024b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00496] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0024c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00498] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0024d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0049a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0024e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0049c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0024f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0049e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00250] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00251] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00252] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00253] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00254] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00255] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00256] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00257] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00258] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00259] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0025a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0025b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0025c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0025d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0025e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0025f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00260] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00261] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00262] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00263] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00264] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00265] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00266] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00267] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00268] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00269] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0026a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0026b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0026c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0026d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0026e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0026f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00270] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00271] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00272] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00273] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00274] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00275] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00276] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00277] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00278] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00279] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0027a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0027b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0027c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0027d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0027e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0027f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h004fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00280] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00500] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00281] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00502] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00282] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00504] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00283] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00506] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00284] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00508] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00285] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0050a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00286] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0050c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00287] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0050e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00288] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00510] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00289] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00512] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0028a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00514] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0028b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00516] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0028c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00518] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0028d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0051a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0028e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0051c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0028f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0051e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00290] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00520] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00291] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00522] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00292] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00524] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00293] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00526] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00294] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00528] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00295] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0052a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00296] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0052c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00297] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0052e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00298] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00530] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00299] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00532] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0029a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00534] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0029b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00536] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0029c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00538] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0029d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0053a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0029e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0053c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0029f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0053e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00540] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00542] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00544] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00546] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00548] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0054a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0054c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0054e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00550] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00552] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00554] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00556] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00558] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0055a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0055c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0055e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00560] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00562] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00564] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00566] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00568] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0056a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0056c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0056e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00570] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00572] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00574] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00576] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00578] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0057a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0057c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0057e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00580] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00582] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00584] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00586] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00588] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0058a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0058c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0058e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00590] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00592] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00594] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00596] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00598] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0059a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0059c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0059e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h002ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h005fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00300] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00600] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00301] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00602] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00302] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00604] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00303] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00606] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00304] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00608] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00305] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0060a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00306] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0060c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00307] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0060e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00308] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00610] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00309] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00612] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0030a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00614] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0030b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00616] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0030c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00618] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0030d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0061a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0030e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0061c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0030f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0061e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00310] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00620] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00311] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00622] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00312] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00624] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00313] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00626] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00314] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00628] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00315] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0062a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00316] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0062c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00317] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0062e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00318] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00630] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00319] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00632] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0031a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00634] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0031b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00636] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0031c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00638] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0031d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0063a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0031e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0063c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0031f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0063e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00320] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00640] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00321] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00642] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00322] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00644] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00323] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00646] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00324] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00648] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00325] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0064a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00326] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0064c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00327] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0064e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00328] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00650] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00329] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00652] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0032a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00654] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0032b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00656] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0032c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00658] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0032d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0065a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0032e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0065c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0032f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0065e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00330] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00660] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00331] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00662] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00332] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00664] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00333] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00666] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00334] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00668] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00335] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0066a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00336] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0066c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00337] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0066e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00338] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00670] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00339] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00672] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0033a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00674] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0033b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00676] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0033c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00678] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0033d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0067a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0033e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0067c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0033f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0067e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00340] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00680] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00341] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00682] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00342] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00684] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00343] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00686] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00344] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00688] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00345] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0068a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00346] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0068c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00347] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0068e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00348] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00690] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00349] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00692] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0034a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00694] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0034b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00696] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0034c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00698] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0034d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0069a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0034e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0069c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0034f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0069e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00350] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00351] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00352] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00353] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00354] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00355] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00356] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00357] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00358] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00359] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0035a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0035b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0035c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0035d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0035e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0035f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00360] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00361] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00362] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00363] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00364] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00365] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00366] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00367] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00368] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00369] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0036a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0036b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0036c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0036d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0036e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0036f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00370] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00371] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00372] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00373] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00374] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00375] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00376] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00377] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00378] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00379] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0037a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0037b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0037c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0037d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0037e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0037f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h006fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00380] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00700] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00381] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00702] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00382] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00704] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00383] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00706] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00384] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00708] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00385] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0070a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00386] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0070c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00387] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0070e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00388] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00710] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00389] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00712] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0038a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00714] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0038b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00716] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0038c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00718] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0038d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0071a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0038e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0071c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0038f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0071e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00390] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00720] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00391] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00722] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00392] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00724] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00393] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00726] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00394] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00728] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00395] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0072a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00396] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0072c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00397] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0072e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00398] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00730] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00399] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00732] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0039a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00734] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0039b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00736] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0039c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00738] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0039d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0073a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0039e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0073c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0039f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0073e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00740] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00742] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00744] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00746] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00748] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0074a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0074c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0074e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00750] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00752] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00754] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00756] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00758] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0075a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0075c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0075e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00760] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00762] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00764] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00766] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00768] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0076a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0076c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0076e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00770] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00772] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00774] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00776] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00778] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0077a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0077c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0077e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00780] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00782] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00784] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00786] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00788] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0078a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0078c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0078e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00790] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00792] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00794] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00796] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00798] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0079a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0079c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0079e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h003ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h007fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00400] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00800] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00401] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00802] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00402] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00804] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00403] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00806] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00404] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00808] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00405] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0080a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00406] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0080c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00407] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0080e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00408] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00810] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00409] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00812] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0040a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00814] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0040b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00816] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0040c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00818] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0040d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0081a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0040e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0081c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0040f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0081e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00410] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00820] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00411] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00822] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00412] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00824] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00413] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00826] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00414] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00828] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00415] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0082a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00416] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0082c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00417] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0082e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00418] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00830] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00419] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00832] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0041a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00834] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0041b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00836] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0041c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00838] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0041d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0083a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0041e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0083c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0041f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0083e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00420] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00840] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00421] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00842] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00422] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00844] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00423] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00846] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00424] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00848] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00425] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0084a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00426] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0084c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00427] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0084e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00428] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00850] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00429] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00852] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0042a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00854] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0042b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00856] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0042c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00858] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0042d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0085a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0042e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0085c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0042f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0085e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00430] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00860] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00431] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00862] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00432] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00864] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00433] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00866] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00434] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00868] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00435] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0086a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00436] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0086c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00437] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0086e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00438] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00870] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00439] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00872] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0043a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00874] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0043b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00876] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0043c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00878] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0043d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0087a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0043e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0087c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0043f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0087e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00440] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00880] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00441] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00882] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00442] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00884] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00443] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00886] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00444] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00888] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00445] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0088a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00446] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0088c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00447] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0088e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00448] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00890] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00449] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00892] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0044a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00894] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0044b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00896] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0044c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00898] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0044d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0089a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0044e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0089c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0044f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0089e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00450] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00451] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00452] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00453] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00454] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00455] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00456] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00457] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00458] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00459] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0045a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0045b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0045c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0045d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0045e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0045f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00460] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00461] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00462] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00463] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00464] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00465] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00466] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00467] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00468] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00469] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0046a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0046b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0046c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0046d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0046e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0046f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00470] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00471] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00472] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00473] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00474] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00475] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00476] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00477] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00478] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00479] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0047a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0047b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0047c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0047d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0047e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0047f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h008fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00480] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00900] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00481] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00902] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00482] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00904] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00483] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00906] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00484] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00908] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00485] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0090a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00486] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0090c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00487] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0090e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00488] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00910] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00489] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00912] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0048a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00914] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0048b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00916] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0048c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00918] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0048d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0091a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0048e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0091c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0048f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0091e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00490] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00920] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00491] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00922] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00492] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00924] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00493] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00926] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00494] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00928] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00495] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0092a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00496] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0092c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00497] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0092e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00498] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00930] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00499] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00932] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0049a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00934] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0049b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00936] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0049c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00938] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0049d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0093a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0049e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0093c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0049f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0093e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00940] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00942] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00944] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00946] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00948] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0094a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0094c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0094e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00950] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00952] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00954] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00956] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00958] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0095a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0095c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0095e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00960] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00962] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00964] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00966] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00968] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0096a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0096c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0096e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00970] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00972] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00974] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00976] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00978] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0097a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0097c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0097e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00980] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00982] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00984] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00986] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00988] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0098a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0098c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0098e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00990] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00992] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00994] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00996] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00998] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0099a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0099c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0099e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h004ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h009fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00500] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00501] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00502] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00503] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00504] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00505] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00506] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00507] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00508] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00509] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0050a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0050b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0050c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0050d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0050e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0050f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00510] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00511] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00512] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00513] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00514] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00515] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00516] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00517] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00518] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00519] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0051a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0051b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0051c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0051d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0051e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0051f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00520] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00521] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00522] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00523] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00524] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00525] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00526] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00527] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00528] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00529] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0052a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0052b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0052c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0052d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0052e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0052f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00530] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00531] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00532] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00533] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00534] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00535] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00536] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00537] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00538] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00539] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0053a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0053b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0053c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0053d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0053e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0053f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00540] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00541] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00542] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00543] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00544] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00545] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00546] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00547] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00548] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00549] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0054a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0054b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0054c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0054d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0054e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0054f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00a9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00550] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00551] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00552] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00553] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00554] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00555] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00556] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00557] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00558] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ab0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00559] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ab2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0055a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ab4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0055b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ab6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0055c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ab8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0055d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0055e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00abc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0055f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00abe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00560] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ac0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00561] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ac2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00562] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ac4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00563] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ac6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00564] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ac8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00565] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00566] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00acc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00567] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ace] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00568] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ad0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00569] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ad2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0056a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ad4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0056b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ad6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0056c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ad8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0056d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ada] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0056e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00adc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0056f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ade] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00570] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ae0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00571] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ae2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00572] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ae4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00573] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ae6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00574] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ae8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00575] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00576] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00577] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00aee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00578] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00af0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00579] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00af2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0057a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00af4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0057b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00af6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0057c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00af8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0057d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00afa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0057e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00afc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0057f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00afe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00580] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00581] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00582] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00583] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00584] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00585] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00586] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00587] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00588] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00589] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0058a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0058b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0058c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0058d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0058e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0058f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00590] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00591] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00592] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00593] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00594] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00595] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00596] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00597] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00598] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00599] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0059a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0059b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0059c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0059d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0059e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0059f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00b9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ba0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ba2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ba4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ba6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ba8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00baa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00be0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00be2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00be4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00be6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00be8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h005ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00bfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00600] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00601] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00602] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00603] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00604] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00605] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00606] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00607] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00608] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00609] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0060a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0060b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0060c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0060d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0060e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0060f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00610] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00611] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00612] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00613] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00614] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00615] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00616] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00617] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00618] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00619] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0061a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0061b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0061c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0061d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0061e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0061f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00620] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00621] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00622] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00623] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00624] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00625] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00626] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00627] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00628] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00629] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0062a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0062b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0062c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0062d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0062e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0062f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00630] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00631] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00632] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00633] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00634] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00635] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00636] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00637] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00638] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00639] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0063a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0063b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0063c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0063d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0063e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0063f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00640] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00641] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00642] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00643] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00644] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00645] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00646] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00647] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00648] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00649] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0064a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0064b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0064c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0064d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0064e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0064f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00c9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00650] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ca0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00651] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ca2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00652] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ca4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00653] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ca6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00654] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ca8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00655] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00caa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00656] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00657] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00658] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00659] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0065a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0065b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0065c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0065d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0065e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0065f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00660] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00661] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00662] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00663] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00664] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00665] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00666] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ccc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00667] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00668] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00669] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0066a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0066b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0066c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0066d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0066e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0066f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00670] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ce0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00671] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ce2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00672] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ce4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00673] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ce6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00674] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ce8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00675] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00676] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00677] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00678] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00679] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0067a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0067b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0067c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0067d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0067e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0067f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00cfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00680] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00681] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00682] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00683] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00684] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00685] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00686] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00687] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00688] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00689] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0068a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0068b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0068c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0068d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0068e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0068f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00690] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00691] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00692] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00693] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00694] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00695] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00696] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00697] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00698] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00699] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0069a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0069b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0069c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0069d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0069e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0069f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00d9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00da0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00da2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00da4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00da6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00da8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00daa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00db0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00db2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00db4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00db6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00db8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ddc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00de0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00de2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00de4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00de6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00de8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00df0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00df2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00df4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00df6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00df8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h006ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00dfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00700] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00701] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00702] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00703] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00704] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00705] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00706] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00707] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00708] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00709] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0070a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0070b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0070c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0070d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0070e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0070f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00710] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00711] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00712] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00713] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00714] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00715] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00716] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00717] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00718] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00719] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0071a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0071b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0071c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0071d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0071e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0071f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00720] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00721] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00722] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00723] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00724] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00725] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00726] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00727] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00728] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00729] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0072a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0072b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0072c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0072d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0072e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0072f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00730] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00731] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00732] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00733] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00734] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00735] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00736] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00737] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00738] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00739] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0073a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0073b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0073c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0073d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0073e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0073f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00740] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00741] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00742] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00743] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00744] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00745] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00746] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00747] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00748] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00749] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0074a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0074b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0074c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0074d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0074e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0074f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00e9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00750] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ea0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00751] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ea2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00752] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ea4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00753] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ea6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00754] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ea8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00755] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00756] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00757] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00758] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00759] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0075a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0075b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0075c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0075d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0075e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ebc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0075f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ebe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00760] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ec0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00761] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ec2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00762] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ec4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00763] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ec6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00764] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ec8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00765] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00766] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ecc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00767] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ece] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00768] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ed0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00769] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ed2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0076a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ed4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0076b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ed6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0076c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ed8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0076d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0076e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00edc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0076f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ede] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00770] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ee0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00771] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ee2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00772] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ee4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00773] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ee6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00774] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ee8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00775] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00776] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00777] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00eee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00778] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ef0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00779] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ef2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0077a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ef4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0077b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ef6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0077c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ef8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0077d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00efa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0077e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00efc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0077f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00efe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00780] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00781] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00782] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00783] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00784] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00785] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00786] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00787] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00788] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00789] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0078a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0078b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0078c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0078d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0078e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0078f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00790] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00791] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00792] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00793] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00794] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00795] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00796] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00797] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00798] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00799] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0079a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0079b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0079c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0079d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0079e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0079f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00f9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00faa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fe0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fe2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fe4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fe6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fe8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00fee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ff0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ff2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ff4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ff6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ff8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ffa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ffc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h007ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h00ffe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00800] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01000] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00801] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01002] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00802] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01004] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00803] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01006] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00804] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01008] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00805] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0100a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00806] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0100c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00807] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0100e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00808] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01010] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00809] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01012] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0080a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01014] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0080b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01016] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0080c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01018] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0080d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0101a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0080e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0101c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0080f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0101e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00810] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01020] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00811] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01022] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00812] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01024] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00813] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01026] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00814] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01028] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00815] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0102a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00816] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0102c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00817] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0102e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00818] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01030] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00819] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01032] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0081a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01034] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0081b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01036] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0081c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01038] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0081d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0103a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0081e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0103c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0081f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0103e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00820] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01040] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00821] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01042] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00822] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01044] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00823] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01046] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00824] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01048] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00825] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0104a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00826] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0104c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00827] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0104e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00828] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01050] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00829] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01052] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0082a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01054] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0082b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01056] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0082c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01058] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0082d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0105a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0082e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0105c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0082f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0105e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00830] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01060] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00831] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01062] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00832] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01064] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00833] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01066] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00834] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01068] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00835] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0106a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00836] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0106c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00837] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0106e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00838] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01070] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00839] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01072] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0083a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01074] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0083b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01076] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0083c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01078] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0083d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0107a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0083e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0107c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0083f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0107e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00840] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01080] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00841] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01082] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00842] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01084] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00843] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01086] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00844] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01088] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00845] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0108a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00846] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0108c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00847] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0108e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00848] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01090] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00849] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01092] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0084a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01094] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0084b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01096] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0084c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01098] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0084d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0109a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0084e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0109c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0084f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0109e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00850] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00851] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00852] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00853] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00854] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00855] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00856] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00857] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00858] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00859] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0085a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0085b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0085c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0085d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0085e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0085f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00860] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00861] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00862] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00863] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00864] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00865] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00866] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00867] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00868] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00869] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0086a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0086b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0086c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0086d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0086e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0086f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00870] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00871] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00872] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00873] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00874] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00875] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00876] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00877] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00878] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00879] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0087a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0087b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0087c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0087d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0087e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0087f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h010fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00880] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01100] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00881] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01102] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00882] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01104] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00883] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01106] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00884] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01108] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00885] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0110a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00886] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0110c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00887] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0110e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00888] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01110] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00889] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01112] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0088a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01114] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0088b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01116] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0088c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01118] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0088d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0111a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0088e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0111c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0088f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0111e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00890] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01120] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00891] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01122] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00892] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01124] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00893] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01126] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00894] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01128] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00895] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0112a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00896] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0112c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00897] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0112e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00898] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01130] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00899] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01132] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0089a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01134] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0089b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01136] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0089c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01138] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0089d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0113a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0089e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0113c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0089f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0113e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01140] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01142] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01144] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01146] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01148] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0114a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0114c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0114e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01150] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01152] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01154] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01156] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01158] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0115a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0115c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0115e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01160] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01162] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01164] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01166] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01168] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0116a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0116c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0116e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01170] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01172] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01174] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01176] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01178] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0117a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0117c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0117e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01180] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01182] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01184] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01186] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01188] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0118a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0118c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0118e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01190] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01192] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01194] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01196] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01198] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0119a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0119c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0119e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h008ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h011fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00900] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01200] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00901] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01202] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00902] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01204] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00903] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01206] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00904] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01208] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00905] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0120a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00906] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0120c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00907] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0120e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00908] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01210] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00909] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01212] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0090a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01214] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0090b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01216] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0090c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01218] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0090d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0121a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0090e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0121c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0090f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0121e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00910] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01220] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00911] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01222] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00912] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01224] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00913] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01226] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00914] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01228] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00915] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0122a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00916] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0122c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00917] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0122e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00918] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01230] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00919] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01232] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0091a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01234] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0091b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01236] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0091c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01238] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0091d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0123a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0091e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0123c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0091f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0123e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00920] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01240] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00921] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01242] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00922] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01244] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00923] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01246] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00924] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01248] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00925] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0124a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00926] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0124c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00927] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0124e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00928] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01250] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00929] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01252] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0092a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01254] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0092b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01256] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0092c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01258] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0092d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0125a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0092e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0125c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0092f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0125e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00930] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01260] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00931] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01262] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00932] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01264] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00933] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01266] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00934] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01268] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00935] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0126a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00936] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0126c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00937] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0126e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00938] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01270] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00939] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01272] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0093a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01274] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0093b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01276] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0093c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01278] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0093d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0127a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0093e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0127c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0093f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0127e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00940] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01280] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00941] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01282] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00942] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01284] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00943] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01286] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00944] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01288] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00945] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0128a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00946] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0128c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00947] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0128e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00948] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01290] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00949] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01292] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0094a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01294] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0094b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01296] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0094c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01298] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0094d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0129a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0094e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0129c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0094f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0129e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00950] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00951] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00952] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00953] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00954] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00955] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00956] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00957] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00958] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00959] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0095a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0095b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0095c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0095d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0095e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0095f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00960] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00961] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00962] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00963] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00964] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00965] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00966] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00967] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00968] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00969] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0096a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0096b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0096c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0096d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0096e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0096f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00970] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00971] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00972] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00973] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00974] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00975] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00976] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00977] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00978] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00979] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0097a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0097b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0097c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0097d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0097e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0097f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h012fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00980] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01300] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00981] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01302] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00982] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01304] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00983] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01306] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00984] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01308] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00985] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0130a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00986] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0130c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00987] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0130e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00988] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01310] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00989] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01312] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0098a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01314] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0098b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01316] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0098c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01318] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0098d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0131a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0098e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0131c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0098f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0131e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00990] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01320] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00991] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01322] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00992] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01324] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00993] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01326] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00994] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01328] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00995] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0132a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00996] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0132c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00997] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0132e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00998] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01330] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00999] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01332] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0099a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01334] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0099b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01336] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0099c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01338] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0099d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0133a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0099e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0133c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0099f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0133e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01340] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01342] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01344] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01346] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01348] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0134a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0134c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0134e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01350] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01352] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01354] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01356] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01358] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0135a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0135c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0135e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01360] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01362] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01364] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01366] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01368] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0136a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0136c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0136e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01370] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01372] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01374] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01376] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01378] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0137a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0137c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0137e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01380] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01382] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01384] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01386] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01388] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0138a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0138c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0138e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01390] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01392] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01394] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01396] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01398] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0139a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0139c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0139e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h009ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h013fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01400] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01402] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01404] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01406] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01408] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0140a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0140c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0140e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01410] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01412] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01414] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01416] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01418] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0141a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0141c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0141e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01420] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01422] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01424] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01426] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01428] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0142a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0142c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0142e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01430] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01432] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01434] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01436] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01438] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0143a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0143c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0143e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01440] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01442] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01444] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01446] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01448] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0144a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0144c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0144e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01450] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01452] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01454] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01456] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01458] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0145a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0145c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0145e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01460] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01462] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01464] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01466] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01468] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0146a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0146c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0146e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01470] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01472] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01474] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01476] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01478] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0147a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0147c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0147e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01480] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01482] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01484] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01486] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01488] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0148a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0148c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0148e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01490] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01492] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01494] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01496] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01498] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0149a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0149c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0149e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h014fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01500] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01502] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01504] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01506] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01508] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0150a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0150c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0150e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01510] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01512] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01514] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01516] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01518] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0151a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0151c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0151e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01520] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01522] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01524] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01526] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01528] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0152a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0152c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0152e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01530] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01532] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01534] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01536] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01538] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0153a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0153c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00a9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0153e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aa0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01540] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aa1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01542] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aa2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01544] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aa3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01546] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aa4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01548] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aa5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0154a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aa6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0154c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aa7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0154e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aa8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01550] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aa9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01552] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aaa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01554] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01556] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01558] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0155a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0155c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aaf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0155e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ab0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01560] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ab1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01562] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ab2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01564] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ab3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01566] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ab4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01568] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ab5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0156a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ab6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0156c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ab7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0156e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ab8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01570] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ab9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01572] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01574] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00abb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01576] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00abc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01578] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00abd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0157a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00abe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0157c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00abf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0157e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ac0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01580] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ac1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01582] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ac2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01584] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ac3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01586] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ac4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01588] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ac5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0158a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ac6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0158c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ac7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0158e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ac8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01590] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ac9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01592] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01594] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00acb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01596] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00acc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01598] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00acd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0159a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ace] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0159c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00acf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0159e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ad0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ad1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ad2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ad3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ad4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ad5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ad6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ad7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ad8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ad9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ada] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00adb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00adc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00add] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ade] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00adf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ae0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ae1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ae2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ae3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ae4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ae5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ae6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ae7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ae8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ae9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aeb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00af0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00af1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00af2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00af3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00af4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00af5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00af6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00af7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00af8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00af9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00afa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00afb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00afc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00afd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00afe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00aff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h015fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01600] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01602] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01604] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01606] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01608] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0160a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0160c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0160e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01610] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01612] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01614] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01616] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01618] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0161a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0161c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0161e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01620] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01622] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01624] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01626] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01628] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0162a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0162c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0162e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01630] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01632] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01634] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01636] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01638] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0163a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0163c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0163e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01640] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01642] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01644] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01646] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01648] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0164a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0164c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0164e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01650] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01652] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01654] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01656] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01658] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0165a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0165c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0165e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01660] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01662] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01664] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01666] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01668] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0166a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0166c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0166e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01670] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01672] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01674] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01676] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01678] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0167a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0167c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0167e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01680] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01682] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01684] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01686] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01688] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0168a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0168c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0168e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01690] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01692] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01694] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01696] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01698] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0169a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0169c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0169e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h016fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01700] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01702] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01704] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01706] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01708] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0170a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0170c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0170e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01710] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01712] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01714] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01716] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01718] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0171a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0171c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0171e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01720] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01722] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01724] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01726] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01728] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0172a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0172c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0172e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01730] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01732] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01734] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01736] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01738] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0173a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0173c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00b9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0173e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ba0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01740] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ba1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01742] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ba2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01744] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ba3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01746] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ba4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01748] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ba5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0174a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ba6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0174c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ba7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0174e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ba8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01750] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ba9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01752] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00baa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01754] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01756] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01758] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0175a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0175c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00baf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0175e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01760] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01762] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01764] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01766] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01768] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0176a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0176c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0176e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01770] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01772] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01774] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01776] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01778] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0177a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0177c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0177e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01780] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01782] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01784] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01786] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01788] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0178a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0178c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0178e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01790] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01792] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01794] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01796] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01798] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0179a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0179c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0179e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00be0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00be1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00be2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00be3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00be4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00be5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00be6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00be7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00be8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00be9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00beb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bf0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bf1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bf2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bf3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bf4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bf5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bf6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bf7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bf8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bf9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00bff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h017fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01800] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01802] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01804] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01806] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01808] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0180a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0180c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0180e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01810] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01812] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01814] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01816] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01818] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0181a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0181c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0181e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01820] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01822] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01824] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01826] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01828] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0182a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0182c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0182e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01830] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01832] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01834] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01836] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01838] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0183a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0183c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0183e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01840] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01842] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01844] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01846] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01848] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0184a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0184c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0184e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01850] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01852] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01854] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01856] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01858] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0185a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0185c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0185e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01860] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01862] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01864] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01866] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01868] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0186a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0186c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0186e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01870] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01872] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01874] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01876] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01878] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0187a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0187c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0187e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01880] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01882] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01884] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01886] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01888] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0188a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0188c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0188e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01890] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01892] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01894] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01896] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01898] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0189a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0189c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0189e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h018fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01900] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01902] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01904] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01906] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01908] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0190a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0190c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0190e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01910] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01912] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01914] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01916] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01918] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0191a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0191c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0191e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01920] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01922] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01924] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01926] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01928] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0192a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0192c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0192e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01930] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01932] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01934] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01936] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01938] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0193a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0193c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00c9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0193e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ca0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01940] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ca1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01942] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ca2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01944] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ca3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01946] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ca4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01948] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ca5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0194a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ca6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0194c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ca7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0194e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ca8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01950] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ca9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01952] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00caa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01954] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01956] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01958] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0195a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0195c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00caf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0195e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01960] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01962] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01964] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01966] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01968] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0196a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0196c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0196e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01970] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01972] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01974] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01976] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01978] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0197a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0197c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0197e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01980] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01982] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01984] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01986] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01988] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0198a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0198c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0198e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01990] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01992] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01994] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ccb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01996] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ccc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01998] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ccd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0199a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0199c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ccf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0199e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ce0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ce1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ce2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ce3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ce4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ce5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ce6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ce7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ce8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ce9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ceb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ced] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cf0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cf1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cf2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cf3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cf4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cf5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cf6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cf7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cf8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cf9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00cff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h019fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01a9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ab0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ab2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ab4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ab6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ab8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01abc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01abe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ac0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ac2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ac4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ac6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ac8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01acc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ace] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ad0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ad2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ad4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ad6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ad8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ada] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01adc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ade] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ae0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ae2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ae4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ae6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ae8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01aee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01af0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01af2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01af4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01af6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01af8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01afa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01afc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01afe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00d9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00da0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00da1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00da2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00da3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00da4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00da5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00da6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00da7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00da8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00da9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00daa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00daf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00db0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00db1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00db2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00db3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00db4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00db5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00db6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00db7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00db8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00db9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01b9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ba0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ba2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ba4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ba6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ba8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01baa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ddb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ddc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ddd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ddf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00de0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00de1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00de2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00de3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00de4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00de5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00de6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00de7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00de8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00de9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00deb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ded] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00def] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00df0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01be0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00df1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01be2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00df2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01be4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00df3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01be6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00df4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01be8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00df5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00df6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00df7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00df8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00df9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00dff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01bfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01c9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ca0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ca2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ca4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ca6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ca8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01caa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ccc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ce0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ce2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ce4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ce6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ce8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01cfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00e9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ea0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ea1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ea2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ea3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ea4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ea5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ea6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ea7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ea8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ea9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eaa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ead] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eaf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ebb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ebc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ebd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ebe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ebf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ec0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ec1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ec2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ec3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ec4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ec5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ec6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ec7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ec8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ec9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ecb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ecc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ecd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ece] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ecf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01d9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ed0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01da0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ed1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01da2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ed2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01da4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ed3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01da6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ed4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01da8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ed5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01daa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ed6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ed7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ed8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01db0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ed9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01db2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01db4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00edb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01db6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00edc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01db8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00edd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ede] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00edf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ee0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ee1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ee2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ee3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ee4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ee5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ee6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ee7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ee8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ee9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eeb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ddc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ef0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01de0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ef1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01de2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ef2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01de4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ef3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01de6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ef4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01de8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ef5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ef6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ef7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ef8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01df0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ef9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01df2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00efa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01df4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00efb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01df6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00efc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01df8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00efd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00efe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00eff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01dfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01e9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ea0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ea2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ea4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ea6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ea8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ebc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ebe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ec0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ec2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ec4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ec6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ec8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ecc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ece] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ed0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ed2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ed4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ed6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ed8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01edc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ede] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ee0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ee2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ee4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ee6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ee8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01eee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ef0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ef2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ef4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ef6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ef8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01efa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01efc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01efe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00f9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fa0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fa1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fa2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fa3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fa4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fa5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fa6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fa7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fa8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fa9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00faa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00faf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01f9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01faa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fe0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fe1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fe2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fe3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fe4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fe5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fe6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fe7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fe8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fe9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00feb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ff0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fe0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ff1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fe2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ff2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fe4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ff3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fe6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ff4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fe8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ff5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ff6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ff7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01fee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ff8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ff0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ff9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ff2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ffa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ff4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ffb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ff6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ffc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ff8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ffd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ffa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00ffe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ffc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h00fff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h01ffe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01000] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02000] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01001] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02002] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01002] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02004] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01003] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02006] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01004] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02008] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01005] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0200a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01006] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0200c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01007] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0200e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01008] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02010] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01009] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02012] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0100a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02014] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0100b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02016] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0100c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02018] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0100d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0201a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0100e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0201c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0100f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0201e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01010] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02020] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01011] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02022] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01012] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02024] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01013] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02026] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01014] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02028] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01015] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0202a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01016] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0202c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01017] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0202e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01018] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02030] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01019] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02032] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0101a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02034] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0101b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02036] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0101c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02038] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0101d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0203a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0101e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0203c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0101f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0203e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01020] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02040] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01021] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02042] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01022] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02044] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01023] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02046] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01024] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02048] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01025] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0204a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01026] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0204c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01027] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0204e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01028] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02050] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01029] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02052] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0102a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02054] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0102b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02056] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0102c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02058] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0102d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0205a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0102e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0205c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0102f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0205e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01030] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02060] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01031] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02062] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01032] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02064] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01033] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02066] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01034] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02068] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01035] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0206a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01036] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0206c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01037] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0206e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01038] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02070] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01039] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02072] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0103a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02074] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0103b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02076] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0103c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02078] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0103d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0207a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0103e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0207c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0103f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0207e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01040] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02080] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01041] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02082] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01042] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02084] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01043] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02086] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01044] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02088] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01045] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0208a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01046] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0208c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01047] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0208e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01048] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02090] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01049] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02092] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0104a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02094] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0104b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02096] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0104c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02098] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0104d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0209a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0104e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0209c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0104f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0209e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01050] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01051] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01052] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01053] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01054] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01055] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01056] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01057] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01058] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01059] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0105a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0105b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0105c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0105d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0105e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0105f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01060] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01061] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01062] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01063] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01064] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01065] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01066] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01067] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01068] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01069] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0106a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0106b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0106c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0106d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0106e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0106f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01070] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01071] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01072] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01073] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01074] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01075] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01076] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01077] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01078] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01079] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0107a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0107b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0107c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0107d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0107e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0107f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h020fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01080] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02100] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01081] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02102] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01082] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02104] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01083] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02106] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01084] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02108] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01085] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0210a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01086] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0210c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01087] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0210e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01088] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02110] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01089] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02112] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0108a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02114] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0108b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02116] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0108c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02118] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0108d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0211a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0108e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0211c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0108f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0211e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01090] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02120] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01091] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02122] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01092] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02124] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01093] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02126] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01094] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02128] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01095] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0212a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01096] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0212c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01097] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0212e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01098] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02130] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01099] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02132] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0109a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02134] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0109b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02136] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0109c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02138] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0109d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0213a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0109e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0213c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0109f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0213e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02140] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02142] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02144] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02146] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02148] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0214a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0214c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0214e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02150] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02152] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02154] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02156] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02158] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0215a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0215c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0215e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02160] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02162] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02164] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02166] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02168] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0216a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0216c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0216e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02170] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02172] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02174] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02176] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02178] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0217a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0217c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0217e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02180] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02182] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02184] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02186] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02188] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0218a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0218c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0218e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02190] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02192] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02194] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02196] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02198] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0219a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0219c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0219e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h010ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h021fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01100] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02200] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01101] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02202] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01102] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02204] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01103] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02206] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01104] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02208] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01105] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0220a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01106] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0220c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01107] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0220e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01108] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02210] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01109] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02212] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0110a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02214] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0110b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02216] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0110c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02218] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0110d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0221a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0110e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0221c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0110f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0221e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01110] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02220] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01111] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02222] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01112] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02224] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01113] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02226] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01114] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02228] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01115] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0222a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01116] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0222c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01117] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0222e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01118] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02230] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01119] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02232] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0111a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02234] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0111b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02236] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0111c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02238] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0111d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0223a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0111e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0223c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0111f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0223e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01120] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02240] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01121] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02242] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01122] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02244] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01123] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02246] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01124] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02248] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01125] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0224a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01126] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0224c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01127] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0224e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01128] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02250] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01129] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02252] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0112a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02254] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0112b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02256] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0112c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02258] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0112d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0225a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0112e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0225c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0112f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0225e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01130] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02260] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01131] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02262] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01132] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02264] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01133] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02266] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01134] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02268] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01135] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0226a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01136] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0226c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01137] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0226e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01138] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02270] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01139] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02272] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0113a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02274] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0113b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02276] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0113c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02278] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0113d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0227a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0113e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0227c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0113f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0227e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01140] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02280] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01141] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02282] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01142] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02284] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01143] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02286] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01144] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02288] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01145] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0228a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01146] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0228c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01147] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0228e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01148] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02290] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01149] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02292] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0114a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02294] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0114b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02296] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0114c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02298] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0114d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0229a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0114e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0229c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0114f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0229e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01150] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01151] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01152] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01153] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01154] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01155] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01156] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01157] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01158] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01159] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0115a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0115b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0115c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0115d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0115e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0115f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01160] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01161] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01162] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01163] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01164] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01165] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01166] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01167] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01168] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01169] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0116a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0116b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0116c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0116d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0116e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0116f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01170] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01171] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01172] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01173] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01174] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01175] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01176] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01177] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01178] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01179] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0117a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0117b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0117c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0117d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0117e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0117f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h022fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01180] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02300] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01181] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02302] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01182] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02304] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01183] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02306] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01184] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02308] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01185] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0230a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01186] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0230c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01187] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0230e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01188] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02310] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01189] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02312] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0118a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02314] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0118b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02316] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0118c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02318] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0118d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0231a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0118e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0231c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0118f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0231e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01190] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02320] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01191] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02322] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01192] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02324] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01193] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02326] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01194] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02328] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01195] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0232a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01196] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0232c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01197] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0232e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01198] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02330] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01199] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02332] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0119a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02334] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0119b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02336] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0119c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02338] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0119d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0233a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0119e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0233c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0119f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0233e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02340] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02342] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02344] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02346] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02348] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0234a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0234c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0234e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02350] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02352] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02354] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02356] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02358] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0235a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0235c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0235e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02360] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02362] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02364] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02366] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02368] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0236a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0236c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0236e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02370] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02372] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02374] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02376] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02378] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0237a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0237c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0237e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02380] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02382] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02384] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02386] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02388] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0238a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0238c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0238e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02390] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02392] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02394] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02396] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02398] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0239a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0239c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0239e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h011ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h023fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01200] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02400] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01201] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02402] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01202] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02404] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01203] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02406] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01204] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02408] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01205] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0240a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01206] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0240c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01207] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0240e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01208] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02410] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01209] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02412] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0120a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02414] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0120b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02416] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0120c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02418] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0120d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0241a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0120e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0241c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0120f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0241e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01210] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02420] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01211] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02422] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01212] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02424] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01213] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02426] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01214] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02428] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01215] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0242a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01216] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0242c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01217] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0242e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01218] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02430] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01219] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02432] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0121a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02434] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0121b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02436] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0121c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02438] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0121d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0243a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0121e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0243c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0121f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0243e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01220] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02440] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01221] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02442] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01222] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02444] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01223] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02446] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01224] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02448] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01225] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0244a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01226] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0244c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01227] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0244e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01228] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02450] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01229] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02452] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0122a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02454] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0122b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02456] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0122c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02458] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0122d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0245a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0122e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0245c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0122f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0245e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01230] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02460] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01231] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02462] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01232] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02464] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01233] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02466] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01234] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02468] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01235] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0246a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01236] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0246c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01237] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0246e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01238] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02470] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01239] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02472] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0123a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02474] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0123b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02476] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0123c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02478] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0123d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0247a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0123e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0247c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0123f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0247e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01240] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02480] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01241] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02482] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01242] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02484] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01243] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02486] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01244] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02488] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01245] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0248a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01246] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0248c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01247] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0248e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01248] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02490] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01249] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02492] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0124a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02494] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0124b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02496] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0124c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02498] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0124d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0249a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0124e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0249c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0124f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0249e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01250] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01251] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01252] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01253] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01254] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01255] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01256] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01257] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01258] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01259] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0125a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0125b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0125c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0125d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0125e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0125f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01260] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01261] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01262] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01263] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01264] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01265] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01266] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01267] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01268] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01269] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0126a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0126b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0126c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0126d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0126e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0126f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01270] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01271] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01272] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01273] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01274] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01275] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01276] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01277] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01278] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01279] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0127a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0127b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0127c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0127d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0127e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0127f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h024fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01280] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02500] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01281] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02502] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01282] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02504] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01283] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02506] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01284] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02508] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01285] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0250a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01286] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0250c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01287] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0250e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01288] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02510] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01289] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02512] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0128a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02514] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0128b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02516] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0128c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02518] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0128d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0251a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0128e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0251c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0128f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0251e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01290] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02520] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01291] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02522] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01292] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02524] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01293] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02526] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01294] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02528] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01295] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0252a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01296] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0252c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01297] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0252e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01298] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02530] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01299] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02532] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0129a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02534] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0129b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02536] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0129c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02538] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0129d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0253a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0129e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0253c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0129f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0253e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02540] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02542] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02544] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02546] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02548] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0254a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0254c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0254e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02550] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02552] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02554] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02556] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02558] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0255a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0255c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0255e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02560] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02562] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02564] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02566] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02568] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0256a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0256c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0256e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02570] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02572] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02574] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02576] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02578] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0257a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0257c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0257e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02580] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02582] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02584] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02586] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02588] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0258a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0258c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0258e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02590] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02592] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02594] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02596] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02598] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0259a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0259c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0259e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h012ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h025fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01300] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02600] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01301] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02602] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01302] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02604] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01303] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02606] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01304] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02608] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01305] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0260a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01306] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0260c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01307] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0260e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01308] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02610] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01309] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02612] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0130a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02614] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0130b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02616] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0130c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02618] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0130d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0261a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0130e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0261c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0130f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0261e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01310] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02620] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01311] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02622] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01312] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02624] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01313] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02626] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01314] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02628] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01315] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0262a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01316] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0262c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01317] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0262e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01318] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02630] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01319] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02632] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0131a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02634] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0131b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02636] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0131c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02638] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0131d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0263a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0131e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0263c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0131f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0263e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01320] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02640] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01321] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02642] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01322] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02644] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01323] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02646] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01324] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02648] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01325] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0264a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01326] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0264c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01327] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0264e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01328] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02650] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01329] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02652] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0132a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02654] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0132b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02656] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0132c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02658] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0132d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0265a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0132e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0265c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0132f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0265e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01330] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02660] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01331] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02662] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01332] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02664] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01333] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02666] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01334] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02668] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01335] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0266a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01336] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0266c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01337] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0266e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01338] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02670] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01339] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02672] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0133a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02674] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0133b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02676] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0133c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02678] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0133d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0267a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0133e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0267c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0133f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0267e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01340] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02680] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01341] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02682] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01342] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02684] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01343] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02686] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01344] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02688] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01345] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0268a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01346] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0268c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01347] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0268e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01348] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02690] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01349] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02692] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0134a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02694] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0134b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02696] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0134c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02698] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0134d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0269a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0134e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0269c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0134f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0269e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01350] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01351] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01352] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01353] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01354] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01355] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01356] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01357] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01358] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01359] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0135a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0135b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0135c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0135d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0135e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0135f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01360] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01361] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01362] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01363] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01364] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01365] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01366] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01367] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01368] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01369] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0136a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0136b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0136c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0136d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0136e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0136f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01370] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01371] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01372] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01373] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01374] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01375] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01376] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01377] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01378] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01379] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0137a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0137b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0137c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0137d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0137e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0137f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h026fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01380] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02700] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01381] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02702] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01382] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02704] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01383] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02706] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01384] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02708] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01385] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0270a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01386] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0270c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01387] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0270e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01388] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02710] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01389] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02712] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0138a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02714] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0138b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02716] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0138c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02718] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0138d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0271a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0138e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0271c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0138f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0271e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01390] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02720] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01391] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02722] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01392] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02724] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01393] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02726] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01394] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02728] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01395] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0272a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01396] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0272c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01397] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0272e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01398] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02730] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01399] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02732] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0139a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02734] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0139b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02736] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0139c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02738] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0139d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0273a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0139e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0273c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0139f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0273e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02740] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02742] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02744] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02746] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02748] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0274a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0274c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0274e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02750] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02752] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02754] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02756] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02758] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0275a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0275c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0275e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02760] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02762] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02764] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02766] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02768] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0276a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0276c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0276e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02770] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02772] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02774] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02776] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02778] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0277a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0277c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0277e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02780] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02782] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02784] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02786] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02788] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0278a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0278c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0278e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02790] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02792] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02794] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02796] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02798] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0279a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0279c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0279e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h013ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h027fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01400] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02800] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01401] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02802] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01402] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02804] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01403] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02806] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01404] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02808] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01405] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0280a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01406] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0280c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01407] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0280e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01408] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02810] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01409] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02812] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0140a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02814] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0140b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02816] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0140c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02818] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0140d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0281a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0140e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0281c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0140f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0281e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01410] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02820] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01411] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02822] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01412] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02824] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01413] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02826] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01414] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02828] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01415] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0282a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01416] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0282c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01417] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0282e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01418] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02830] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01419] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02832] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0141a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02834] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0141b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02836] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0141c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02838] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0141d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0283a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0141e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0283c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0141f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0283e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01420] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02840] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01421] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02842] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01422] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02844] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01423] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02846] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01424] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02848] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01425] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0284a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01426] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0284c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01427] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0284e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01428] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02850] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01429] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02852] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0142a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02854] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0142b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02856] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0142c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02858] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0142d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0285a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0142e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0285c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0142f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0285e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01430] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02860] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01431] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02862] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01432] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02864] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01433] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02866] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01434] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02868] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01435] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0286a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01436] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0286c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01437] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0286e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01438] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02870] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01439] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02872] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0143a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02874] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0143b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02876] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0143c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02878] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0143d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0287a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0143e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0287c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0143f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0287e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01440] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02880] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01441] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02882] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01442] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02884] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01443] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02886] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01444] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02888] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01445] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0288a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01446] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0288c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01447] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0288e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01448] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02890] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01449] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02892] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0144a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02894] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0144b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02896] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0144c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02898] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0144d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0289a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0144e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0289c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0144f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0289e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01450] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01451] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01452] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01453] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01454] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01455] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01456] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01457] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01458] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01459] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0145a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0145b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0145c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0145d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0145e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0145f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01460] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01461] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01462] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01463] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01464] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01465] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01466] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01467] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01468] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01469] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0146a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0146b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0146c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0146d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0146e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0146f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01470] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01471] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01472] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01473] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01474] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01475] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01476] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01477] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01478] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01479] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0147a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0147b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0147c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0147d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0147e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0147f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h028fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01480] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02900] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01481] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02902] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01482] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02904] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01483] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02906] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01484] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02908] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01485] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0290a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01486] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0290c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01487] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0290e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01488] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02910] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01489] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02912] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0148a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02914] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0148b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02916] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0148c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02918] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0148d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0291a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0148e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0291c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0148f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0291e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01490] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02920] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01491] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02922] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01492] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02924] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01493] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02926] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01494] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02928] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01495] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0292a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01496] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0292c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01497] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0292e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01498] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02930] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01499] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02932] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0149a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02934] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0149b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02936] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0149c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02938] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0149d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0293a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0149e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0293c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0149f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0293e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02940] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02942] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02944] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02946] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02948] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0294a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0294c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0294e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02950] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02952] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02954] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02956] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02958] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0295a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0295c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0295e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02960] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02962] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02964] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02966] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02968] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0296a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0296c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0296e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02970] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02972] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02974] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02976] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02978] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0297a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0297c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0297e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02980] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02982] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02984] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02986] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02988] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0298a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0298c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0298e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02990] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02992] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02994] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02996] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02998] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0299a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0299c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0299e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h014ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h029fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01500] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01501] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01502] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01503] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01504] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01505] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01506] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01507] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01508] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01509] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0150a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0150b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0150c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0150d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0150e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0150f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01510] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01511] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01512] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01513] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01514] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01515] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01516] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01517] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01518] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01519] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0151a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0151b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0151c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0151d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0151e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0151f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01520] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01521] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01522] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01523] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01524] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01525] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01526] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01527] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01528] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01529] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0152a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0152b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0152c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0152d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0152e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0152f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01530] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01531] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01532] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01533] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01534] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01535] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01536] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01537] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01538] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01539] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0153a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0153b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0153c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0153d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0153e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0153f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01540] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01541] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01542] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01543] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01544] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01545] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01546] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01547] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01548] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01549] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0154a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0154b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0154c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0154d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0154e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0154f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02a9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01550] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01551] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01552] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01553] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01554] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01555] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01556] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01557] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01558] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ab0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01559] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ab2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0155a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ab4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0155b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ab6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0155c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ab8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0155d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0155e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02abc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0155f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02abe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01560] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ac0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01561] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ac2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01562] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ac4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01563] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ac6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01564] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ac8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01565] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01566] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02acc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01567] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ace] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01568] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ad0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01569] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ad2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0156a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ad4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0156b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ad6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0156c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ad8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0156d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ada] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0156e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02adc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0156f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ade] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01570] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ae0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01571] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ae2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01572] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ae4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01573] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ae6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01574] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ae8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01575] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01576] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01577] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02aee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01578] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02af0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01579] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02af2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0157a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02af4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0157b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02af6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0157c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02af8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0157d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02afa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0157e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02afc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0157f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02afe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01580] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01581] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01582] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01583] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01584] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01585] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01586] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01587] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01588] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01589] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0158a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0158b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0158c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0158d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0158e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0158f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01590] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01591] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01592] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01593] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01594] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01595] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01596] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01597] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01598] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01599] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0159a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0159b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0159c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0159d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0159e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0159f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02b9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ba0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ba2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ba4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ba6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ba8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02baa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02be0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02be2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02be4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02be6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02be8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h015ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02bfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01600] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01601] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01602] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01603] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01604] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01605] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01606] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01607] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01608] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01609] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0160a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0160b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0160c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0160d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0160e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0160f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01610] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01611] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01612] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01613] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01614] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01615] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01616] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01617] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01618] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01619] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0161a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0161b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0161c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0161d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0161e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0161f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01620] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01621] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01622] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01623] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01624] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01625] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01626] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01627] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01628] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01629] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0162a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0162b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0162c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0162d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0162e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0162f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01630] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01631] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01632] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01633] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01634] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01635] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01636] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01637] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01638] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01639] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0163a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0163b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0163c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0163d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0163e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0163f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01640] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01641] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01642] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01643] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01644] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01645] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01646] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01647] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01648] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01649] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0164a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0164b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0164c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0164d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0164e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0164f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02c9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01650] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ca0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01651] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ca2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01652] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ca4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01653] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ca6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01654] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ca8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01655] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02caa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01656] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01657] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01658] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01659] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0165a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0165b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0165c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0165d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0165e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0165f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01660] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01661] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01662] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01663] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01664] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01665] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01666] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ccc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01667] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01668] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01669] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0166a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0166b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0166c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0166d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0166e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0166f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01670] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ce0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01671] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ce2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01672] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ce4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01673] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ce6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01674] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ce8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01675] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01676] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01677] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01678] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01679] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0167a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0167b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0167c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0167d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0167e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0167f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02cfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01680] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01681] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01682] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01683] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01684] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01685] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01686] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01687] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01688] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01689] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0168a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0168b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0168c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0168d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0168e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0168f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01690] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01691] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01692] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01693] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01694] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01695] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01696] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01697] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01698] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01699] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0169a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0169b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0169c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0169d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0169e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0169f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02d9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02da0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02da2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02da4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02da6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02da8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02daa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02db0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02db2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02db4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02db6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02db8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ddc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02de0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02de2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02de4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02de6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02de8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02df0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02df2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02df4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02df6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02df8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h016ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02dfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01700] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01701] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01702] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01703] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01704] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01705] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01706] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01707] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01708] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01709] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0170a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0170b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0170c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0170d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0170e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0170f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01710] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01711] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01712] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01713] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01714] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01715] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01716] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01717] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01718] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01719] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0171a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0171b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0171c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0171d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0171e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0171f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01720] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01721] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01722] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01723] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01724] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01725] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01726] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01727] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01728] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01729] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0172a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0172b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0172c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0172d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0172e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0172f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01730] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01731] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01732] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01733] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01734] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01735] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01736] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01737] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01738] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01739] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0173a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0173b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0173c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0173d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0173e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0173f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01740] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01741] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01742] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01743] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01744] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01745] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01746] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01747] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01748] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01749] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0174a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0174b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0174c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0174d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0174e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0174f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02e9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01750] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ea0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01751] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ea2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01752] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ea4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01753] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ea6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01754] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ea8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01755] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01756] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01757] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01758] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01759] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0175a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0175b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0175c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0175d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0175e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ebc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0175f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ebe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01760] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ec0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01761] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ec2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01762] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ec4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01763] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ec6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01764] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ec8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01765] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01766] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ecc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01767] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ece] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01768] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ed0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01769] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ed2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0176a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ed4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0176b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ed6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0176c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ed8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0176d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0176e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02edc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0176f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ede] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01770] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ee0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01771] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ee2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01772] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ee4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01773] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ee6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01774] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ee8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01775] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01776] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01777] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02eee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01778] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ef0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01779] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ef2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0177a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ef4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0177b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ef6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0177c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ef8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0177d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02efa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0177e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02efc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0177f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02efe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01780] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01781] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01782] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01783] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01784] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01785] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01786] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01787] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01788] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01789] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0178a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0178b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0178c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0178d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0178e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0178f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01790] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01791] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01792] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01793] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01794] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01795] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01796] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01797] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01798] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01799] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0179a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0179b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0179c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0179d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0179e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0179f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02f9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02faa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fe0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fe2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fe4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fe6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fe8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02fee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ff0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ff2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ff4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ff6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ff8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ffa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ffc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h017ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h02ffe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01800] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03000] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01801] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03002] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01802] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03004] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01803] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03006] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01804] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03008] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01805] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0300a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01806] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0300c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01807] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0300e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01808] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03010] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01809] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03012] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0180a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03014] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0180b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03016] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0180c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03018] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0180d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0301a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0180e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0301c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0180f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0301e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01810] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03020] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01811] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03022] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01812] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03024] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01813] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03026] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01814] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03028] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01815] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0302a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01816] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0302c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01817] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0302e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01818] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03030] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01819] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03032] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0181a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03034] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0181b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03036] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0181c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03038] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0181d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0303a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0181e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0303c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0181f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0303e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01820] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03040] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01821] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03042] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01822] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03044] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01823] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03046] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01824] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03048] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01825] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0304a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01826] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0304c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01827] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0304e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01828] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03050] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01829] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03052] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0182a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03054] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0182b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03056] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0182c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03058] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0182d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0305a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0182e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0305c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0182f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0305e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01830] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03060] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01831] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03062] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01832] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03064] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01833] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03066] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01834] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03068] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01835] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0306a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01836] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0306c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01837] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0306e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01838] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03070] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01839] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03072] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0183a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03074] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0183b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03076] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0183c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03078] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0183d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0307a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0183e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0307c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0183f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0307e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01840] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03080] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01841] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03082] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01842] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03084] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01843] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03086] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01844] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03088] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01845] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0308a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01846] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0308c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01847] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0308e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01848] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03090] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01849] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03092] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0184a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03094] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0184b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03096] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0184c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03098] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0184d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0309a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0184e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0309c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0184f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0309e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01850] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01851] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01852] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01853] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01854] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01855] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01856] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01857] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01858] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01859] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0185a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0185b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0185c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0185d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0185e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0185f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01860] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01861] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01862] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01863] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01864] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01865] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01866] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01867] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01868] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01869] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0186a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0186b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0186c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0186d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0186e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0186f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01870] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01871] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01872] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01873] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01874] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01875] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01876] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01877] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01878] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01879] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0187a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0187b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0187c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0187d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0187e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0187f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h030fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01880] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03100] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01881] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03102] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01882] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03104] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01883] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03106] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01884] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03108] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01885] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0310a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01886] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0310c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01887] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0310e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01888] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03110] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01889] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03112] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0188a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03114] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0188b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03116] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0188c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03118] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0188d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0311a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0188e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0311c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0188f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0311e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01890] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03120] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01891] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03122] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01892] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03124] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01893] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03126] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01894] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03128] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01895] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0312a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01896] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0312c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01897] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0312e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01898] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03130] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01899] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03132] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0189a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03134] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0189b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03136] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0189c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03138] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0189d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0313a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0189e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0313c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0189f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0313e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03140] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03142] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03144] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03146] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03148] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0314a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0314c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0314e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03150] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03152] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03154] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03156] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03158] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0315a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0315c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0315e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03160] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03162] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03164] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03166] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03168] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0316a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0316c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0316e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03170] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03172] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03174] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03176] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03178] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0317a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0317c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0317e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03180] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03182] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03184] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03186] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03188] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0318a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0318c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0318e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03190] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03192] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03194] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03196] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03198] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0319a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0319c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0319e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h018ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h031fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01900] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03200] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01901] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03202] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01902] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03204] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01903] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03206] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01904] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03208] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01905] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0320a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01906] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0320c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01907] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0320e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01908] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03210] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01909] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03212] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0190a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03214] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0190b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03216] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0190c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03218] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0190d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0321a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0190e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0321c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0190f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0321e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01910] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03220] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01911] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03222] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01912] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03224] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01913] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03226] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01914] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03228] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01915] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0322a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01916] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0322c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01917] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0322e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01918] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03230] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01919] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03232] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0191a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03234] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0191b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03236] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0191c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03238] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0191d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0323a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0191e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0323c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0191f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0323e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01920] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03240] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01921] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03242] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01922] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03244] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01923] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03246] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01924] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03248] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01925] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0324a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01926] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0324c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01927] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0324e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01928] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03250] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01929] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03252] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0192a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03254] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0192b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03256] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0192c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03258] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0192d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0325a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0192e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0325c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0192f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0325e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01930] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03260] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01931] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03262] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01932] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03264] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01933] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03266] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01934] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03268] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01935] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0326a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01936] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0326c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01937] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0326e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01938] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03270] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01939] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03272] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0193a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03274] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0193b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03276] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0193c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03278] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0193d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0327a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0193e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0327c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0193f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0327e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01940] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03280] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01941] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03282] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01942] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03284] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01943] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03286] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01944] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03288] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01945] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0328a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01946] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0328c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01947] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0328e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01948] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03290] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01949] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03292] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0194a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03294] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0194b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03296] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0194c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03298] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0194d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0329a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0194e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0329c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0194f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0329e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01950] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01951] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01952] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01953] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01954] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01955] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01956] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01957] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01958] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01959] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0195a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0195b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0195c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0195d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0195e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0195f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01960] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01961] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01962] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01963] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01964] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01965] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01966] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01967] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01968] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01969] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0196a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0196b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0196c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0196d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0196e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0196f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01970] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01971] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01972] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01973] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01974] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01975] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01976] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01977] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01978] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01979] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0197a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0197b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0197c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0197d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0197e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0197f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h032fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01980] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03300] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01981] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03302] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01982] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03304] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01983] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03306] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01984] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03308] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01985] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0330a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01986] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0330c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01987] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0330e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01988] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03310] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01989] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03312] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0198a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03314] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0198b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03316] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0198c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03318] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0198d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0331a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0198e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0331c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0198f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0331e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01990] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03320] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01991] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03322] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01992] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03324] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01993] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03326] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01994] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03328] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01995] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0332a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01996] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0332c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01997] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0332e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01998] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03330] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01999] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03332] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0199a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03334] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0199b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03336] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0199c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03338] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0199d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0333a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0199e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0333c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0199f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0333e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03340] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03342] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03344] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03346] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03348] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0334a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0334c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0334e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03350] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03352] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03354] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03356] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03358] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0335a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0335c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0335e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03360] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03362] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03364] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03366] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03368] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0336a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0336c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0336e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03370] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03372] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03374] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03376] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03378] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0337a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0337c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0337e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03380] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03382] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03384] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03386] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03388] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0338a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0338c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0338e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03390] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03392] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03394] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03396] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03398] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0339a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0339c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0339e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h019ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h033fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03400] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03402] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03404] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03406] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03408] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0340a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0340c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0340e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03410] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03412] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03414] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03416] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03418] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0341a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0341c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0341e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03420] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03422] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03424] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03426] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03428] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0342a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0342c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0342e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03430] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03432] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03434] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03436] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03438] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0343a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0343c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0343e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03440] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03442] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03444] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03446] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03448] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0344a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0344c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0344e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03450] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03452] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03454] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03456] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03458] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0345a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0345c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0345e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03460] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03462] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03464] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03466] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03468] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0346a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0346c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0346e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03470] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03472] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03474] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03476] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03478] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0347a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0347c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0347e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03480] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03482] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03484] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03486] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03488] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0348a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0348c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0348e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03490] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03492] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03494] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03496] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03498] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0349a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0349c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0349e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h034fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03500] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03502] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03504] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03506] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03508] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0350a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0350c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0350e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03510] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03512] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03514] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03516] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03518] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0351a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0351c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0351e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03520] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03522] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03524] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03526] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03528] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0352a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0352c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0352e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03530] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03532] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03534] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03536] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03538] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0353a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0353c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01a9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0353e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aa0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03540] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aa1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03542] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aa2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03544] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aa3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03546] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aa4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03548] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aa5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0354a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aa6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0354c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aa7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0354e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aa8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03550] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aa9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03552] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aaa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03554] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03556] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03558] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0355a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0355c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aaf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0355e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ab0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03560] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ab1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03562] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ab2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03564] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ab3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03566] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ab4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03568] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ab5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0356a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ab6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0356c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ab7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0356e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ab8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03570] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ab9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03572] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03574] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01abb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03576] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01abc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03578] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01abd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0357a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01abe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0357c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01abf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0357e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ac0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03580] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ac1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03582] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ac2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03584] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ac3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03586] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ac4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03588] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ac5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0358a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ac6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0358c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ac7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0358e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ac8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03590] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ac9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03592] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03594] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01acb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03596] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01acc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03598] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01acd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0359a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ace] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0359c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01acf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0359e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ad0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ad1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ad2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ad3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ad4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ad5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ad6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ad7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ad8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ad9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ada] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01adb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01adc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01add] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ade] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01adf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ae0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ae1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ae2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ae3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ae4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ae5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ae6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ae7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ae8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ae9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aeb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01af0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01af1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01af2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01af3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01af4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01af5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01af6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01af7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01af8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01af9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01afa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01afb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01afc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01afd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01afe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01aff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h035fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03600] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03602] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03604] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03606] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03608] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0360a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0360c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0360e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03610] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03612] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03614] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03616] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03618] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0361a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0361c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0361e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03620] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03622] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03624] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03626] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03628] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0362a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0362c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0362e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03630] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03632] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03634] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03636] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03638] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0363a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0363c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0363e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03640] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03642] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03644] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03646] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03648] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0364a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0364c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0364e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03650] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03652] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03654] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03656] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03658] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0365a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0365c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0365e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03660] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03662] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03664] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03666] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03668] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0366a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0366c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0366e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03670] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03672] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03674] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03676] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03678] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0367a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0367c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0367e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03680] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03682] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03684] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03686] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03688] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0368a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0368c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0368e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03690] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03692] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03694] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03696] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03698] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0369a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0369c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0369e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h036fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03700] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03702] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03704] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03706] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03708] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0370a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0370c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0370e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03710] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03712] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03714] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03716] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03718] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0371a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0371c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0371e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03720] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03722] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03724] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03726] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03728] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0372a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0372c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0372e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03730] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03732] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03734] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03736] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03738] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0373a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0373c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01b9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0373e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ba0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03740] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ba1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03742] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ba2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03744] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ba3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03746] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ba4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03748] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ba5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0374a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ba6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0374c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ba7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0374e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ba8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03750] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ba9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03752] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01baa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03754] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03756] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03758] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0375a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0375c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01baf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0375e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03760] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03762] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03764] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03766] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03768] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0376a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0376c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0376e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03770] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03772] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03774] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03776] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03778] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0377a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0377c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0377e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03780] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03782] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03784] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03786] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03788] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0378a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0378c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0378e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03790] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03792] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03794] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03796] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03798] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0379a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0379c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0379e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01be0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01be1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01be2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01be3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01be4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01be5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01be6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01be7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01be8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01be9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01beb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bf0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bf1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bf2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bf3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bf4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bf5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bf6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bf7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bf8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bf9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01bff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h037fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03800] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03802] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03804] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03806] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03808] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0380a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0380c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0380e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03810] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03812] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03814] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03816] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03818] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0381a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0381c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0381e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03820] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03822] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03824] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03826] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03828] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0382a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0382c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0382e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03830] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03832] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03834] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03836] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03838] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0383a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0383c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0383e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03840] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03842] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03844] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03846] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03848] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0384a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0384c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0384e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03850] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03852] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03854] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03856] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03858] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0385a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0385c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0385e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03860] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03862] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03864] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03866] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03868] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0386a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0386c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0386e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03870] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03872] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03874] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03876] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03878] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0387a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0387c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0387e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03880] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03882] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03884] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03886] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03888] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0388a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0388c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0388e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03890] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03892] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03894] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03896] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03898] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0389a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0389c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0389e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h038fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03900] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03902] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03904] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03906] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03908] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0390a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0390c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0390e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03910] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03912] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03914] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03916] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03918] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0391a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0391c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0391e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03920] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03922] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03924] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03926] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03928] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0392a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0392c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0392e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03930] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03932] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03934] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03936] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03938] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0393a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0393c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01c9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0393e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ca0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03940] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ca1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03942] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ca2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03944] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ca3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03946] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ca4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03948] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ca5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0394a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ca6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0394c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ca7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0394e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ca8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03950] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ca9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03952] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01caa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03954] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03956] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03958] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0395a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0395c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01caf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0395e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03960] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03962] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03964] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03966] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03968] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0396a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0396c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0396e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03970] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03972] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03974] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03976] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03978] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0397a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0397c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0397e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03980] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03982] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03984] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03986] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03988] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0398a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0398c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0398e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03990] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03992] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03994] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ccb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03996] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ccc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03998] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ccd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0399a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0399c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ccf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0399e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ce0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ce1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ce2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ce3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ce4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ce5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ce6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ce7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ce8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ce9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ceb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ced] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cf0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cf1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cf2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cf3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cf4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cf5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cf6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cf7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cf8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cf9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01cff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h039fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03a9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ab0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ab2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ab4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ab6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ab8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03abc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03abe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ac0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ac2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ac4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ac6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ac8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03acc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ace] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ad0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ad2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ad4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ad6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ad8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ada] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03adc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ade] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ae0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ae2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ae4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ae6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ae8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03aee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03af0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03af2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03af4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03af6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03af8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03afa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03afc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03afe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01d9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01da0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01da1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01da2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01da3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01da4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01da5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01da6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01da7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01da8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01da9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01daa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01daf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01db0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01db1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01db2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01db3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01db4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01db5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01db6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01db7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01db8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01db9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03b9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ba0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ba2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ba4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ba6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ba8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03baa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ddb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ddc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ddd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ddf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01de0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01de1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01de2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01de3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01de4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01de5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01de6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01de7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01de8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01de9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01deb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ded] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01def] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01df0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03be0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01df1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03be2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01df2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03be4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01df3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03be6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01df4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03be8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01df5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01df6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01df7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01df8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01df9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01dff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03bfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03c9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ca0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ca2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ca4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ca6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ca8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03caa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ccc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ce0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ce2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ce4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ce6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ce8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03cfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01e9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ea0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ea1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ea2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ea3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ea4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ea5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ea6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ea7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ea8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ea9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eaa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ead] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eaf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ebb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ebc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ebd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ebe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ebf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ec0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ec1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ec2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ec3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ec4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ec5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ec6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ec7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ec8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ec9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ecb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ecc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ecd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ece] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ecf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03d9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ed0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03da0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ed1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03da2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ed2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03da4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ed3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03da6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ed4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03da8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ed5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03daa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ed6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ed7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ed8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03db0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ed9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03db2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03db4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01edb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03db6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01edc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03db8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01edd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ede] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01edf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ee0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ee1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ee2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ee3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ee4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ee5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ee6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ee7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ee8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ee9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eeb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ddc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ef0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03de0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ef1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03de2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ef2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03de4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ef3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03de6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ef4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03de8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ef5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ef6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ef7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ef8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03df0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ef9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03df2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01efa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03df4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01efb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03df6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01efc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03df8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01efd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01efe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01eff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03dfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03e9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ea0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ea2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ea4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ea6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ea8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ebc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ebe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ec0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ec2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ec4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ec6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ec8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ecc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ece] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ed0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ed2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ed4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ed6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ed8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03edc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ede] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ee0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ee2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ee4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ee6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ee8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03eee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ef0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ef2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ef4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ef6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ef8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03efa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03efc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03efe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01f9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fa0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fa1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fa2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fa3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fa4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fa5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fa6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fa7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fa8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fa9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01faa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01faf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03f9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03faa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fe0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fe1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fe2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fe3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fe4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fe5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fe6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fe7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fe8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fe9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01feb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ff0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fe0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ff1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fe2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ff2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fe4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ff3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fe6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ff4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fe8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ff5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ff6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ff7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03fee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ff8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ff0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ff9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ff2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ffa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ff4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ffb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ff6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ffc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ff8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ffd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ffa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01ffe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ffc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h01fff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h03ffe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02000] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04000] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02001] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04002] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02002] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04004] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02003] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04006] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02004] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04008] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02005] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0400a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02006] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0400c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02007] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0400e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02008] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04010] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02009] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04012] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0200a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04014] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0200b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04016] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0200c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04018] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0200d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0401a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0200e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0401c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0200f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0401e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02010] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04020] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02011] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04022] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02012] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04024] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02013] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04026] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02014] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04028] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02015] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0402a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02016] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0402c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02017] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0402e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02018] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04030] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02019] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04032] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0201a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04034] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0201b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04036] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0201c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04038] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0201d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0403a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0201e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0403c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0201f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0403e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02020] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04040] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02021] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04042] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02022] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04044] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02023] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04046] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02024] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04048] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02025] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0404a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02026] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0404c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02027] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0404e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02028] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04050] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02029] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04052] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0202a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04054] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0202b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04056] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0202c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04058] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0202d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0405a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0202e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0405c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0202f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0405e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02030] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04060] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02031] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04062] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02032] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04064] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02033] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04066] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02034] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04068] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02035] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0406a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02036] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0406c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02037] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0406e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02038] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04070] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02039] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04072] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0203a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04074] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0203b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04076] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0203c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04078] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0203d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0407a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0203e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0407c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0203f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0407e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02040] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04080] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02041] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04082] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02042] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04084] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02043] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04086] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02044] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04088] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02045] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0408a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02046] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0408c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02047] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0408e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02048] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04090] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02049] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04092] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0204a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04094] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0204b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04096] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0204c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04098] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0204d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0409a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0204e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0409c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0204f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0409e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02050] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02051] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02052] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02053] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02054] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02055] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02056] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02057] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02058] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02059] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0205a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0205b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0205c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0205d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0205e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0205f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02060] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02061] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02062] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02063] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02064] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02065] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02066] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02067] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02068] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02069] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0206a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0206b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0206c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0206d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0206e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0206f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02070] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02071] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02072] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02073] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02074] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02075] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02076] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02077] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02078] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02079] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0207a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0207b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0207c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0207d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0207e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0207f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h040fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02080] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04100] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02081] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04102] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02082] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04104] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02083] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04106] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02084] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04108] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02085] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0410a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02086] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0410c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02087] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0410e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02088] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04110] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02089] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04112] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0208a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04114] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0208b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04116] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0208c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04118] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0208d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0411a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0208e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0411c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0208f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0411e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02090] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04120] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02091] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04122] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02092] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04124] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02093] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04126] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02094] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04128] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02095] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0412a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02096] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0412c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02097] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0412e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02098] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04130] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02099] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04132] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0209a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04134] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0209b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04136] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0209c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04138] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0209d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0413a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0209e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0413c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0209f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0413e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04140] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04142] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04144] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04146] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04148] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0414a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0414c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0414e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04150] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04152] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04154] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04156] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04158] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0415a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0415c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0415e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04160] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04162] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04164] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04166] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04168] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0416a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0416c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0416e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04170] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04172] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04174] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04176] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04178] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0417a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0417c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0417e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04180] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04182] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04184] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04186] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04188] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0418a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0418c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0418e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04190] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04192] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04194] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04196] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04198] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0419a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0419c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0419e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h020ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h041fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02100] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04200] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02101] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04202] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02102] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04204] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02103] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04206] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02104] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04208] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02105] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0420a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02106] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0420c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02107] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0420e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02108] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04210] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02109] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04212] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0210a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04214] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0210b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04216] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0210c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04218] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0210d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0421a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0210e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0421c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0210f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0421e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02110] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04220] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02111] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04222] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02112] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04224] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02113] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04226] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02114] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04228] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02115] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0422a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02116] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0422c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02117] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0422e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02118] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04230] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02119] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04232] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0211a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04234] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0211b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04236] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0211c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04238] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0211d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0423a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0211e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0423c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0211f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0423e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02120] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04240] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02121] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04242] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02122] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04244] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02123] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04246] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02124] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04248] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02125] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0424a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02126] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0424c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02127] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0424e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02128] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04250] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02129] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04252] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0212a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04254] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0212b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04256] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0212c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04258] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0212d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0425a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0212e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0425c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0212f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0425e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02130] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04260] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02131] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04262] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02132] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04264] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02133] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04266] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02134] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04268] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02135] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0426a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02136] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0426c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02137] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0426e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02138] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04270] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02139] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04272] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0213a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04274] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0213b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04276] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0213c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04278] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0213d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0427a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0213e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0427c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0213f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0427e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02140] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04280] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02141] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04282] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02142] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04284] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02143] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04286] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02144] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04288] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02145] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0428a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02146] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0428c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02147] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0428e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02148] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04290] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02149] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04292] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0214a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04294] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0214b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04296] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0214c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04298] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0214d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0429a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0214e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0429c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0214f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0429e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02150] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02151] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02152] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02153] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02154] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02155] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02156] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02157] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02158] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02159] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0215a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0215b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0215c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0215d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0215e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0215f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02160] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02161] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02162] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02163] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02164] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02165] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02166] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02167] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02168] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02169] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0216a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0216b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0216c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0216d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0216e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0216f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02170] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02171] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02172] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02173] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02174] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02175] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02176] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02177] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02178] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02179] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0217a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0217b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0217c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0217d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0217e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0217f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h042fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02180] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04300] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02181] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04302] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02182] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04304] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02183] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04306] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02184] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04308] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02185] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0430a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02186] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0430c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02187] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0430e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02188] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04310] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02189] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04312] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0218a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04314] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0218b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04316] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0218c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04318] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0218d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0431a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0218e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0431c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0218f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0431e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02190] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04320] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02191] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04322] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02192] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04324] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02193] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04326] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02194] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04328] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02195] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0432a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02196] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0432c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02197] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0432e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02198] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04330] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02199] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04332] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0219a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04334] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0219b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04336] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0219c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04338] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0219d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0433a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0219e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0433c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0219f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0433e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04340] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04342] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04344] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04346] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04348] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0434a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0434c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0434e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04350] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04352] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04354] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04356] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04358] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0435a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0435c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0435e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04360] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04362] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04364] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04366] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04368] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0436a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0436c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0436e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04370] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04372] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04374] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04376] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04378] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0437a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0437c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0437e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04380] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04382] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04384] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04386] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04388] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0438a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0438c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0438e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04390] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04392] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04394] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04396] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04398] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0439a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0439c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0439e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h021ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h043fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02200] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04400] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02201] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04402] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02202] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04404] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02203] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04406] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02204] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04408] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02205] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0440a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02206] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0440c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02207] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0440e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02208] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04410] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02209] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04412] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0220a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04414] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0220b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04416] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0220c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04418] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0220d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0441a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0220e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0441c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0220f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0441e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02210] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04420] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02211] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04422] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02212] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04424] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02213] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04426] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02214] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04428] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02215] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0442a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02216] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0442c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02217] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0442e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02218] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04430] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02219] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04432] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0221a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04434] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0221b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04436] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0221c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04438] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0221d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0443a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0221e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0443c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0221f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0443e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02220] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04440] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02221] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04442] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02222] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04444] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02223] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04446] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02224] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04448] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02225] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0444a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02226] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0444c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02227] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0444e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02228] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04450] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02229] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04452] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0222a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04454] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0222b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04456] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0222c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04458] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0222d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0445a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0222e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0445c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0222f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0445e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02230] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04460] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02231] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04462] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02232] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04464] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02233] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04466] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02234] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04468] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02235] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0446a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02236] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0446c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02237] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0446e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02238] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04470] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02239] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04472] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0223a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04474] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0223b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04476] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0223c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04478] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0223d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0447a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0223e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0447c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0223f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0447e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02240] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04480] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02241] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04482] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02242] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04484] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02243] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04486] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02244] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04488] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02245] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0448a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02246] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0448c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02247] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0448e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02248] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04490] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02249] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04492] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0224a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04494] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0224b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04496] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0224c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04498] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0224d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0449a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0224e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0449c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0224f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0449e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02250] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02251] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02252] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02253] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02254] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02255] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02256] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02257] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02258] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02259] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0225a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0225b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0225c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0225d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0225e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0225f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02260] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02261] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02262] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02263] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02264] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02265] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02266] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02267] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02268] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02269] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0226a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0226b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0226c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0226d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0226e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0226f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02270] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02271] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02272] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02273] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02274] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02275] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02276] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02277] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02278] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02279] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0227a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0227b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0227c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0227d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0227e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0227f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h044fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02280] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04500] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02281] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04502] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02282] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04504] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02283] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04506] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02284] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04508] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02285] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0450a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02286] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0450c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02287] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0450e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02288] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04510] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02289] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04512] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0228a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04514] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0228b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04516] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0228c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04518] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0228d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0451a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0228e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0451c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0228f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0451e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02290] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04520] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02291] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04522] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02292] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04524] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02293] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04526] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02294] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04528] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02295] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0452a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02296] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0452c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02297] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0452e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02298] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04530] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02299] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04532] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0229a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04534] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0229b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04536] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0229c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04538] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0229d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0453a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0229e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0453c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0229f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0453e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04540] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04542] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04544] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04546] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04548] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0454a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0454c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0454e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04550] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04552] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04554] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04556] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04558] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0455a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0455c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0455e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04560] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04562] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04564] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04566] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04568] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0456a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0456c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0456e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04570] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04572] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04574] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04576] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04578] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0457a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0457c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0457e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04580] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04582] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04584] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04586] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04588] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0458a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0458c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0458e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04590] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04592] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04594] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04596] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04598] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0459a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0459c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0459e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h022ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h045fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02300] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04600] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02301] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04602] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02302] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04604] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02303] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04606] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02304] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04608] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02305] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0460a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02306] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0460c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02307] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0460e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02308] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04610] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02309] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04612] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0230a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04614] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0230b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04616] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0230c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04618] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0230d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0461a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0230e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0461c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0230f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0461e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02310] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04620] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02311] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04622] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02312] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04624] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02313] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04626] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02314] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04628] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02315] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0462a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02316] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0462c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02317] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0462e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02318] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04630] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02319] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04632] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0231a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04634] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0231b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04636] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0231c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04638] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0231d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0463a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0231e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0463c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0231f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0463e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02320] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04640] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02321] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04642] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02322] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04644] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02323] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04646] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02324] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04648] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02325] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0464a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02326] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0464c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02327] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0464e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02328] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04650] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02329] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04652] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0232a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04654] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0232b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04656] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0232c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04658] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0232d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0465a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0232e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0465c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0232f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0465e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02330] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04660] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02331] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04662] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02332] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04664] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02333] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04666] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02334] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04668] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02335] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0466a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02336] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0466c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02337] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0466e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02338] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04670] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02339] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04672] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0233a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04674] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0233b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04676] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0233c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04678] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0233d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0467a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0233e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0467c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0233f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0467e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02340] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04680] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02341] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04682] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02342] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04684] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02343] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04686] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02344] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04688] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02345] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0468a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02346] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0468c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02347] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0468e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02348] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04690] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02349] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04692] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0234a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04694] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0234b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04696] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0234c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04698] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0234d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0469a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0234e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0469c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0234f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0469e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02350] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02351] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02352] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02353] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02354] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02355] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02356] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02357] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02358] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02359] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0235a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0235b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0235c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0235d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0235e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0235f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02360] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02361] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02362] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02363] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02364] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02365] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02366] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02367] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02368] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02369] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0236a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0236b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0236c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0236d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0236e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0236f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02370] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02371] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02372] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02373] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02374] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02375] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02376] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02377] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02378] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02379] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0237a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0237b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0237c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0237d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0237e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0237f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h046fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02380] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04700] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02381] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04702] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02382] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04704] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02383] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04706] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02384] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04708] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02385] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0470a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02386] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0470c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02387] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0470e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02388] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04710] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02389] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04712] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0238a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04714] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0238b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04716] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0238c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04718] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0238d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0471a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0238e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0471c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0238f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0471e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02390] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04720] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02391] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04722] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02392] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04724] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02393] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04726] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02394] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04728] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02395] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0472a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02396] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0472c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02397] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0472e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02398] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04730] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02399] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04732] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0239a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04734] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0239b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04736] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0239c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04738] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0239d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0473a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0239e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0473c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0239f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0473e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04740] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04742] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04744] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04746] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04748] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0474a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0474c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0474e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04750] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04752] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04754] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04756] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04758] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0475a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0475c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0475e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04760] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04762] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04764] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04766] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04768] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0476a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0476c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0476e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04770] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04772] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04774] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04776] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04778] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0477a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0477c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0477e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04780] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04782] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04784] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04786] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04788] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0478a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0478c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0478e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04790] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04792] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04794] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04796] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04798] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0479a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0479c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0479e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h023ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h047fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02400] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04800] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02401] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04802] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02402] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04804] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02403] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04806] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02404] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04808] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02405] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0480a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02406] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0480c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02407] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0480e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02408] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04810] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02409] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04812] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0240a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04814] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0240b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04816] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0240c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04818] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0240d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0481a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0240e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0481c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0240f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0481e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02410] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04820] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02411] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04822] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02412] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04824] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02413] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04826] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02414] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04828] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02415] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0482a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02416] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0482c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02417] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0482e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02418] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04830] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02419] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04832] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0241a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04834] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0241b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04836] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0241c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04838] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0241d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0483a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0241e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0483c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0241f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0483e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02420] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04840] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02421] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04842] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02422] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04844] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02423] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04846] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02424] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04848] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02425] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0484a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02426] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0484c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02427] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0484e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02428] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04850] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02429] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04852] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0242a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04854] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0242b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04856] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0242c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04858] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0242d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0485a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0242e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0485c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0242f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0485e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02430] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04860] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02431] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04862] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02432] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04864] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02433] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04866] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02434] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04868] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02435] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0486a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02436] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0486c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02437] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0486e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02438] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04870] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02439] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04872] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0243a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04874] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0243b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04876] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0243c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04878] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0243d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0487a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0243e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0487c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0243f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0487e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02440] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04880] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02441] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04882] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02442] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04884] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02443] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04886] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02444] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04888] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02445] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0488a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02446] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0488c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02447] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0488e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02448] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04890] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02449] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04892] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0244a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04894] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0244b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04896] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0244c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04898] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0244d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0489a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0244e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0489c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0244f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0489e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02450] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02451] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02452] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02453] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02454] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02455] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02456] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02457] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02458] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02459] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0245a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0245b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0245c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0245d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0245e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0245f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02460] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02461] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02462] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02463] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02464] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02465] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02466] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02467] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02468] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02469] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0246a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0246b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0246c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0246d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0246e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0246f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02470] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02471] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02472] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02473] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02474] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02475] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02476] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02477] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02478] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02479] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0247a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0247b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0247c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0247d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0247e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0247f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h048fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02480] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04900] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02481] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04902] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02482] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04904] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02483] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04906] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02484] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04908] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02485] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0490a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02486] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0490c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02487] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0490e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02488] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04910] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02489] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04912] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0248a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04914] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0248b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04916] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0248c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04918] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0248d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0491a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0248e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0491c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0248f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0491e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02490] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04920] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02491] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04922] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02492] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04924] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02493] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04926] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02494] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04928] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02495] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0492a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02496] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0492c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02497] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0492e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02498] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04930] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02499] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04932] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0249a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04934] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0249b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04936] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0249c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04938] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0249d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0493a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0249e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0493c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0249f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0493e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04940] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04942] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04944] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04946] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04948] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0494a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0494c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0494e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04950] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04952] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04954] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04956] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04958] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0495a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0495c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0495e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04960] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04962] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04964] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04966] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04968] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0496a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0496c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0496e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04970] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04972] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04974] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04976] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04978] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0497a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0497c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0497e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04980] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04982] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04984] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04986] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04988] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0498a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0498c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0498e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04990] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04992] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04994] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04996] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04998] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0499a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0499c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0499e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h024ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h049fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02500] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02501] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02502] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02503] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02504] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02505] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02506] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02507] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02508] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02509] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0250a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0250b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0250c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0250d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0250e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0250f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02510] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02511] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02512] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02513] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02514] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02515] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02516] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02517] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02518] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02519] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0251a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0251b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0251c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0251d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0251e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0251f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02520] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02521] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02522] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02523] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02524] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02525] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02526] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02527] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02528] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02529] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0252a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0252b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0252c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0252d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0252e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0252f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02530] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02531] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02532] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02533] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02534] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02535] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02536] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02537] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02538] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02539] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0253a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0253b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0253c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0253d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0253e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0253f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02540] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02541] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02542] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02543] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02544] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02545] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02546] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02547] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02548] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02549] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0254a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0254b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0254c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0254d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0254e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0254f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04a9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02550] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02551] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02552] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02553] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02554] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02555] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02556] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02557] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02558] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ab0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02559] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ab2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0255a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ab4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0255b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ab6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0255c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ab8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0255d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0255e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04abc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0255f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04abe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02560] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ac0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02561] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ac2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02562] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ac4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02563] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ac6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02564] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ac8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02565] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02566] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04acc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02567] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ace] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02568] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ad0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02569] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ad2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0256a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ad4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0256b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ad6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0256c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ad8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0256d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ada] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0256e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04adc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0256f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ade] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02570] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ae0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02571] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ae2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02572] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ae4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02573] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ae6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02574] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ae8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02575] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02576] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02577] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04aee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02578] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04af0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02579] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04af2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0257a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04af4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0257b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04af6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0257c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04af8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0257d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04afa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0257e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04afc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0257f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04afe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02580] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02581] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02582] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02583] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02584] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02585] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02586] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02587] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02588] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02589] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0258a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0258b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0258c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0258d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0258e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0258f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02590] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02591] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02592] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02593] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02594] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02595] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02596] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02597] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02598] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02599] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0259a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0259b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0259c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0259d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0259e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0259f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04b9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ba0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ba2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ba4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ba6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ba8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04baa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04be0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04be2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04be4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04be6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04be8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h025ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04bfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02600] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02601] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02602] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02603] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02604] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02605] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02606] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02607] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02608] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02609] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0260a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0260b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0260c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0260d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0260e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0260f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02610] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02611] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02612] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02613] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02614] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02615] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02616] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02617] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02618] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02619] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0261a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0261b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0261c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0261d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0261e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0261f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02620] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02621] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02622] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02623] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02624] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02625] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02626] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02627] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02628] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02629] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0262a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0262b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0262c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0262d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0262e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0262f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02630] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02631] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02632] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02633] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02634] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02635] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02636] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02637] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02638] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02639] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0263a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0263b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0263c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0263d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0263e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0263f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02640] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02641] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02642] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02643] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02644] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02645] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02646] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02647] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02648] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02649] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0264a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0264b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0264c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0264d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0264e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0264f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04c9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02650] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ca0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02651] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ca2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02652] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ca4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02653] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ca6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02654] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ca8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02655] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04caa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02656] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02657] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02658] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02659] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0265a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0265b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0265c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0265d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0265e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0265f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02660] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02661] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02662] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02663] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02664] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02665] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02666] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ccc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02667] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02668] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02669] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0266a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0266b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0266c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0266d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0266e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0266f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02670] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ce0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02671] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ce2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02672] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ce4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02673] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ce6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02674] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ce8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02675] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02676] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02677] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02678] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02679] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0267a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0267b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0267c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0267d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0267e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0267f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04cfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02680] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02681] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02682] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02683] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02684] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02685] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02686] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02687] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02688] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02689] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0268a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0268b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0268c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0268d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0268e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0268f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02690] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02691] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02692] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02693] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02694] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02695] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02696] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02697] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02698] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02699] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0269a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0269b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0269c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0269d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0269e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0269f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04d9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04da0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04da2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04da4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04da6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04da8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04daa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04db0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04db2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04db4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04db6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04db8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ddc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04de0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04de2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04de4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04de6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04de8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04df0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04df2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04df4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04df6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04df8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h026ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04dfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02700] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02701] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02702] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02703] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02704] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02705] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02706] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02707] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02708] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02709] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0270a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0270b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0270c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0270d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0270e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0270f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02710] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02711] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02712] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02713] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02714] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02715] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02716] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02717] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02718] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02719] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0271a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0271b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0271c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0271d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0271e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0271f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02720] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02721] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02722] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02723] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02724] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02725] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02726] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02727] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02728] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02729] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0272a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0272b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0272c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0272d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0272e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0272f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02730] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02731] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02732] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02733] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02734] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02735] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02736] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02737] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02738] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02739] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0273a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0273b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0273c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0273d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0273e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0273f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02740] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02741] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02742] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02743] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02744] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02745] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02746] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02747] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02748] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02749] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0274a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0274b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0274c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0274d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0274e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0274f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04e9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02750] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ea0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02751] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ea2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02752] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ea4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02753] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ea6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02754] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ea8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02755] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02756] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02757] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02758] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02759] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0275a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0275b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0275c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0275d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0275e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ebc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0275f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ebe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02760] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ec0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02761] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ec2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02762] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ec4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02763] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ec6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02764] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ec8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02765] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02766] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ecc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02767] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ece] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02768] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ed0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02769] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ed2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0276a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ed4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0276b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ed6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0276c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ed8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0276d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0276e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04edc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0276f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ede] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02770] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ee0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02771] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ee2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02772] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ee4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02773] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ee6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02774] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ee8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02775] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02776] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02777] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04eee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02778] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ef0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02779] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ef2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0277a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ef4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0277b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ef6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0277c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ef8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0277d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04efa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0277e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04efc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0277f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04efe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02780] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02781] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02782] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02783] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02784] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02785] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02786] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02787] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02788] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02789] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0278a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0278b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0278c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0278d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0278e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0278f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02790] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02791] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02792] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02793] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02794] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02795] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02796] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02797] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02798] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02799] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0279a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0279b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0279c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0279d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0279e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0279f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04f9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04faa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fe0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fe2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fe4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fe6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fe8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04fee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ff0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ff2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ff4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ff6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ff8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ffa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ffc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h027ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h04ffe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02800] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05000] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02801] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05002] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02802] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05004] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02803] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05006] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02804] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05008] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02805] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0500a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02806] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0500c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02807] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0500e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02808] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05010] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02809] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05012] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0280a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05014] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0280b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05016] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0280c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05018] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0280d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0501a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0280e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0501c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0280f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0501e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02810] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05020] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02811] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05022] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02812] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05024] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02813] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05026] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02814] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05028] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02815] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0502a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02816] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0502c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02817] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0502e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02818] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05030] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02819] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05032] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0281a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05034] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0281b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05036] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0281c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05038] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0281d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0503a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0281e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0503c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0281f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0503e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02820] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05040] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02821] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05042] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02822] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05044] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02823] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05046] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02824] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05048] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02825] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0504a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02826] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0504c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02827] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0504e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02828] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05050] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02829] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05052] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0282a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05054] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0282b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05056] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0282c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05058] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0282d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0505a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0282e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0505c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0282f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0505e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02830] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05060] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02831] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05062] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02832] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05064] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02833] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05066] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02834] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05068] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02835] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0506a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02836] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0506c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02837] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0506e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02838] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05070] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02839] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05072] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0283a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05074] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0283b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05076] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0283c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05078] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0283d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0507a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0283e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0507c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0283f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0507e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02840] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05080] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02841] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05082] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02842] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05084] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02843] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05086] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02844] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05088] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02845] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0508a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02846] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0508c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02847] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0508e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02848] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05090] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02849] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05092] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0284a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05094] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0284b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05096] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0284c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05098] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0284d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0509a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0284e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0509c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0284f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0509e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02850] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02851] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02852] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02853] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02854] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02855] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02856] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02857] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02858] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02859] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0285a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0285b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0285c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0285d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0285e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0285f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02860] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02861] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02862] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02863] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02864] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02865] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02866] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02867] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02868] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02869] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0286a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0286b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0286c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0286d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0286e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0286f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02870] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02871] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02872] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02873] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02874] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02875] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02876] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02877] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02878] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02879] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0287a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0287b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0287c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0287d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0287e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0287f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h050fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02880] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05100] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02881] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05102] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02882] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05104] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02883] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05106] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02884] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05108] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02885] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0510a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02886] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0510c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02887] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0510e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02888] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05110] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02889] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05112] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0288a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05114] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0288b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05116] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0288c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05118] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0288d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0511a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0288e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0511c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0288f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0511e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02890] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05120] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02891] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05122] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02892] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05124] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02893] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05126] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02894] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05128] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02895] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0512a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02896] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0512c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02897] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0512e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02898] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05130] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02899] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05132] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0289a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05134] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0289b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05136] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0289c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05138] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0289d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0513a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0289e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0513c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0289f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0513e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05140] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05142] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05144] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05146] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05148] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0514a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0514c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0514e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05150] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05152] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05154] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05156] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05158] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0515a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0515c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0515e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05160] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05162] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05164] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05166] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05168] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0516a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0516c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0516e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05170] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05172] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05174] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05176] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05178] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0517a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0517c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0517e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05180] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05182] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05184] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05186] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05188] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0518a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0518c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0518e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05190] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05192] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05194] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05196] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05198] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0519a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0519c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0519e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h028ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h051fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02900] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05200] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02901] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05202] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02902] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05204] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02903] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05206] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02904] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05208] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02905] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0520a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02906] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0520c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02907] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0520e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02908] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05210] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02909] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05212] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0290a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05214] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0290b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05216] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0290c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05218] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0290d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0521a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0290e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0521c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0290f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0521e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02910] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05220] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02911] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05222] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02912] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05224] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02913] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05226] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02914] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05228] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02915] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0522a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02916] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0522c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02917] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0522e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02918] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05230] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02919] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05232] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0291a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05234] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0291b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05236] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0291c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05238] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0291d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0523a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0291e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0523c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0291f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0523e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02920] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05240] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02921] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05242] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02922] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05244] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02923] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05246] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02924] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05248] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02925] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0524a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02926] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0524c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02927] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0524e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02928] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05250] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02929] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05252] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0292a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05254] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0292b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05256] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0292c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05258] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0292d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0525a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0292e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0525c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0292f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0525e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02930] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05260] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02931] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05262] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02932] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05264] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02933] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05266] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02934] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05268] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02935] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0526a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02936] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0526c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02937] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0526e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02938] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05270] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02939] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05272] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0293a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05274] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0293b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05276] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0293c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05278] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0293d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0527a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0293e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0527c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0293f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0527e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02940] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05280] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02941] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05282] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02942] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05284] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02943] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05286] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02944] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05288] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02945] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0528a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02946] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0528c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02947] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0528e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02948] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05290] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02949] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05292] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0294a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05294] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0294b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05296] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0294c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05298] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0294d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0529a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0294e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0529c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0294f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0529e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02950] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02951] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02952] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02953] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02954] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02955] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02956] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02957] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02958] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02959] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0295a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0295b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0295c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0295d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0295e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0295f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02960] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02961] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02962] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02963] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02964] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02965] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02966] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02967] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02968] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02969] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0296a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0296b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0296c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0296d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0296e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0296f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02970] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02971] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02972] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02973] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02974] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02975] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02976] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02977] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02978] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02979] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0297a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0297b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0297c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0297d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0297e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0297f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h052fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02980] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05300] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02981] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05302] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02982] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05304] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02983] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05306] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02984] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05308] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02985] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0530a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02986] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0530c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02987] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0530e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02988] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05310] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02989] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05312] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0298a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05314] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0298b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05316] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0298c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05318] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0298d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0531a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0298e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0531c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0298f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0531e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02990] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05320] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02991] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05322] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02992] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05324] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02993] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05326] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02994] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05328] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02995] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0532a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02996] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0532c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02997] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0532e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02998] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05330] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02999] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05332] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0299a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05334] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0299b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05336] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0299c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05338] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0299d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0533a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0299e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0533c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0299f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0533e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05340] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05342] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05344] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05346] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05348] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0534a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0534c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0534e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05350] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05352] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05354] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05356] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05358] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0535a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0535c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0535e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05360] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05362] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05364] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05366] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05368] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0536a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0536c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0536e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05370] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05372] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05374] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05376] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05378] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0537a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0537c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0537e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05380] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05382] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05384] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05386] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05388] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0538a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0538c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0538e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05390] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05392] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05394] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05396] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05398] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0539a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0539c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0539e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h029ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h053fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05400] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05402] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05404] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05406] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05408] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0540a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0540c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0540e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05410] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05412] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05414] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05416] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05418] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0541a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0541c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0541e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05420] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05422] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05424] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05426] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05428] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0542a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0542c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0542e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05430] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05432] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05434] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05436] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05438] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0543a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0543c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0543e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05440] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05442] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05444] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05446] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05448] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0544a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0544c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0544e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05450] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05452] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05454] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05456] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05458] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0545a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0545c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0545e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05460] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05462] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05464] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05466] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05468] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0546a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0546c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0546e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05470] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05472] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05474] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05476] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05478] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0547a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0547c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0547e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05480] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05482] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05484] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05486] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05488] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0548a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0548c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0548e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05490] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05492] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05494] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05496] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05498] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0549a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0549c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0549e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h054fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05500] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05502] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05504] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05506] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05508] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0550a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0550c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0550e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05510] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05512] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05514] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05516] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05518] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0551a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0551c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0551e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05520] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05522] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05524] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05526] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05528] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0552a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0552c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0552e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05530] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05532] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05534] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05536] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05538] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0553a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0553c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02a9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0553e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aa0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05540] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aa1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05542] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aa2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05544] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aa3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05546] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aa4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05548] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aa5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0554a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aa6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0554c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aa7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0554e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aa8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05550] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aa9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05552] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aaa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05554] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05556] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05558] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0555a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0555c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aaf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0555e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ab0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05560] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ab1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05562] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ab2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05564] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ab3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05566] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ab4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05568] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ab5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0556a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ab6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0556c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ab7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0556e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ab8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05570] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ab9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05572] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05574] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02abb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05576] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02abc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05578] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02abd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0557a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02abe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0557c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02abf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0557e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ac0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05580] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ac1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05582] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ac2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05584] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ac3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05586] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ac4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05588] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ac5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0558a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ac6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0558c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ac7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0558e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ac8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05590] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ac9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05592] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05594] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02acb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05596] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02acc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05598] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02acd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0559a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ace] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0559c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02acf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0559e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ad0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ad1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ad2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ad3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ad4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ad5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ad6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ad7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ad8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ad9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ada] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02adb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02adc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02add] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ade] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02adf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ae0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ae1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ae2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ae3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ae4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ae5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ae6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ae7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ae8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ae9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aeb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02af0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02af1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02af2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02af3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02af4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02af5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02af6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02af7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02af8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02af9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02afa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02afb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02afc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02afd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02afe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02aff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h055fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05600] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05602] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05604] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05606] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05608] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0560a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0560c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0560e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05610] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05612] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05614] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05616] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05618] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0561a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0561c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0561e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05620] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05622] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05624] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05626] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05628] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0562a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0562c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0562e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05630] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05632] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05634] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05636] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05638] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0563a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0563c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0563e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05640] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05642] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05644] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05646] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05648] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0564a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0564c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0564e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05650] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05652] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05654] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05656] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05658] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0565a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0565c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0565e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05660] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05662] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05664] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05666] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05668] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0566a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0566c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0566e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05670] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05672] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05674] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05676] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05678] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0567a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0567c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0567e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05680] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05682] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05684] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05686] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05688] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0568a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0568c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0568e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05690] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05692] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05694] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05696] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05698] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0569a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0569c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0569e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h056fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05700] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05702] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05704] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05706] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05708] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0570a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0570c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0570e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05710] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05712] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05714] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05716] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05718] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0571a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0571c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0571e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05720] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05722] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05724] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05726] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05728] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0572a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0572c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0572e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05730] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05732] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05734] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05736] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05738] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0573a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0573c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02b9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0573e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ba0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05740] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ba1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05742] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ba2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05744] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ba3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05746] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ba4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05748] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ba5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0574a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ba6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0574c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ba7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0574e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ba8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05750] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ba9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05752] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02baa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05754] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05756] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05758] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0575a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0575c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02baf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0575e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05760] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05762] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05764] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05766] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05768] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0576a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0576c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0576e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05770] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05772] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05774] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05776] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05778] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0577a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0577c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0577e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05780] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05782] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05784] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05786] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05788] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0578a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0578c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0578e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05790] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05792] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05794] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05796] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05798] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0579a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0579c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0579e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02be0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02be1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02be2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02be3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02be4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02be5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02be6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02be7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02be8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02be9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02beb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bf0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bf1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bf2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bf3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bf4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bf5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bf6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bf7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bf8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bf9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02bff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h057fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05800] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05802] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05804] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05806] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05808] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0580a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0580c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0580e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05810] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05812] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05814] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05816] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05818] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0581a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0581c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0581e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05820] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05822] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05824] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05826] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05828] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0582a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0582c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0582e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05830] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05832] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05834] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05836] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05838] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0583a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0583c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0583e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05840] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05842] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05844] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05846] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05848] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0584a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0584c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0584e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05850] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05852] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05854] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05856] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05858] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0585a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0585c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0585e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05860] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05862] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05864] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05866] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05868] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0586a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0586c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0586e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05870] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05872] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05874] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05876] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05878] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0587a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0587c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0587e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05880] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05882] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05884] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05886] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05888] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0588a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0588c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0588e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05890] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05892] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05894] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05896] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05898] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0589a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0589c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0589e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h058fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05900] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05902] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05904] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05906] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05908] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0590a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0590c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0590e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05910] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05912] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05914] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05916] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05918] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0591a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0591c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0591e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05920] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05922] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05924] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05926] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05928] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0592a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0592c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0592e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05930] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05932] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05934] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05936] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05938] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0593a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0593c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02c9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0593e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ca0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05940] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ca1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05942] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ca2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05944] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ca3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05946] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ca4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05948] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ca5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0594a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ca6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0594c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ca7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0594e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ca8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05950] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ca9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05952] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02caa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05954] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05956] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05958] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0595a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0595c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02caf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0595e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05960] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05962] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05964] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05966] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05968] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0596a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0596c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0596e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05970] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05972] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05974] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05976] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05978] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0597a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0597c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0597e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05980] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05982] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05984] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05986] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05988] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0598a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0598c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0598e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05990] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05992] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05994] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ccb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05996] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ccc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05998] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ccd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0599a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0599c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ccf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0599e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ce0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ce1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ce2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ce3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ce4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ce5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ce6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ce7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ce8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ce9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ceb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ced] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cf0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cf1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cf2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cf3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cf4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cf5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cf6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cf7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cf8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cf9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02cff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h059fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05a9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ab0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ab2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ab4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ab6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ab8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05abc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05abe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ac0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ac2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ac4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ac6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ac8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05acc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ace] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ad0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ad2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ad4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ad6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ad8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ada] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05adc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ade] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ae0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ae2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ae4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ae6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ae8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05aee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05af0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05af2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05af4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05af6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05af8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05afa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05afc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05afe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02d9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02da0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02da1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02da2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02da3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02da4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02da5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02da6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02da7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02da8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02da9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02daa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02daf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02db0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02db1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02db2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02db3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02db4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02db5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02db6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02db7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02db8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02db9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05b9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ba0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ba2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ba4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ba6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ba8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05baa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ddb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ddc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ddd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ddf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02de0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02de1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02de2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02de3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02de4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02de5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02de6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02de7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02de8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02de9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02deb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ded] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02def] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02df0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05be0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02df1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05be2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02df2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05be4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02df3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05be6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02df4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05be8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02df5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02df6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02df7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02df8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02df9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02dff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05bfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05c9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ca0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ca2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ca4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ca6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ca8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05caa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ccc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ce0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ce2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ce4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ce6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ce8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05cfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02e9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ea0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ea1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ea2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ea3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ea4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ea5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ea6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ea7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ea8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ea9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eaa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ead] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eaf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ebb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ebc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ebd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ebe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ebf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ec0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ec1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ec2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ec3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ec4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ec5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ec6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ec7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ec8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ec9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ecb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ecc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ecd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ece] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ecf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05d9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ed0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05da0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ed1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05da2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ed2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05da4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ed3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05da6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ed4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05da8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ed5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05daa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ed6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ed7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ed8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05db0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ed9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05db2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05db4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02edb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05db6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02edc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05db8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02edd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ede] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02edf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ee0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ee1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ee2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ee3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ee4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ee5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ee6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ee7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ee8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ee9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eeb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ddc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ef0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05de0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ef1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05de2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ef2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05de4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ef3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05de6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ef4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05de8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ef5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ef6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ef7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ef8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05df0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ef9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05df2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02efa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05df4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02efb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05df6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02efc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05df8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02efd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02efe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02eff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05dfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05e9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ea0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ea2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ea4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ea6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ea8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ebc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ebe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ec0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ec2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ec4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ec6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ec8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ecc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ece] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ed0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ed2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ed4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ed6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ed8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05edc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ede] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ee0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ee2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ee4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ee6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ee8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05eee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ef0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ef2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ef4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ef6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ef8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05efa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05efc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05efe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02f9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fa0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fa1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fa2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fa3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fa4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fa5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fa6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fa7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fa8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fa9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02faa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02faf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05f9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05faa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fe0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fe1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fe2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fe3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fe4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fe5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fe6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fe7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fe8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fe9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02feb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ff0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fe0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ff1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fe2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ff2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fe4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ff3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fe6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ff4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fe8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ff5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ff6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ff7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05fee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ff8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ff0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ff9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ff2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ffa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ff4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ffb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ff6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ffc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ff8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ffd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ffa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02ffe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ffc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h02fff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h05ffe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03000] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06000] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03001] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06002] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03002] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06004] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03003] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06006] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03004] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06008] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03005] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0600a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03006] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0600c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03007] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0600e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03008] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06010] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03009] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06012] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0300a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06014] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0300b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06016] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0300c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06018] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0300d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0601a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0300e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0601c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0300f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0601e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03010] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06020] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03011] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06022] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03012] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06024] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03013] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06026] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03014] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06028] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03015] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0602a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03016] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0602c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03017] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0602e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03018] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06030] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03019] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06032] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0301a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06034] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0301b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06036] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0301c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06038] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0301d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0603a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0301e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0603c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0301f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0603e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03020] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06040] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03021] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06042] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03022] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06044] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03023] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06046] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03024] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06048] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03025] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0604a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03026] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0604c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03027] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0604e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03028] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06050] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03029] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06052] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0302a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06054] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0302b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06056] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0302c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06058] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0302d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0605a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0302e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0605c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0302f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0605e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03030] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06060] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03031] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06062] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03032] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06064] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03033] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06066] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03034] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06068] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03035] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0606a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03036] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0606c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03037] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0606e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03038] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06070] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03039] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06072] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0303a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06074] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0303b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06076] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0303c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06078] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0303d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0607a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0303e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0607c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0303f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0607e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03040] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06080] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03041] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06082] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03042] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06084] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03043] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06086] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03044] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06088] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03045] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0608a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03046] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0608c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03047] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0608e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03048] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06090] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03049] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06092] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0304a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06094] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0304b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06096] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0304c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06098] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0304d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0609a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0304e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0609c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0304f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0609e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03050] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03051] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03052] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03053] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03054] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03055] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03056] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03057] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03058] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03059] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0305a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0305b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0305c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0305d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0305e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0305f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03060] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03061] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03062] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03063] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03064] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03065] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03066] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03067] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03068] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03069] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0306a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0306b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0306c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0306d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0306e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0306f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03070] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03071] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03072] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03073] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03074] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03075] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03076] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03077] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03078] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03079] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0307a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0307b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0307c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0307d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0307e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0307f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h060fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03080] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06100] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03081] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06102] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03082] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06104] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03083] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06106] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03084] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06108] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03085] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0610a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03086] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0610c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03087] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0610e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03088] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06110] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03089] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06112] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0308a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06114] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0308b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06116] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0308c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06118] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0308d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0611a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0308e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0611c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0308f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0611e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03090] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06120] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03091] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06122] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03092] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06124] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03093] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06126] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03094] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06128] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03095] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0612a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03096] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0612c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03097] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0612e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03098] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06130] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03099] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06132] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0309a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06134] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0309b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06136] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0309c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06138] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0309d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0613a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0309e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0613c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0309f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0613e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06140] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06142] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06144] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06146] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06148] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0614a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0614c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0614e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06150] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06152] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06154] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06156] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06158] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0615a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0615c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0615e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06160] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06162] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06164] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06166] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06168] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0616a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0616c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0616e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06170] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06172] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06174] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06176] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06178] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0617a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0617c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0617e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06180] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06182] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06184] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06186] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06188] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0618a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0618c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0618e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06190] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06192] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06194] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06196] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06198] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0619a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0619c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0619e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h030ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h061fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03100] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06200] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03101] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06202] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03102] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06204] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03103] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06206] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03104] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06208] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03105] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0620a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03106] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0620c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03107] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0620e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03108] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06210] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03109] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06212] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0310a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06214] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0310b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06216] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0310c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06218] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0310d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0621a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0310e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0621c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0310f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0621e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03110] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06220] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03111] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06222] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03112] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06224] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03113] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06226] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03114] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06228] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03115] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0622a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03116] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0622c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03117] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0622e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03118] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06230] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03119] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06232] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0311a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06234] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0311b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06236] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0311c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06238] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0311d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0623a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0311e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0623c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0311f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0623e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03120] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06240] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03121] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06242] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03122] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06244] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03123] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06246] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03124] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06248] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03125] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0624a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03126] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0624c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03127] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0624e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03128] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06250] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03129] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06252] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0312a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06254] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0312b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06256] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0312c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06258] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0312d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0625a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0312e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0625c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0312f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0625e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03130] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06260] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03131] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06262] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03132] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06264] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03133] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06266] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03134] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06268] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03135] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0626a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03136] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0626c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03137] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0626e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03138] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06270] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03139] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06272] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0313a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06274] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0313b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06276] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0313c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06278] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0313d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0627a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0313e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0627c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0313f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0627e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03140] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06280] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03141] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06282] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03142] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06284] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03143] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06286] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03144] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06288] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03145] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0628a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03146] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0628c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03147] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0628e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03148] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06290] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03149] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06292] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0314a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06294] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0314b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06296] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0314c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06298] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0314d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0629a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0314e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0629c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0314f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0629e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03150] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03151] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03152] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03153] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03154] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03155] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03156] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03157] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03158] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03159] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0315a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0315b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0315c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0315d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0315e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0315f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03160] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03161] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03162] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03163] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03164] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03165] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03166] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03167] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03168] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03169] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0316a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0316b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0316c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0316d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0316e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0316f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03170] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03171] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03172] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03173] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03174] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03175] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03176] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03177] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03178] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03179] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0317a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0317b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0317c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0317d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0317e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0317f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h062fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03180] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06300] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03181] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06302] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03182] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06304] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03183] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06306] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03184] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06308] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03185] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0630a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03186] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0630c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03187] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0630e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03188] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06310] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03189] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06312] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0318a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06314] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0318b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06316] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0318c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06318] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0318d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0631a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0318e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0631c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0318f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0631e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03190] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06320] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03191] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06322] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03192] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06324] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03193] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06326] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03194] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06328] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03195] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0632a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03196] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0632c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03197] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0632e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03198] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06330] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03199] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06332] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0319a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06334] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0319b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06336] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0319c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06338] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0319d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0633a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0319e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0633c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0319f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0633e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06340] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06342] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06344] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06346] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06348] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0634a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0634c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0634e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06350] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06352] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06354] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06356] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06358] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0635a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0635c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0635e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06360] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06362] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06364] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06366] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06368] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0636a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0636c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0636e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06370] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06372] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06374] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06376] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06378] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0637a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0637c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0637e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06380] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06382] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06384] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06386] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06388] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0638a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0638c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0638e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06390] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06392] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06394] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06396] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06398] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0639a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0639c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0639e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h031ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h063fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03200] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06400] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03201] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06402] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03202] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06404] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03203] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06406] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03204] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06408] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03205] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0640a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03206] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0640c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03207] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0640e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03208] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06410] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03209] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06412] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0320a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06414] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0320b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06416] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0320c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06418] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0320d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0641a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0320e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0641c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0320f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0641e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03210] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06420] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03211] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06422] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03212] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06424] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03213] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06426] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03214] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06428] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03215] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0642a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03216] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0642c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03217] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0642e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03218] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06430] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03219] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06432] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0321a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06434] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0321b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06436] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0321c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06438] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0321d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0643a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0321e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0643c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0321f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0643e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03220] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06440] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03221] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06442] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03222] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06444] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03223] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06446] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03224] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06448] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03225] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0644a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03226] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0644c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03227] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0644e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03228] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06450] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03229] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06452] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0322a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06454] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0322b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06456] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0322c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06458] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0322d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0645a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0322e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0645c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0322f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0645e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03230] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06460] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03231] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06462] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03232] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06464] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03233] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06466] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03234] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06468] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03235] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0646a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03236] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0646c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03237] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0646e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03238] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06470] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03239] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06472] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0323a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06474] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0323b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06476] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0323c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06478] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0323d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0647a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0323e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0647c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0323f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0647e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03240] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06480] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03241] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06482] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03242] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06484] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03243] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06486] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03244] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06488] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03245] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0648a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03246] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0648c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03247] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0648e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03248] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06490] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03249] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06492] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0324a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06494] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0324b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06496] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0324c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06498] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0324d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0649a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0324e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0649c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0324f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0649e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03250] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03251] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03252] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03253] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03254] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03255] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03256] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03257] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03258] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03259] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0325a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0325b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0325c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0325d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0325e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0325f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03260] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03261] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03262] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03263] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03264] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03265] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03266] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03267] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03268] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03269] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0326a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0326b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0326c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0326d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0326e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0326f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03270] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03271] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03272] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03273] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03274] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03275] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03276] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03277] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03278] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03279] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0327a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0327b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0327c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0327d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0327e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0327f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h064fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03280] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06500] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03281] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06502] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03282] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06504] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03283] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06506] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03284] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06508] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03285] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0650a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03286] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0650c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03287] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0650e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03288] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06510] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03289] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06512] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0328a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06514] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0328b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06516] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0328c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06518] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0328d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0651a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0328e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0651c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0328f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0651e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03290] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06520] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03291] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06522] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03292] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06524] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03293] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06526] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03294] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06528] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03295] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0652a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03296] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0652c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03297] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0652e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03298] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06530] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03299] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06532] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0329a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06534] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0329b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06536] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0329c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06538] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0329d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0653a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0329e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0653c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0329f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0653e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06540] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06542] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06544] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06546] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06548] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0654a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0654c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0654e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06550] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06552] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06554] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06556] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06558] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0655a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0655c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0655e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06560] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06562] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06564] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06566] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06568] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0656a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0656c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0656e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06570] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06572] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06574] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06576] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06578] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0657a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0657c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0657e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06580] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06582] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06584] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06586] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06588] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0658a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0658c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0658e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06590] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06592] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06594] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06596] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06598] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0659a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0659c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0659e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h032ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h065fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03300] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06600] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03301] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06602] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03302] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06604] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03303] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06606] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03304] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06608] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03305] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0660a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03306] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0660c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03307] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0660e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03308] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06610] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03309] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06612] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0330a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06614] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0330b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06616] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0330c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06618] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0330d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0661a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0330e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0661c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0330f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0661e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03310] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06620] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03311] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06622] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03312] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06624] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03313] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06626] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03314] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06628] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03315] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0662a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03316] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0662c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03317] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0662e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03318] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06630] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03319] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06632] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0331a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06634] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0331b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06636] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0331c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06638] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0331d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0663a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0331e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0663c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0331f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0663e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03320] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06640] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03321] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06642] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03322] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06644] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03323] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06646] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03324] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06648] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03325] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0664a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03326] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0664c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03327] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0664e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03328] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06650] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03329] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06652] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0332a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06654] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0332b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06656] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0332c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06658] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0332d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0665a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0332e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0665c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0332f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0665e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03330] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06660] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03331] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06662] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03332] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06664] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03333] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06666] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03334] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06668] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03335] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0666a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03336] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0666c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03337] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0666e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03338] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06670] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03339] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06672] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0333a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06674] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0333b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06676] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0333c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06678] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0333d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0667a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0333e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0667c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0333f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0667e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03340] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06680] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03341] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06682] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03342] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06684] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03343] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06686] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03344] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06688] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03345] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0668a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03346] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0668c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03347] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0668e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03348] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06690] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03349] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06692] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0334a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06694] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0334b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06696] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0334c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06698] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0334d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0669a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0334e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0669c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0334f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0669e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03350] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03351] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03352] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03353] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03354] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03355] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03356] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03357] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03358] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03359] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0335a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0335b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0335c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0335d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0335e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0335f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03360] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03361] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03362] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03363] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03364] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03365] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03366] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03367] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03368] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03369] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0336a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0336b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0336c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0336d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0336e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0336f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03370] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03371] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03372] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03373] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03374] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03375] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03376] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03377] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03378] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03379] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0337a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0337b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0337c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0337d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0337e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0337f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h066fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03380] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06700] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03381] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06702] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03382] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06704] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03383] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06706] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03384] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06708] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03385] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0670a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03386] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0670c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03387] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0670e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03388] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06710] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03389] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06712] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0338a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06714] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0338b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06716] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0338c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06718] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0338d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0671a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0338e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0671c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0338f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0671e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03390] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06720] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03391] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06722] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03392] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06724] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03393] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06726] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03394] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06728] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03395] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0672a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03396] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0672c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03397] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0672e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03398] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06730] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03399] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06732] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0339a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06734] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0339b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06736] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0339c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06738] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0339d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0673a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0339e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0673c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0339f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0673e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06740] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06742] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06744] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06746] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06748] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0674a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0674c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0674e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06750] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06752] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06754] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06756] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06758] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0675a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0675c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0675e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06760] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06762] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06764] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06766] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06768] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0676a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0676c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0676e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06770] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06772] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06774] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06776] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06778] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0677a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0677c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0677e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06780] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06782] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06784] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06786] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06788] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0678a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0678c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0678e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06790] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06792] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06794] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06796] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06798] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0679a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0679c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0679e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h033ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h067fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03400] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06800] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03401] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06802] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03402] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06804] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03403] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06806] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03404] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06808] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03405] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0680a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03406] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0680c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03407] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0680e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03408] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06810] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03409] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06812] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0340a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06814] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0340b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06816] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0340c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06818] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0340d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0681a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0340e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0681c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0340f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0681e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03410] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06820] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03411] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06822] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03412] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06824] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03413] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06826] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03414] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06828] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03415] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0682a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03416] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0682c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03417] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0682e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03418] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06830] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03419] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06832] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0341a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06834] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0341b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06836] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0341c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06838] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0341d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0683a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0341e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0683c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0341f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0683e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03420] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06840] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03421] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06842] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03422] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06844] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03423] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06846] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03424] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06848] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03425] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0684a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03426] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0684c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03427] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0684e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03428] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06850] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03429] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06852] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0342a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06854] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0342b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06856] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0342c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06858] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0342d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0685a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0342e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0685c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0342f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0685e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03430] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06860] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03431] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06862] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03432] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06864] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03433] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06866] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03434] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06868] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03435] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0686a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03436] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0686c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03437] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0686e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03438] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06870] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03439] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06872] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0343a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06874] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0343b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06876] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0343c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06878] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0343d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0687a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0343e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0687c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0343f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0687e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03440] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06880] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03441] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06882] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03442] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06884] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03443] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06886] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03444] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06888] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03445] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0688a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03446] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0688c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03447] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0688e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03448] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06890] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03449] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06892] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0344a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06894] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0344b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06896] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0344c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06898] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0344d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0689a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0344e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0689c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0344f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0689e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03450] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03451] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03452] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03453] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03454] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03455] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03456] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03457] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03458] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03459] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0345a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0345b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0345c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0345d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0345e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0345f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03460] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03461] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03462] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03463] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03464] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03465] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03466] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03467] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03468] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03469] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0346a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0346b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0346c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0346d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0346e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0346f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03470] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03471] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03472] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03473] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03474] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03475] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03476] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03477] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03478] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03479] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0347a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0347b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0347c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0347d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0347e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0347f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h068fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03480] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06900] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03481] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06902] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03482] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06904] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03483] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06906] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03484] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06908] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03485] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0690a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03486] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0690c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03487] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0690e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03488] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06910] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03489] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06912] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0348a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06914] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0348b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06916] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0348c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06918] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0348d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0691a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0348e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0691c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0348f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0691e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03490] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06920] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03491] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06922] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03492] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06924] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03493] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06926] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03494] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06928] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03495] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0692a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03496] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0692c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03497] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0692e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03498] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06930] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03499] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06932] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0349a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06934] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0349b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06936] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0349c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06938] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0349d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0693a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0349e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0693c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0349f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0693e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06940] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06942] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06944] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06946] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06948] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0694a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0694c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0694e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06950] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06952] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06954] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06956] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06958] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0695a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0695c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0695e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06960] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06962] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06964] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06966] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06968] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0696a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0696c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0696e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06970] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06972] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06974] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06976] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06978] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0697a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0697c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0697e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06980] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06982] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06984] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06986] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06988] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0698a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0698c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0698e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06990] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06992] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06994] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06996] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06998] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0699a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0699c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0699e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h034ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h069fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03500] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03501] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03502] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03503] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03504] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03505] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03506] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03507] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03508] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03509] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0350a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0350b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0350c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0350d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0350e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0350f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03510] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03511] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03512] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03513] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03514] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03515] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03516] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03517] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03518] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03519] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0351a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0351b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0351c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0351d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0351e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0351f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03520] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03521] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03522] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03523] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03524] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03525] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03526] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03527] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03528] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03529] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0352a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0352b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0352c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0352d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0352e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0352f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03530] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03531] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03532] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03533] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03534] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03535] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03536] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03537] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03538] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03539] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0353a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0353b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0353c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0353d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0353e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0353f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03540] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03541] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03542] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03543] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03544] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03545] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03546] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03547] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03548] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03549] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0354a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0354b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0354c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0354d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0354e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0354f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06a9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03550] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03551] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03552] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03553] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03554] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03555] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03556] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03557] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03558] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ab0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03559] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ab2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0355a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ab4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0355b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ab6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0355c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ab8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0355d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0355e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06abc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0355f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06abe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03560] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ac0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03561] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ac2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03562] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ac4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03563] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ac6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03564] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ac8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03565] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03566] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06acc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03567] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ace] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03568] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ad0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03569] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ad2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0356a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ad4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0356b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ad6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0356c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ad8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0356d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ada] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0356e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06adc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0356f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ade] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03570] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ae0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03571] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ae2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03572] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ae4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03573] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ae6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03574] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ae8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03575] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03576] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03577] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06aee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03578] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06af0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03579] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06af2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0357a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06af4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0357b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06af6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0357c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06af8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0357d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06afa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0357e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06afc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0357f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06afe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03580] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03581] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03582] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03583] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03584] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03585] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03586] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03587] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03588] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03589] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0358a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0358b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0358c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0358d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0358e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0358f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03590] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03591] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03592] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03593] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03594] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03595] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03596] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03597] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03598] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03599] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0359a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0359b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0359c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0359d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0359e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0359f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06b9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ba0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ba2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ba4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ba6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ba8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06baa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06be0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06be2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06be4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06be6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06be8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h035ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06bfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03600] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03601] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03602] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03603] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03604] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03605] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03606] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03607] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03608] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03609] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0360a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0360b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0360c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0360d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0360e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0360f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03610] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03611] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03612] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03613] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03614] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03615] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03616] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03617] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03618] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03619] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0361a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0361b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0361c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0361d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0361e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0361f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03620] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03621] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03622] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03623] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03624] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03625] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03626] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03627] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03628] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03629] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0362a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0362b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0362c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0362d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0362e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0362f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03630] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03631] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03632] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03633] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03634] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03635] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03636] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03637] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03638] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03639] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0363a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0363b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0363c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0363d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0363e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0363f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03640] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03641] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03642] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03643] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03644] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03645] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03646] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03647] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03648] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03649] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0364a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0364b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0364c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0364d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0364e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0364f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06c9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03650] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ca0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03651] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ca2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03652] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ca4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03653] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ca6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03654] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ca8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03655] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06caa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03656] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03657] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03658] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03659] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0365a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0365b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0365c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0365d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0365e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0365f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03660] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03661] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03662] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03663] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03664] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03665] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03666] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ccc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03667] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03668] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03669] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0366a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0366b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0366c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0366d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0366e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0366f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03670] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ce0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03671] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ce2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03672] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ce4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03673] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ce6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03674] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ce8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03675] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03676] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03677] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03678] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03679] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0367a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0367b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0367c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0367d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0367e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0367f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06cfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03680] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03681] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03682] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03683] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03684] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03685] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03686] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03687] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03688] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03689] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0368a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0368b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0368c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0368d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0368e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0368f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03690] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03691] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03692] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03693] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03694] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03695] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03696] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03697] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03698] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03699] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0369a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0369b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0369c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0369d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0369e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0369f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06d9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06da0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06da2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06da4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06da6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06da8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06daa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06db0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06db2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06db4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06db6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06db8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ddc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06de0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06de2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06de4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06de6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06de8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06df0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06df2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06df4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06df6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06df8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h036ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06dfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03700] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03701] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03702] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03703] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03704] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03705] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03706] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03707] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03708] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03709] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0370a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0370b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0370c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0370d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0370e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0370f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03710] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03711] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03712] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03713] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03714] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03715] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03716] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03717] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03718] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03719] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0371a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0371b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0371c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0371d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0371e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0371f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03720] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03721] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03722] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03723] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03724] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03725] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03726] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03727] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03728] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03729] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0372a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0372b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0372c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0372d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0372e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0372f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03730] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03731] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03732] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03733] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03734] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03735] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03736] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03737] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03738] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03739] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0373a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0373b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0373c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0373d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0373e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0373f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03740] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03741] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03742] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03743] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03744] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03745] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03746] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03747] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03748] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03749] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0374a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0374b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0374c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0374d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0374e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0374f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06e9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03750] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ea0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03751] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ea2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03752] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ea4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03753] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ea6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03754] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ea8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03755] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03756] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03757] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03758] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03759] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0375a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0375b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0375c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0375d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0375e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ebc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0375f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ebe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03760] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ec0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03761] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ec2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03762] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ec4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03763] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ec6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03764] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ec8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03765] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03766] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ecc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03767] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ece] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03768] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ed0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03769] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ed2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0376a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ed4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0376b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ed6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0376c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ed8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0376d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0376e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06edc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0376f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ede] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03770] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ee0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03771] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ee2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03772] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ee4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03773] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ee6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03774] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ee8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03775] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03776] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03777] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06eee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03778] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ef0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03779] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ef2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0377a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ef4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0377b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ef6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0377c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ef8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0377d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06efa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0377e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06efc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0377f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06efe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03780] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03781] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03782] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03783] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03784] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03785] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03786] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03787] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03788] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03789] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0378a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0378b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0378c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0378d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0378e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0378f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03790] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03791] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03792] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03793] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03794] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03795] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03796] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03797] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03798] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03799] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0379a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0379b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0379c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0379d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0379e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0379f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06f9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06faa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fe0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fe2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fe4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fe6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fe8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06fee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ff0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ff2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ff4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ff6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ff8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ffa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ffc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h037ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h06ffe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03800] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07000] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03801] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07002] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03802] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07004] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03803] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07006] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03804] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07008] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03805] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0700a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03806] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0700c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03807] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0700e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03808] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07010] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03809] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07012] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0380a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07014] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0380b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07016] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0380c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07018] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0380d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0701a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0380e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0701c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0380f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0701e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03810] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07020] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03811] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07022] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03812] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07024] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03813] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07026] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03814] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07028] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03815] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0702a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03816] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0702c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03817] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0702e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03818] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07030] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03819] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07032] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0381a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07034] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0381b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07036] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0381c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07038] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0381d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0703a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0381e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0703c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0381f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0703e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03820] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07040] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03821] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07042] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03822] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07044] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03823] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07046] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03824] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07048] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03825] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0704a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03826] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0704c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03827] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0704e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03828] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07050] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03829] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07052] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0382a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07054] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0382b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07056] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0382c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07058] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0382d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0705a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0382e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0705c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0382f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0705e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03830] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07060] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03831] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07062] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03832] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07064] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03833] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07066] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03834] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07068] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03835] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0706a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03836] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0706c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03837] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0706e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03838] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07070] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03839] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07072] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0383a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07074] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0383b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07076] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0383c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07078] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0383d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0707a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0383e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0707c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0383f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0707e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03840] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07080] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03841] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07082] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03842] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07084] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03843] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07086] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03844] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07088] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03845] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0708a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03846] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0708c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03847] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0708e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03848] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07090] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03849] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07092] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0384a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07094] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0384b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07096] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0384c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07098] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0384d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0709a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0384e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0709c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0384f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0709e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03850] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03851] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03852] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03853] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03854] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03855] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03856] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03857] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03858] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03859] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0385a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0385b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0385c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0385d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0385e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0385f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03860] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03861] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03862] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03863] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03864] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03865] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03866] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03867] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03868] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03869] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0386a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0386b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0386c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0386d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0386e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0386f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03870] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03871] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03872] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03873] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03874] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03875] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03876] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03877] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03878] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03879] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0387a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0387b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0387c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0387d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0387e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0387f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h070fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03880] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07100] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03881] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07102] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03882] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07104] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03883] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07106] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03884] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07108] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03885] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0710a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03886] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0710c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03887] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0710e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03888] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07110] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03889] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07112] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0388a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07114] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0388b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07116] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0388c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07118] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0388d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0711a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0388e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0711c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0388f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0711e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03890] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07120] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03891] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07122] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03892] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07124] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03893] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07126] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03894] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07128] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03895] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0712a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03896] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0712c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03897] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0712e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03898] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07130] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03899] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07132] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0389a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07134] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0389b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07136] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0389c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07138] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0389d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0713a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0389e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0713c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0389f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0713e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07140] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07142] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07144] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07146] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07148] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0714a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0714c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0714e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07150] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07152] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07154] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07156] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07158] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0715a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0715c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0715e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07160] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07162] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07164] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07166] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07168] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0716a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0716c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0716e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07170] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07172] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07174] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07176] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07178] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0717a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0717c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0717e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07180] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07182] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07184] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07186] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07188] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0718a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0718c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0718e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07190] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07192] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07194] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07196] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07198] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0719a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0719c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0719e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h038ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h071fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03900] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07200] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03901] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07202] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03902] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07204] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03903] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07206] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03904] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07208] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03905] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0720a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03906] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0720c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03907] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0720e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03908] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07210] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03909] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07212] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0390a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07214] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0390b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07216] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0390c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07218] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0390d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0721a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0390e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0721c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0390f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0721e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03910] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07220] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03911] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07222] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03912] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07224] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03913] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07226] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03914] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07228] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03915] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0722a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03916] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0722c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03917] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0722e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03918] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07230] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03919] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07232] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0391a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07234] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0391b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07236] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0391c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07238] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0391d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0723a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0391e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0723c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0391f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0723e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03920] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07240] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03921] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07242] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03922] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07244] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03923] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07246] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03924] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07248] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03925] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0724a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03926] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0724c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03927] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0724e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03928] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07250] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03929] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07252] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0392a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07254] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0392b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07256] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0392c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07258] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0392d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0725a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0392e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0725c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0392f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0725e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03930] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07260] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03931] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07262] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03932] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07264] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03933] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07266] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03934] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07268] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03935] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0726a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03936] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0726c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03937] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0726e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03938] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07270] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03939] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07272] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0393a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07274] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0393b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07276] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0393c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07278] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0393d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0727a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0393e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0727c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0393f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0727e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03940] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07280] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03941] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07282] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03942] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07284] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03943] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07286] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03944] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07288] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03945] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0728a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03946] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0728c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03947] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0728e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03948] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07290] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03949] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07292] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0394a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07294] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0394b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07296] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0394c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07298] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0394d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0729a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0394e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0729c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0394f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0729e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03950] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03951] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03952] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03953] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03954] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03955] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03956] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03957] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03958] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03959] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0395a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0395b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0395c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0395d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0395e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0395f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03960] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03961] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03962] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03963] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03964] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03965] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03966] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03967] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03968] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03969] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0396a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0396b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0396c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0396d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0396e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0396f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03970] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03971] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03972] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03973] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03974] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03975] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03976] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03977] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03978] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03979] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0397a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0397b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0397c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0397d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0397e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0397f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h072fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03980] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07300] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03981] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07302] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03982] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07304] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03983] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07306] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03984] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07308] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03985] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0730a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03986] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0730c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03987] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0730e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03988] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07310] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03989] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07312] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0398a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07314] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0398b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07316] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0398c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07318] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0398d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0731a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0398e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0731c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0398f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0731e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03990] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07320] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03991] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07322] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03992] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07324] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03993] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07326] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03994] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07328] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03995] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0732a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03996] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0732c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03997] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0732e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03998] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07330] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03999] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07332] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0399a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07334] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0399b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07336] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0399c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07338] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0399d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0733a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0399e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0733c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h0399f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0733e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039a0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07340] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039a1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07342] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039a2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07344] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039a3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07346] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039a4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07348] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039a5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0734a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039a6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0734c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039a7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0734e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039a8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07350] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039a9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07352] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039aa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07354] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07356] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07358] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0735a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0735c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039af] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0735e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039b0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07360] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039b1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07362] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039b2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07364] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039b3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07366] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039b4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07368] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039b5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0736a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039b6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0736c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039b7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0736e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039b8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07370] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039b9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07372] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07374] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039bb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07376] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039bc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07378] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039bd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0737a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039be] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0737c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039bf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0737e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039c0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07380] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039c1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07382] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039c2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07384] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039c3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07386] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039c4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07388] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039c5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0738a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039c6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0738c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039c7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0738e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039c8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07390] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039c9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07392] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07394] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039cb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07396] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039cc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07398] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039cd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0739a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0739c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039cf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0739e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039d0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039d1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039d2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039d3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039d4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039d5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039d6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039d7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039d8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039d9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039da] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039db] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039dc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039dd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039de] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039df] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039e0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039e1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039e2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039e3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039e4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039e5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039e6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039e7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039e8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039e9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039eb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039f0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039f1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039f2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039f3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039f4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039f5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039f6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039f7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039f8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039f9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039fa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039fb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039fc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039fd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039fe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h039ff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h073fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07400] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07402] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07404] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07406] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07408] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0740a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0740c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0740e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07410] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07412] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07414] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07416] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07418] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0741a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0741c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0741e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07420] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07422] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07424] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07426] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07428] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0742a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0742c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0742e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07430] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07432] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07434] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07436] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07438] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0743a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0743c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0743e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07440] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07442] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07444] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07446] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07448] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0744a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0744c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0744e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07450] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07452] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07454] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07456] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07458] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0745a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0745c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0745e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07460] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07462] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07464] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07466] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07468] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0746a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0746c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0746e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07470] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07472] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07474] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07476] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07478] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0747a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0747c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0747e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07480] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07482] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07484] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07486] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07488] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0748a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0748c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0748e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07490] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07492] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07494] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07496] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07498] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0749a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0749c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0749e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h074fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07500] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07502] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07504] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07506] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07508] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0750a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0750c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0750e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07510] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07512] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07514] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07516] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07518] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0751a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0751c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0751e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07520] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07522] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07524] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07526] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07528] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0752a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0752c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0752e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07530] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07532] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07534] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07536] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07538] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0753a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0753c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03a9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0753e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aa0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07540] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aa1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07542] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aa2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07544] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aa3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07546] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aa4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07548] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aa5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0754a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aa6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0754c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aa7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0754e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aa8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07550] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aa9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07552] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aaa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07554] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07556] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07558] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0755a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0755c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aaf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0755e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ab0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07560] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ab1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07562] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ab2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07564] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ab3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07566] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ab4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07568] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ab5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0756a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ab6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0756c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ab7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0756e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ab8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07570] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ab9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07572] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07574] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03abb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07576] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03abc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07578] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03abd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0757a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03abe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0757c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03abf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0757e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ac0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07580] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ac1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07582] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ac2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07584] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ac3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07586] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ac4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07588] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ac5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0758a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ac6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0758c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ac7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0758e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ac8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07590] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ac9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07592] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07594] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03acb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07596] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03acc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07598] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03acd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0759a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ace] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0759c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03acf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0759e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ad0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ad1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ad2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ad3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ad4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ad5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ad6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ad7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ad8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ad9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ada] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03adb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03adc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03add] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ade] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03adf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ae0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ae1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ae2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ae3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ae4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ae5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ae6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ae7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ae8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ae9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aeb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03af0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03af1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03af2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03af3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03af4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03af5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03af6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03af7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03af8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03af9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03afa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03afb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03afc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03afd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03afe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03aff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h075fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07600] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07602] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07604] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07606] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07608] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0760a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0760c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0760e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07610] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07612] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07614] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07616] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07618] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0761a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0761c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0761e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07620] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07622] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07624] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07626] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07628] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0762a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0762c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0762e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07630] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07632] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07634] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07636] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07638] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0763a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0763c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0763e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07640] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07642] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07644] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07646] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07648] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0764a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0764c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0764e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07650] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07652] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07654] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07656] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07658] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0765a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0765c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0765e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07660] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07662] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07664] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07666] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07668] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0766a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0766c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0766e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07670] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07672] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07674] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07676] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07678] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0767a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0767c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0767e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07680] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07682] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07684] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07686] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07688] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0768a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0768c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0768e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07690] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07692] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07694] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07696] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07698] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0769a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0769c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0769e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h076fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07700] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07702] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07704] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07706] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07708] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0770a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0770c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0770e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07710] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07712] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07714] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07716] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07718] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0771a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0771c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0771e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07720] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07722] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07724] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07726] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07728] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0772a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0772c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0772e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07730] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07732] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07734] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07736] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07738] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0773a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0773c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03b9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0773e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ba0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07740] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ba1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07742] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ba2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07744] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ba3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07746] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ba4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07748] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ba5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0774a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ba6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0774c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ba7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0774e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ba8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07750] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ba9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07752] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03baa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07754] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07756] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07758] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0775a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0775c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03baf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0775e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07760] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07762] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07764] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07766] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07768] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0776a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0776c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0776e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07770] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07772] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07774] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07776] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07778] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0777a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0777c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0777e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07780] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07782] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07784] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07786] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07788] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0778a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0778c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0778e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07790] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07792] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07794] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07796] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07798] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0779a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0779c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0779e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03be0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03be1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03be2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03be3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03be4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03be5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03be6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03be7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03be8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03be9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03beb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bf0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bf1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bf2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bf3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bf4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bf5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bf6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bf7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bf8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bf9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03bff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h077fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07800] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07802] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07804] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07806] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07808] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0780a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0780c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0780e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07810] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07812] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07814] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07816] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07818] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0781a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0781c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0781e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07820] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07822] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07824] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07826] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07828] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0782a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0782c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0782e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07830] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07832] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07834] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07836] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07838] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0783a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0783c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0783e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07840] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07842] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07844] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07846] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07848] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0784a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0784c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0784e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07850] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07852] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07854] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07856] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07858] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0785a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0785c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0785e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07860] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07862] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07864] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07866] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07868] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0786a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0786c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0786e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07870] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07872] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07874] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07876] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07878] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0787a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0787c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0787e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07880] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07882] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07884] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07886] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07888] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0788a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0788c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0788e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07890] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07892] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07894] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07896] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07898] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0789a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0789c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0789e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h078fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07900] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07902] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07904] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07906] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07908] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0790a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0790c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0790e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07910] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07912] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07914] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07916] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07918] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0791a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0791c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0791e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07920] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07922] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07924] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07926] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07928] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0792a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0792c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0792e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07930] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07932] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07934] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07936] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07938] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0793a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0793c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03c9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0793e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ca0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07940] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ca1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07942] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ca2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07944] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ca3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07946] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ca4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07948] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ca5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0794a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ca6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0794c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ca7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0794e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ca8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07950] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ca9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07952] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03caa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07954] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07956] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07958] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0795a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0795c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03caf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0795e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07960] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07962] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07964] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07966] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07968] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0796a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0796c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0796e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07970] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07972] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07974] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07976] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07978] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0797a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0797c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0797e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07980] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07982] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07984] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07986] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07988] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0798a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0798c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0798e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07990] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07992] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07994] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ccb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07996] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ccc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07998] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ccd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0799a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0799c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ccf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h0799e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079a0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079a2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079a4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079a6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079a8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079aa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079ac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079ae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079b0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079b2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079b4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079b6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079b8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079ba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079bc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079be] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ce0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079c0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ce1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079c2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ce2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079c4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ce3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079c6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ce4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079c8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ce5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079ca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ce6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079cc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ce7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079ce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ce8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079d0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ce9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079d2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079d4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ceb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079d6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079d8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ced] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079da] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079dc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079de] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cf0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079e0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cf1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079e2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cf2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079e4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cf3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079e6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cf4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079e8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cf5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079ea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cf6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079ec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cf7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079ee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cf8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079f0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cf9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079f2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079f4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079f6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079f8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079fa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079fc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03cff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h079fe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07a9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ab0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ab2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ab4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ab6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ab8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07abc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07abe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ac0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ac2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ac4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ac6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ac8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07acc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ace] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ad0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ad2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ad4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ad6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ad8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ada] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07adc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ade] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ae0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ae2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ae4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ae6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ae8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07aee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07af0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07af2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07af4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07af6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07af8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07afa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07afc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07afe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03d9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03da0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03da1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03da2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03da3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03da4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03da5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03da6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03da7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03da8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03da9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03daa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03daf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03db0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03db1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03db2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03db3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03db4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03db5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03db6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03db7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03db8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03db9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07b9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ba0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ba2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ba4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ba6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ba8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07baa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ddb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ddc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ddd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ddf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03de0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03de1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03de2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03de3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03de4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03de5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03de6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03de7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03de8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03de9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03deb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ded] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03def] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03df0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07be0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03df1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07be2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03df2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07be4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03df3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07be6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03df4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07be8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03df5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03df6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03df7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03df8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03df9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dfa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dfb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dfc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dfd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dfe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03dff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07bfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07c9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ca0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ca2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ca4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ca6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ca8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07caa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ccc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ce0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ce2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ce4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ce6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ce8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cf0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cf2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cf4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cf6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cf8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07cfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03e9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ea0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ea1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ea2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ea3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ea4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ea5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ea6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ea7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ea8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ea9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eaa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ead] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eaf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ebb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ebc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ebd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ebe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ebf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ec0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ec1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ec2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ec3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ec4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ec5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ec6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ec7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ec8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ec9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ecb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ecc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ecd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ece] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ecf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07d9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ed0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07da0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ed1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07da2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ed2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07da4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ed3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07da6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ed4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07da8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ed5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07daa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ed6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ed7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ed8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07db0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ed9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07db2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07db4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03edb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07db6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03edc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07db8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03edd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ede] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03edf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ee0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ee1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ee2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ee3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ee4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ee5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ee6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ee7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ee8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ee9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eeb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ddc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ef0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07de0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ef1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07de2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ef2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07de4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ef3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07de6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ef4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07de8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ef5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ef6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ef7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ef8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07df0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ef9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07df2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03efa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07df4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03efb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07df6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03efc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07df8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03efd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dfa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03efe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dfc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03eff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07dfe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f00] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f01] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f02] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f03] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f04] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f05] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f06] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f07] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f08] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f09] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f0a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f0b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f0c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f0d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f0e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f0f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f10] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f11] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f12] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f13] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f14] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f15] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f16] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f17] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f18] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f19] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f1a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f1b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f1c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f1d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f1e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f1f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f20] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f21] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f22] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f23] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f24] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f25] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f26] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f27] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f28] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f29] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f2a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f2b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f2c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f2d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f2e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f2f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f30] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f31] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f32] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f33] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f34] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f35] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f36] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f37] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f38] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f39] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f3a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f3b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f3c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f3d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f3e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f3f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f40] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f41] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f42] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f43] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f44] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f45] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f46] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f47] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f48] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f49] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f4a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f4b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f4c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f4d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f4e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f4f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07e9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f50] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ea0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f51] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ea2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f52] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ea4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f53] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ea6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f54] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ea8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f55] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eaa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f56] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f57] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f58] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f59] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f5a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f5b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f5c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f5d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f5e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ebc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f5f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ebe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f60] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ec0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f61] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ec2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f62] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ec4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f63] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ec6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f64] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ec8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f65] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f66] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ecc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f67] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ece] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f68] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ed0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f69] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ed2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f6a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ed4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f6b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ed6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f6c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ed8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f6d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f6e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07edc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f6f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ede] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f70] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ee0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f71] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ee2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f72] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ee4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f73] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ee6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f74] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ee8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f75] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f76] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f77] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07eee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f78] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ef0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f79] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ef2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f7a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ef4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f7b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ef6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f7c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ef8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f7d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07efa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f7e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07efc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f7f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07efe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f80] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f00] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f81] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f02] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f82] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f04] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f83] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f06] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f84] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f08] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f85] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f0a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f86] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f0c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f87] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f0e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f88] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f10] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f89] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f12] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f8a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f14] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f8b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f16] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f8c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f18] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f8d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f1a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f8e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f1c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f8f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f1e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f90] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f20] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f91] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f22] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f92] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f24] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f93] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f26] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f94] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f28] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f95] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f2a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f96] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f2c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f97] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f2e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f98] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f30] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f99] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f32] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f9a] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f34] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f9b] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f36] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f9c] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f38] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f9d] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f3a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f9e] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f3c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03f9f] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f3e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fa0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f40] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fa1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f42] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fa2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f44] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fa3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f46] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fa4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f48] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fa5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f4a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fa6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f4c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fa7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f4e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fa8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f50] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fa9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f52] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03faa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f54] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fab] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f56] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fac] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f58] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fad] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f5a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fae] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f5c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03faf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f5e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fb0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f60] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fb1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f62] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fb2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f64] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fb3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f66] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fb4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f68] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fb5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f6a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fb6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f6c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fb7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f6e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fb8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f70] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fb9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f72] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fba] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f74] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fbb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f76] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fbc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f78] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fbd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f7a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fbe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f7c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fbf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f7e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fc0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f80] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fc1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f82] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fc2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f84] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fc3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f86] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fc4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f88] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fc5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f8a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fc6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f8c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fc7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f8e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fc8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f90] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fc9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f92] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fca] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f94] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fcb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f96] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fcc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f98] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fcd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f9a] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fce] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f9c] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fcf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07f9e] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fd0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fa0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fd1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fa2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fd2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fa4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fd3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fa6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fd4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fa8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fd5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07faa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fd6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fac] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fd7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fae] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fd8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fb0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fd9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fb2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fda] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fb4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fdb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fb6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fdc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fb8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fdd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fba] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fde] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fbc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fdf] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fbe] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fe0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fc0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fe1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fc2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fe2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fc4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fe3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fc6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fe4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fc8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fe5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fca] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fe6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fcc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fe7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fce] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fe8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fd0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fe9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fd2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fea] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fd4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03feb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fd6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fec] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fd8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fed] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fda] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fee] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fdc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fef] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fde] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ff0] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fe0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ff1] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fe2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ff2] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fe4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ff3] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fe6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ff4] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fe8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ff5] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fea] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ff6] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fec] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ff7] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07fee] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ff8] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ff0] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ff9] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ff2] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ffa] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ff4] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ffb] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ff6] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ffc] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ff8] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ffd] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ffa] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03ffe] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ffc] ;
//end
//always_comb begin // 
               Ifd35529b44c957737bf422127283c08e['h03fff] =  I6eb3a3e04397efbe48cc2f5809bfcb98['h07ffe] ;
//end
