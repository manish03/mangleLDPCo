//`include "GF2_LDPC_fgallag_0x00006_assign_inc.sv"
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00000] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00000] : //%
                       If409768b648a33a7ed878a070d4f6251['h00001] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00001] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00002] : //%
                       If409768b648a33a7ed878a070d4f6251['h00003] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00002] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00004] : //%
                       If409768b648a33a7ed878a070d4f6251['h00005] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00003] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00006] : //%
                       If409768b648a33a7ed878a070d4f6251['h00007] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00004] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00008] : //%
                       If409768b648a33a7ed878a070d4f6251['h00009] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00005] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0000a] : //%
                       If409768b648a33a7ed878a070d4f6251['h0000b] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00006] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0000c] : //%
                       If409768b648a33a7ed878a070d4f6251['h0000d] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00007] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0000e] : //%
                       If409768b648a33a7ed878a070d4f6251['h0000f] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00008] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00010] : //%
                       If409768b648a33a7ed878a070d4f6251['h00011] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00009] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00012] : //%
                       If409768b648a33a7ed878a070d4f6251['h00013] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0000a] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00014] : //%
                       If409768b648a33a7ed878a070d4f6251['h00015] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0000b] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00016] : //%
                       If409768b648a33a7ed878a070d4f6251['h00017] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0000c] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00018] : //%
                       If409768b648a33a7ed878a070d4f6251['h00019] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0000d] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0001a] : //%
                       If409768b648a33a7ed878a070d4f6251['h0001b] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0000e] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0001c] : //%
                       If409768b648a33a7ed878a070d4f6251['h0001d] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0000f] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0001e] : //%
                       If409768b648a33a7ed878a070d4f6251['h0001f] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00010] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00020] : //%
                       If409768b648a33a7ed878a070d4f6251['h00021] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00011] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00022] : //%
                       If409768b648a33a7ed878a070d4f6251['h00023] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00012] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00024] : //%
                       If409768b648a33a7ed878a070d4f6251['h00025] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00013] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00026] : //%
                       If409768b648a33a7ed878a070d4f6251['h00027] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00014] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00028] : //%
                       If409768b648a33a7ed878a070d4f6251['h00029] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00015] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0002a] : //%
                       If409768b648a33a7ed878a070d4f6251['h0002b] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00016] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0002c] : //%
                       If409768b648a33a7ed878a070d4f6251['h0002d] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00017] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0002e] : //%
                       If409768b648a33a7ed878a070d4f6251['h0002f] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00018] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00030] : //%
                       If409768b648a33a7ed878a070d4f6251['h00031] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00019] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00032] : //%
                       If409768b648a33a7ed878a070d4f6251['h00033] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0001a] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00034] : //%
                       If409768b648a33a7ed878a070d4f6251['h00035] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0001b] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00036] : //%
                       If409768b648a33a7ed878a070d4f6251['h00037] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0001c] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00038] : //%
                       If409768b648a33a7ed878a070d4f6251['h00039] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0001d] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0003a] : //%
                       If409768b648a33a7ed878a070d4f6251['h0003b] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0001e] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0003c] : //%
                       If409768b648a33a7ed878a070d4f6251['h0003d] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0001f] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0003e] : //%
                       If409768b648a33a7ed878a070d4f6251['h0003f] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00020] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00040] : //%
                       If409768b648a33a7ed878a070d4f6251['h00041] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00021] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00042] : //%
                       If409768b648a33a7ed878a070d4f6251['h00043] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00022] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00044] : //%
                       If409768b648a33a7ed878a070d4f6251['h00045] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00023] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00046] : //%
                       If409768b648a33a7ed878a070d4f6251['h00047] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00024] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00048] : //%
                       If409768b648a33a7ed878a070d4f6251['h00049] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00025] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0004a] : //%
                       If409768b648a33a7ed878a070d4f6251['h0004b] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00026] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0004c] : //%
                       If409768b648a33a7ed878a070d4f6251['h0004d] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00027] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0004e] : //%
                       If409768b648a33a7ed878a070d4f6251['h0004f] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00028] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00050] : //%
                       If409768b648a33a7ed878a070d4f6251['h00051] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00029] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00052] : //%
                       If409768b648a33a7ed878a070d4f6251['h00053] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0002a] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00054] : //%
                       If409768b648a33a7ed878a070d4f6251['h00055] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0002b] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00056] : //%
                       If409768b648a33a7ed878a070d4f6251['h00057] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0002c] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00058] : //%
                       If409768b648a33a7ed878a070d4f6251['h00059] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0002d] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0005a] : //%
                       If409768b648a33a7ed878a070d4f6251['h0005b] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0002e] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0005c] : //%
                       If409768b648a33a7ed878a070d4f6251['h0005d] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0002f] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0005e] : //%
                       If409768b648a33a7ed878a070d4f6251['h0005f] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00030] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00060] : //%
                       If409768b648a33a7ed878a070d4f6251['h00061] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00031] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00062] : //%
                       If409768b648a33a7ed878a070d4f6251['h00063] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00032] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00064] : //%
                       If409768b648a33a7ed878a070d4f6251['h00065] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00033] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00066] : //%
                       If409768b648a33a7ed878a070d4f6251['h00067] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00034] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00068] : //%
                       If409768b648a33a7ed878a070d4f6251['h00069] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00035] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0006a] : //%
                       If409768b648a33a7ed878a070d4f6251['h0006b] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00036] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0006c] : //%
                       If409768b648a33a7ed878a070d4f6251['h0006d] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00037] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0006e] : //%
                       If409768b648a33a7ed878a070d4f6251['h0006f] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00038] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00070] : //%
                       If409768b648a33a7ed878a070d4f6251['h00071] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00039] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00072] : //%
                       If409768b648a33a7ed878a070d4f6251['h00073] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0003a] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00074] : //%
                       If409768b648a33a7ed878a070d4f6251['h00075] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0003b] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00076] : //%
                       If409768b648a33a7ed878a070d4f6251['h00077] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0003c] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00078] : //%
                       If409768b648a33a7ed878a070d4f6251['h00079] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0003d] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0007a] : //%
                       If409768b648a33a7ed878a070d4f6251['h0007b] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0003e] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0007c] : //%
                       If409768b648a33a7ed878a070d4f6251['h0007d] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0003f] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0007e] : //%
                       If409768b648a33a7ed878a070d4f6251['h0007f] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00040] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00080] : //%
                       If409768b648a33a7ed878a070d4f6251['h00081] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00041] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00082] : //%
                       If409768b648a33a7ed878a070d4f6251['h00083] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00042] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00084] : //%
                       If409768b648a33a7ed878a070d4f6251['h00085] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00043] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00086] : //%
                       If409768b648a33a7ed878a070d4f6251['h00087] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00044] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00088] : //%
                       If409768b648a33a7ed878a070d4f6251['h00089] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00045] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0008a] : //%
                       If409768b648a33a7ed878a070d4f6251['h0008b] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00046] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0008c] : //%
                       If409768b648a33a7ed878a070d4f6251['h0008d] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00047] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0008e] : //%
                       If409768b648a33a7ed878a070d4f6251['h0008f] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00048] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00090] : //%
                       If409768b648a33a7ed878a070d4f6251['h00091] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00049] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00092] : //%
                       If409768b648a33a7ed878a070d4f6251['h00093] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0004a] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00094] : //%
                       If409768b648a33a7ed878a070d4f6251['h00095] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0004b] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00096] : //%
                       If409768b648a33a7ed878a070d4f6251['h00097] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0004c] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00098] : //%
                       If409768b648a33a7ed878a070d4f6251['h00099] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0004d] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0009a] : //%
                       If409768b648a33a7ed878a070d4f6251['h0009b] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0004e] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0009c] : //%
                       If409768b648a33a7ed878a070d4f6251['h0009d] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0004f] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h0009e] : //%
                       If409768b648a33a7ed878a070d4f6251['h0009f] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00050] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000a0] : //%
                       If409768b648a33a7ed878a070d4f6251['h000a1] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00051] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000a2] : //%
                       If409768b648a33a7ed878a070d4f6251['h000a3] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00052] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000a4] : //%
                       If409768b648a33a7ed878a070d4f6251['h000a5] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00053] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000a6] : //%
                       If409768b648a33a7ed878a070d4f6251['h000a7] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00054] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000a8] : //%
                       If409768b648a33a7ed878a070d4f6251['h000a9] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00055] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000aa] : //%
                       If409768b648a33a7ed878a070d4f6251['h000ab] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00056] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000ac] : //%
                       If409768b648a33a7ed878a070d4f6251['h000ad] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00057] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000ae] : //%
                       If409768b648a33a7ed878a070d4f6251['h000af] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00058] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000b0] : //%
                       If409768b648a33a7ed878a070d4f6251['h000b1] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00059] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000b2] : //%
                       If409768b648a33a7ed878a070d4f6251['h000b3] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0005a] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000b4] : //%
                       If409768b648a33a7ed878a070d4f6251['h000b5] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0005b] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000b6] : //%
                       If409768b648a33a7ed878a070d4f6251['h000b7] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0005c] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000b8] : //%
                       If409768b648a33a7ed878a070d4f6251['h000b9] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0005d] =  If409768b648a33a7ed878a070d4f6251['h000ba] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0005e] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000bc] : //%
                       If409768b648a33a7ed878a070d4f6251['h000bd] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0005f] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000be] : //%
                       If409768b648a33a7ed878a070d4f6251['h000bf] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00060] =  If409768b648a33a7ed878a070d4f6251['h000c0] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00061] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000c2] : //%
                       If409768b648a33a7ed878a070d4f6251['h000c3] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00062] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000c4] : //%
                       If409768b648a33a7ed878a070d4f6251['h000c5] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00063] =  If409768b648a33a7ed878a070d4f6251['h000c6] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00064] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000c8] : //%
                       If409768b648a33a7ed878a070d4f6251['h000c9] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00065] =  If409768b648a33a7ed878a070d4f6251['h000ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00066] =  If409768b648a33a7ed878a070d4f6251['h000cc] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00067] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000ce] : //%
                       If409768b648a33a7ed878a070d4f6251['h000cf] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00068] =  If409768b648a33a7ed878a070d4f6251['h000d0] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00069] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000d2] : //%
                       If409768b648a33a7ed878a070d4f6251['h000d3] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0006a] =  If409768b648a33a7ed878a070d4f6251['h000d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0006b] =  If409768b648a33a7ed878a070d4f6251['h000d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0006c] =  If409768b648a33a7ed878a070d4f6251['h000d8] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0006d] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000da] : //%
                       If409768b648a33a7ed878a070d4f6251['h000db] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0006e] =  If409768b648a33a7ed878a070d4f6251['h000dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0006f] =  If409768b648a33a7ed878a070d4f6251['h000de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00070] =  If409768b648a33a7ed878a070d4f6251['h000e0] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00071] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000e2] : //%
                       If409768b648a33a7ed878a070d4f6251['h000e3] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00072] =  If409768b648a33a7ed878a070d4f6251['h000e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00073] =  If409768b648a33a7ed878a070d4f6251['h000e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00074] =  If409768b648a33a7ed878a070d4f6251['h000e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00075] =  If409768b648a33a7ed878a070d4f6251['h000ea] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00076] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000ec] : //%
                       If409768b648a33a7ed878a070d4f6251['h000ed] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00077] =  If409768b648a33a7ed878a070d4f6251['h000ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00078] =  If409768b648a33a7ed878a070d4f6251['h000f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00079] =  If409768b648a33a7ed878a070d4f6251['h000f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0007a] =  If409768b648a33a7ed878a070d4f6251['h000f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0007b] =  If409768b648a33a7ed878a070d4f6251['h000f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0007c] =  If409768b648a33a7ed878a070d4f6251['h000f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0007d] =  If409768b648a33a7ed878a070d4f6251['h000fa] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h0007e] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h000fc] : //%
                       If409768b648a33a7ed878a070d4f6251['h000fd] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0007f] =  If409768b648a33a7ed878a070d4f6251['h000fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00080] =  If409768b648a33a7ed878a070d4f6251['h00100] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00081] =  If409768b648a33a7ed878a070d4f6251['h00102] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00082] =  If409768b648a33a7ed878a070d4f6251['h00104] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00083] =  If409768b648a33a7ed878a070d4f6251['h00106] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00084] =  If409768b648a33a7ed878a070d4f6251['h00108] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00085] =  If409768b648a33a7ed878a070d4f6251['h0010a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00086] =  If409768b648a33a7ed878a070d4f6251['h0010c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00087] =  If409768b648a33a7ed878a070d4f6251['h0010e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00088] =  If409768b648a33a7ed878a070d4f6251['h00110] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00089] =  If409768b648a33a7ed878a070d4f6251['h00112] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0008a] =  If409768b648a33a7ed878a070d4f6251['h00114] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0008b] =  If409768b648a33a7ed878a070d4f6251['h00116] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0008c] =  If409768b648a33a7ed878a070d4f6251['h00118] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0008d] =  If409768b648a33a7ed878a070d4f6251['h0011a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0008e] =  If409768b648a33a7ed878a070d4f6251['h0011c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0008f] =  If409768b648a33a7ed878a070d4f6251['h0011e] ;
//end
//always_comb begin
              Ic8a4ab93493bd6cdd4939054e46d2247['h00090] = 
          (!fgallag_sel['h00006]) ? 
                       If409768b648a33a7ed878a070d4f6251['h00120] : //%
                       If409768b648a33a7ed878a070d4f6251['h00121] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00091] =  If409768b648a33a7ed878a070d4f6251['h00122] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00092] =  If409768b648a33a7ed878a070d4f6251['h00124] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00093] =  If409768b648a33a7ed878a070d4f6251['h00126] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00094] =  If409768b648a33a7ed878a070d4f6251['h00128] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00095] =  If409768b648a33a7ed878a070d4f6251['h0012a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00096] =  If409768b648a33a7ed878a070d4f6251['h0012c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00097] =  If409768b648a33a7ed878a070d4f6251['h0012e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00098] =  If409768b648a33a7ed878a070d4f6251['h00130] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00099] =  If409768b648a33a7ed878a070d4f6251['h00132] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0009a] =  If409768b648a33a7ed878a070d4f6251['h00134] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0009b] =  If409768b648a33a7ed878a070d4f6251['h00136] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0009c] =  If409768b648a33a7ed878a070d4f6251['h00138] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0009d] =  If409768b648a33a7ed878a070d4f6251['h0013a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0009e] =  If409768b648a33a7ed878a070d4f6251['h0013c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0009f] =  If409768b648a33a7ed878a070d4f6251['h0013e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000a0] =  If409768b648a33a7ed878a070d4f6251['h00140] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000a1] =  If409768b648a33a7ed878a070d4f6251['h00142] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000a2] =  If409768b648a33a7ed878a070d4f6251['h00144] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000a3] =  If409768b648a33a7ed878a070d4f6251['h00146] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000a4] =  If409768b648a33a7ed878a070d4f6251['h00148] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000a5] =  If409768b648a33a7ed878a070d4f6251['h0014a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000a6] =  If409768b648a33a7ed878a070d4f6251['h0014c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000a7] =  If409768b648a33a7ed878a070d4f6251['h0014e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000a8] =  If409768b648a33a7ed878a070d4f6251['h00150] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000a9] =  If409768b648a33a7ed878a070d4f6251['h00152] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000aa] =  If409768b648a33a7ed878a070d4f6251['h00154] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ab] =  If409768b648a33a7ed878a070d4f6251['h00156] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ac] =  If409768b648a33a7ed878a070d4f6251['h00158] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ad] =  If409768b648a33a7ed878a070d4f6251['h0015a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ae] =  If409768b648a33a7ed878a070d4f6251['h0015c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000af] =  If409768b648a33a7ed878a070d4f6251['h0015e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000b0] =  If409768b648a33a7ed878a070d4f6251['h00160] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000b1] =  If409768b648a33a7ed878a070d4f6251['h00162] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000b2] =  If409768b648a33a7ed878a070d4f6251['h00164] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000b3] =  If409768b648a33a7ed878a070d4f6251['h00166] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000b4] =  If409768b648a33a7ed878a070d4f6251['h00168] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000b5] =  If409768b648a33a7ed878a070d4f6251['h0016a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000b6] =  If409768b648a33a7ed878a070d4f6251['h0016c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000b7] =  If409768b648a33a7ed878a070d4f6251['h0016e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000b8] =  If409768b648a33a7ed878a070d4f6251['h00170] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000b9] =  If409768b648a33a7ed878a070d4f6251['h00172] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ba] =  If409768b648a33a7ed878a070d4f6251['h00174] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000bb] =  If409768b648a33a7ed878a070d4f6251['h00176] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000bc] =  If409768b648a33a7ed878a070d4f6251['h00178] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000bd] =  If409768b648a33a7ed878a070d4f6251['h0017a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000be] =  If409768b648a33a7ed878a070d4f6251['h0017c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000bf] =  If409768b648a33a7ed878a070d4f6251['h0017e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000c0] =  If409768b648a33a7ed878a070d4f6251['h00180] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000c1] =  If409768b648a33a7ed878a070d4f6251['h00182] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000c2] =  If409768b648a33a7ed878a070d4f6251['h00184] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000c3] =  If409768b648a33a7ed878a070d4f6251['h00186] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000c4] =  If409768b648a33a7ed878a070d4f6251['h00188] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000c5] =  If409768b648a33a7ed878a070d4f6251['h0018a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000c6] =  If409768b648a33a7ed878a070d4f6251['h0018c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000c7] =  If409768b648a33a7ed878a070d4f6251['h0018e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000c8] =  If409768b648a33a7ed878a070d4f6251['h00190] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000c9] =  If409768b648a33a7ed878a070d4f6251['h00192] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ca] =  If409768b648a33a7ed878a070d4f6251['h00194] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000cb] =  If409768b648a33a7ed878a070d4f6251['h00196] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000cc] =  If409768b648a33a7ed878a070d4f6251['h00198] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000cd] =  If409768b648a33a7ed878a070d4f6251['h0019a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ce] =  If409768b648a33a7ed878a070d4f6251['h0019c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000cf] =  If409768b648a33a7ed878a070d4f6251['h0019e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000d0] =  If409768b648a33a7ed878a070d4f6251['h001a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000d1] =  If409768b648a33a7ed878a070d4f6251['h001a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000d2] =  If409768b648a33a7ed878a070d4f6251['h001a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000d3] =  If409768b648a33a7ed878a070d4f6251['h001a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000d4] =  If409768b648a33a7ed878a070d4f6251['h001a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000d5] =  If409768b648a33a7ed878a070d4f6251['h001aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000d6] =  If409768b648a33a7ed878a070d4f6251['h001ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000d7] =  If409768b648a33a7ed878a070d4f6251['h001ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000d8] =  If409768b648a33a7ed878a070d4f6251['h001b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000d9] =  If409768b648a33a7ed878a070d4f6251['h001b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000da] =  If409768b648a33a7ed878a070d4f6251['h001b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000db] =  If409768b648a33a7ed878a070d4f6251['h001b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000dc] =  If409768b648a33a7ed878a070d4f6251['h001b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000dd] =  If409768b648a33a7ed878a070d4f6251['h001ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000de] =  If409768b648a33a7ed878a070d4f6251['h001bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000df] =  If409768b648a33a7ed878a070d4f6251['h001be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000e0] =  If409768b648a33a7ed878a070d4f6251['h001c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000e1] =  If409768b648a33a7ed878a070d4f6251['h001c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000e2] =  If409768b648a33a7ed878a070d4f6251['h001c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000e3] =  If409768b648a33a7ed878a070d4f6251['h001c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000e4] =  If409768b648a33a7ed878a070d4f6251['h001c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000e5] =  If409768b648a33a7ed878a070d4f6251['h001ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000e6] =  If409768b648a33a7ed878a070d4f6251['h001cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000e7] =  If409768b648a33a7ed878a070d4f6251['h001ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000e8] =  If409768b648a33a7ed878a070d4f6251['h001d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000e9] =  If409768b648a33a7ed878a070d4f6251['h001d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ea] =  If409768b648a33a7ed878a070d4f6251['h001d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000eb] =  If409768b648a33a7ed878a070d4f6251['h001d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ec] =  If409768b648a33a7ed878a070d4f6251['h001d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ed] =  If409768b648a33a7ed878a070d4f6251['h001da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ee] =  If409768b648a33a7ed878a070d4f6251['h001dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ef] =  If409768b648a33a7ed878a070d4f6251['h001de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000f0] =  If409768b648a33a7ed878a070d4f6251['h001e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000f1] =  If409768b648a33a7ed878a070d4f6251['h001e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000f2] =  If409768b648a33a7ed878a070d4f6251['h001e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000f3] =  If409768b648a33a7ed878a070d4f6251['h001e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000f4] =  If409768b648a33a7ed878a070d4f6251['h001e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000f5] =  If409768b648a33a7ed878a070d4f6251['h001ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000f6] =  If409768b648a33a7ed878a070d4f6251['h001ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000f7] =  If409768b648a33a7ed878a070d4f6251['h001ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000f8] =  If409768b648a33a7ed878a070d4f6251['h001f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000f9] =  If409768b648a33a7ed878a070d4f6251['h001f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000fa] =  If409768b648a33a7ed878a070d4f6251['h001f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000fb] =  If409768b648a33a7ed878a070d4f6251['h001f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000fc] =  If409768b648a33a7ed878a070d4f6251['h001f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000fd] =  If409768b648a33a7ed878a070d4f6251['h001fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000fe] =  If409768b648a33a7ed878a070d4f6251['h001fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h000ff] =  If409768b648a33a7ed878a070d4f6251['h001fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00100] =  If409768b648a33a7ed878a070d4f6251['h00200] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00101] =  If409768b648a33a7ed878a070d4f6251['h00202] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00102] =  If409768b648a33a7ed878a070d4f6251['h00204] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00103] =  If409768b648a33a7ed878a070d4f6251['h00206] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00104] =  If409768b648a33a7ed878a070d4f6251['h00208] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00105] =  If409768b648a33a7ed878a070d4f6251['h0020a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00106] =  If409768b648a33a7ed878a070d4f6251['h0020c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00107] =  If409768b648a33a7ed878a070d4f6251['h0020e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00108] =  If409768b648a33a7ed878a070d4f6251['h00210] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00109] =  If409768b648a33a7ed878a070d4f6251['h00212] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0010a] =  If409768b648a33a7ed878a070d4f6251['h00214] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0010b] =  If409768b648a33a7ed878a070d4f6251['h00216] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0010c] =  If409768b648a33a7ed878a070d4f6251['h00218] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0010d] =  If409768b648a33a7ed878a070d4f6251['h0021a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0010e] =  If409768b648a33a7ed878a070d4f6251['h0021c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0010f] =  If409768b648a33a7ed878a070d4f6251['h0021e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00110] =  If409768b648a33a7ed878a070d4f6251['h00220] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00111] =  If409768b648a33a7ed878a070d4f6251['h00222] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00112] =  If409768b648a33a7ed878a070d4f6251['h00224] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00113] =  If409768b648a33a7ed878a070d4f6251['h00226] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00114] =  If409768b648a33a7ed878a070d4f6251['h00228] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00115] =  If409768b648a33a7ed878a070d4f6251['h0022a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00116] =  If409768b648a33a7ed878a070d4f6251['h0022c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00117] =  If409768b648a33a7ed878a070d4f6251['h0022e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00118] =  If409768b648a33a7ed878a070d4f6251['h00230] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00119] =  If409768b648a33a7ed878a070d4f6251['h00232] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0011a] =  If409768b648a33a7ed878a070d4f6251['h00234] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0011b] =  If409768b648a33a7ed878a070d4f6251['h00236] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0011c] =  If409768b648a33a7ed878a070d4f6251['h00238] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0011d] =  If409768b648a33a7ed878a070d4f6251['h0023a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0011e] =  If409768b648a33a7ed878a070d4f6251['h0023c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0011f] =  If409768b648a33a7ed878a070d4f6251['h0023e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00120] =  If409768b648a33a7ed878a070d4f6251['h00240] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00121] =  If409768b648a33a7ed878a070d4f6251['h00242] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00122] =  If409768b648a33a7ed878a070d4f6251['h00244] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00123] =  If409768b648a33a7ed878a070d4f6251['h00246] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00124] =  If409768b648a33a7ed878a070d4f6251['h00248] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00125] =  If409768b648a33a7ed878a070d4f6251['h0024a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00126] =  If409768b648a33a7ed878a070d4f6251['h0024c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00127] =  If409768b648a33a7ed878a070d4f6251['h0024e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00128] =  If409768b648a33a7ed878a070d4f6251['h00250] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00129] =  If409768b648a33a7ed878a070d4f6251['h00252] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0012a] =  If409768b648a33a7ed878a070d4f6251['h00254] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0012b] =  If409768b648a33a7ed878a070d4f6251['h00256] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0012c] =  If409768b648a33a7ed878a070d4f6251['h00258] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0012d] =  If409768b648a33a7ed878a070d4f6251['h0025a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0012e] =  If409768b648a33a7ed878a070d4f6251['h0025c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0012f] =  If409768b648a33a7ed878a070d4f6251['h0025e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00130] =  If409768b648a33a7ed878a070d4f6251['h00260] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00131] =  If409768b648a33a7ed878a070d4f6251['h00262] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00132] =  If409768b648a33a7ed878a070d4f6251['h00264] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00133] =  If409768b648a33a7ed878a070d4f6251['h00266] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00134] =  If409768b648a33a7ed878a070d4f6251['h00268] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00135] =  If409768b648a33a7ed878a070d4f6251['h0026a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00136] =  If409768b648a33a7ed878a070d4f6251['h0026c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00137] =  If409768b648a33a7ed878a070d4f6251['h0026e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00138] =  If409768b648a33a7ed878a070d4f6251['h00270] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00139] =  If409768b648a33a7ed878a070d4f6251['h00272] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0013a] =  If409768b648a33a7ed878a070d4f6251['h00274] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0013b] =  If409768b648a33a7ed878a070d4f6251['h00276] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0013c] =  If409768b648a33a7ed878a070d4f6251['h00278] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0013d] =  If409768b648a33a7ed878a070d4f6251['h0027a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0013e] =  If409768b648a33a7ed878a070d4f6251['h0027c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0013f] =  If409768b648a33a7ed878a070d4f6251['h0027e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00140] =  If409768b648a33a7ed878a070d4f6251['h00280] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00141] =  If409768b648a33a7ed878a070d4f6251['h00282] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00142] =  If409768b648a33a7ed878a070d4f6251['h00284] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00143] =  If409768b648a33a7ed878a070d4f6251['h00286] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00144] =  If409768b648a33a7ed878a070d4f6251['h00288] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00145] =  If409768b648a33a7ed878a070d4f6251['h0028a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00146] =  If409768b648a33a7ed878a070d4f6251['h0028c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00147] =  If409768b648a33a7ed878a070d4f6251['h0028e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00148] =  If409768b648a33a7ed878a070d4f6251['h00290] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00149] =  If409768b648a33a7ed878a070d4f6251['h00292] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0014a] =  If409768b648a33a7ed878a070d4f6251['h00294] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0014b] =  If409768b648a33a7ed878a070d4f6251['h00296] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0014c] =  If409768b648a33a7ed878a070d4f6251['h00298] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0014d] =  If409768b648a33a7ed878a070d4f6251['h0029a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0014e] =  If409768b648a33a7ed878a070d4f6251['h0029c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0014f] =  If409768b648a33a7ed878a070d4f6251['h0029e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00150] =  If409768b648a33a7ed878a070d4f6251['h002a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00151] =  If409768b648a33a7ed878a070d4f6251['h002a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00152] =  If409768b648a33a7ed878a070d4f6251['h002a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00153] =  If409768b648a33a7ed878a070d4f6251['h002a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00154] =  If409768b648a33a7ed878a070d4f6251['h002a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00155] =  If409768b648a33a7ed878a070d4f6251['h002aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00156] =  If409768b648a33a7ed878a070d4f6251['h002ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00157] =  If409768b648a33a7ed878a070d4f6251['h002ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00158] =  If409768b648a33a7ed878a070d4f6251['h002b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00159] =  If409768b648a33a7ed878a070d4f6251['h002b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0015a] =  If409768b648a33a7ed878a070d4f6251['h002b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0015b] =  If409768b648a33a7ed878a070d4f6251['h002b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0015c] =  If409768b648a33a7ed878a070d4f6251['h002b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0015d] =  If409768b648a33a7ed878a070d4f6251['h002ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0015e] =  If409768b648a33a7ed878a070d4f6251['h002bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0015f] =  If409768b648a33a7ed878a070d4f6251['h002be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00160] =  If409768b648a33a7ed878a070d4f6251['h002c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00161] =  If409768b648a33a7ed878a070d4f6251['h002c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00162] =  If409768b648a33a7ed878a070d4f6251['h002c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00163] =  If409768b648a33a7ed878a070d4f6251['h002c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00164] =  If409768b648a33a7ed878a070d4f6251['h002c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00165] =  If409768b648a33a7ed878a070d4f6251['h002ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00166] =  If409768b648a33a7ed878a070d4f6251['h002cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00167] =  If409768b648a33a7ed878a070d4f6251['h002ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00168] =  If409768b648a33a7ed878a070d4f6251['h002d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00169] =  If409768b648a33a7ed878a070d4f6251['h002d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0016a] =  If409768b648a33a7ed878a070d4f6251['h002d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0016b] =  If409768b648a33a7ed878a070d4f6251['h002d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0016c] =  If409768b648a33a7ed878a070d4f6251['h002d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0016d] =  If409768b648a33a7ed878a070d4f6251['h002da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0016e] =  If409768b648a33a7ed878a070d4f6251['h002dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0016f] =  If409768b648a33a7ed878a070d4f6251['h002de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00170] =  If409768b648a33a7ed878a070d4f6251['h002e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00171] =  If409768b648a33a7ed878a070d4f6251['h002e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00172] =  If409768b648a33a7ed878a070d4f6251['h002e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00173] =  If409768b648a33a7ed878a070d4f6251['h002e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00174] =  If409768b648a33a7ed878a070d4f6251['h002e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00175] =  If409768b648a33a7ed878a070d4f6251['h002ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00176] =  If409768b648a33a7ed878a070d4f6251['h002ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00177] =  If409768b648a33a7ed878a070d4f6251['h002ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00178] =  If409768b648a33a7ed878a070d4f6251['h002f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00179] =  If409768b648a33a7ed878a070d4f6251['h002f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0017a] =  If409768b648a33a7ed878a070d4f6251['h002f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0017b] =  If409768b648a33a7ed878a070d4f6251['h002f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0017c] =  If409768b648a33a7ed878a070d4f6251['h002f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0017d] =  If409768b648a33a7ed878a070d4f6251['h002fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0017e] =  If409768b648a33a7ed878a070d4f6251['h002fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0017f] =  If409768b648a33a7ed878a070d4f6251['h002fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00180] =  If409768b648a33a7ed878a070d4f6251['h00300] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00181] =  If409768b648a33a7ed878a070d4f6251['h00302] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00182] =  If409768b648a33a7ed878a070d4f6251['h00304] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00183] =  If409768b648a33a7ed878a070d4f6251['h00306] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00184] =  If409768b648a33a7ed878a070d4f6251['h00308] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00185] =  If409768b648a33a7ed878a070d4f6251['h0030a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00186] =  If409768b648a33a7ed878a070d4f6251['h0030c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00187] =  If409768b648a33a7ed878a070d4f6251['h0030e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00188] =  If409768b648a33a7ed878a070d4f6251['h00310] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00189] =  If409768b648a33a7ed878a070d4f6251['h00312] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0018a] =  If409768b648a33a7ed878a070d4f6251['h00314] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0018b] =  If409768b648a33a7ed878a070d4f6251['h00316] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0018c] =  If409768b648a33a7ed878a070d4f6251['h00318] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0018d] =  If409768b648a33a7ed878a070d4f6251['h0031a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0018e] =  If409768b648a33a7ed878a070d4f6251['h0031c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0018f] =  If409768b648a33a7ed878a070d4f6251['h0031e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00190] =  If409768b648a33a7ed878a070d4f6251['h00320] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00191] =  If409768b648a33a7ed878a070d4f6251['h00322] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00192] =  If409768b648a33a7ed878a070d4f6251['h00324] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00193] =  If409768b648a33a7ed878a070d4f6251['h00326] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00194] =  If409768b648a33a7ed878a070d4f6251['h00328] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00195] =  If409768b648a33a7ed878a070d4f6251['h0032a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00196] =  If409768b648a33a7ed878a070d4f6251['h0032c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00197] =  If409768b648a33a7ed878a070d4f6251['h0032e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00198] =  If409768b648a33a7ed878a070d4f6251['h00330] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00199] =  If409768b648a33a7ed878a070d4f6251['h00332] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0019a] =  If409768b648a33a7ed878a070d4f6251['h00334] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0019b] =  If409768b648a33a7ed878a070d4f6251['h00336] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0019c] =  If409768b648a33a7ed878a070d4f6251['h00338] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0019d] =  If409768b648a33a7ed878a070d4f6251['h0033a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0019e] =  If409768b648a33a7ed878a070d4f6251['h0033c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0019f] =  If409768b648a33a7ed878a070d4f6251['h0033e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001a0] =  If409768b648a33a7ed878a070d4f6251['h00340] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001a1] =  If409768b648a33a7ed878a070d4f6251['h00342] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001a2] =  If409768b648a33a7ed878a070d4f6251['h00344] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001a3] =  If409768b648a33a7ed878a070d4f6251['h00346] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001a4] =  If409768b648a33a7ed878a070d4f6251['h00348] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001a5] =  If409768b648a33a7ed878a070d4f6251['h0034a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001a6] =  If409768b648a33a7ed878a070d4f6251['h0034c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001a7] =  If409768b648a33a7ed878a070d4f6251['h0034e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001a8] =  If409768b648a33a7ed878a070d4f6251['h00350] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001a9] =  If409768b648a33a7ed878a070d4f6251['h00352] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001aa] =  If409768b648a33a7ed878a070d4f6251['h00354] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ab] =  If409768b648a33a7ed878a070d4f6251['h00356] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ac] =  If409768b648a33a7ed878a070d4f6251['h00358] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ad] =  If409768b648a33a7ed878a070d4f6251['h0035a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ae] =  If409768b648a33a7ed878a070d4f6251['h0035c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001af] =  If409768b648a33a7ed878a070d4f6251['h0035e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001b0] =  If409768b648a33a7ed878a070d4f6251['h00360] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001b1] =  If409768b648a33a7ed878a070d4f6251['h00362] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001b2] =  If409768b648a33a7ed878a070d4f6251['h00364] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001b3] =  If409768b648a33a7ed878a070d4f6251['h00366] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001b4] =  If409768b648a33a7ed878a070d4f6251['h00368] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001b5] =  If409768b648a33a7ed878a070d4f6251['h0036a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001b6] =  If409768b648a33a7ed878a070d4f6251['h0036c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001b7] =  If409768b648a33a7ed878a070d4f6251['h0036e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001b8] =  If409768b648a33a7ed878a070d4f6251['h00370] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001b9] =  If409768b648a33a7ed878a070d4f6251['h00372] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ba] =  If409768b648a33a7ed878a070d4f6251['h00374] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001bb] =  If409768b648a33a7ed878a070d4f6251['h00376] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001bc] =  If409768b648a33a7ed878a070d4f6251['h00378] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001bd] =  If409768b648a33a7ed878a070d4f6251['h0037a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001be] =  If409768b648a33a7ed878a070d4f6251['h0037c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001bf] =  If409768b648a33a7ed878a070d4f6251['h0037e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001c0] =  If409768b648a33a7ed878a070d4f6251['h00380] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001c1] =  If409768b648a33a7ed878a070d4f6251['h00382] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001c2] =  If409768b648a33a7ed878a070d4f6251['h00384] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001c3] =  If409768b648a33a7ed878a070d4f6251['h00386] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001c4] =  If409768b648a33a7ed878a070d4f6251['h00388] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001c5] =  If409768b648a33a7ed878a070d4f6251['h0038a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001c6] =  If409768b648a33a7ed878a070d4f6251['h0038c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001c7] =  If409768b648a33a7ed878a070d4f6251['h0038e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001c8] =  If409768b648a33a7ed878a070d4f6251['h00390] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001c9] =  If409768b648a33a7ed878a070d4f6251['h00392] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ca] =  If409768b648a33a7ed878a070d4f6251['h00394] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001cb] =  If409768b648a33a7ed878a070d4f6251['h00396] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001cc] =  If409768b648a33a7ed878a070d4f6251['h00398] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001cd] =  If409768b648a33a7ed878a070d4f6251['h0039a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ce] =  If409768b648a33a7ed878a070d4f6251['h0039c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001cf] =  If409768b648a33a7ed878a070d4f6251['h0039e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001d0] =  If409768b648a33a7ed878a070d4f6251['h003a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001d1] =  If409768b648a33a7ed878a070d4f6251['h003a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001d2] =  If409768b648a33a7ed878a070d4f6251['h003a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001d3] =  If409768b648a33a7ed878a070d4f6251['h003a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001d4] =  If409768b648a33a7ed878a070d4f6251['h003a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001d5] =  If409768b648a33a7ed878a070d4f6251['h003aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001d6] =  If409768b648a33a7ed878a070d4f6251['h003ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001d7] =  If409768b648a33a7ed878a070d4f6251['h003ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001d8] =  If409768b648a33a7ed878a070d4f6251['h003b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001d9] =  If409768b648a33a7ed878a070d4f6251['h003b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001da] =  If409768b648a33a7ed878a070d4f6251['h003b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001db] =  If409768b648a33a7ed878a070d4f6251['h003b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001dc] =  If409768b648a33a7ed878a070d4f6251['h003b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001dd] =  If409768b648a33a7ed878a070d4f6251['h003ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001de] =  If409768b648a33a7ed878a070d4f6251['h003bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001df] =  If409768b648a33a7ed878a070d4f6251['h003be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001e0] =  If409768b648a33a7ed878a070d4f6251['h003c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001e1] =  If409768b648a33a7ed878a070d4f6251['h003c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001e2] =  If409768b648a33a7ed878a070d4f6251['h003c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001e3] =  If409768b648a33a7ed878a070d4f6251['h003c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001e4] =  If409768b648a33a7ed878a070d4f6251['h003c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001e5] =  If409768b648a33a7ed878a070d4f6251['h003ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001e6] =  If409768b648a33a7ed878a070d4f6251['h003cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001e7] =  If409768b648a33a7ed878a070d4f6251['h003ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001e8] =  If409768b648a33a7ed878a070d4f6251['h003d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001e9] =  If409768b648a33a7ed878a070d4f6251['h003d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ea] =  If409768b648a33a7ed878a070d4f6251['h003d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001eb] =  If409768b648a33a7ed878a070d4f6251['h003d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ec] =  If409768b648a33a7ed878a070d4f6251['h003d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ed] =  If409768b648a33a7ed878a070d4f6251['h003da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ee] =  If409768b648a33a7ed878a070d4f6251['h003dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ef] =  If409768b648a33a7ed878a070d4f6251['h003de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001f0] =  If409768b648a33a7ed878a070d4f6251['h003e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001f1] =  If409768b648a33a7ed878a070d4f6251['h003e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001f2] =  If409768b648a33a7ed878a070d4f6251['h003e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001f3] =  If409768b648a33a7ed878a070d4f6251['h003e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001f4] =  If409768b648a33a7ed878a070d4f6251['h003e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001f5] =  If409768b648a33a7ed878a070d4f6251['h003ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001f6] =  If409768b648a33a7ed878a070d4f6251['h003ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001f7] =  If409768b648a33a7ed878a070d4f6251['h003ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001f8] =  If409768b648a33a7ed878a070d4f6251['h003f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001f9] =  If409768b648a33a7ed878a070d4f6251['h003f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001fa] =  If409768b648a33a7ed878a070d4f6251['h003f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001fb] =  If409768b648a33a7ed878a070d4f6251['h003f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001fc] =  If409768b648a33a7ed878a070d4f6251['h003f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001fd] =  If409768b648a33a7ed878a070d4f6251['h003fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001fe] =  If409768b648a33a7ed878a070d4f6251['h003fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h001ff] =  If409768b648a33a7ed878a070d4f6251['h003fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00200] =  If409768b648a33a7ed878a070d4f6251['h00400] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00201] =  If409768b648a33a7ed878a070d4f6251['h00402] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00202] =  If409768b648a33a7ed878a070d4f6251['h00404] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00203] =  If409768b648a33a7ed878a070d4f6251['h00406] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00204] =  If409768b648a33a7ed878a070d4f6251['h00408] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00205] =  If409768b648a33a7ed878a070d4f6251['h0040a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00206] =  If409768b648a33a7ed878a070d4f6251['h0040c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00207] =  If409768b648a33a7ed878a070d4f6251['h0040e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00208] =  If409768b648a33a7ed878a070d4f6251['h00410] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00209] =  If409768b648a33a7ed878a070d4f6251['h00412] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0020a] =  If409768b648a33a7ed878a070d4f6251['h00414] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0020b] =  If409768b648a33a7ed878a070d4f6251['h00416] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0020c] =  If409768b648a33a7ed878a070d4f6251['h00418] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0020d] =  If409768b648a33a7ed878a070d4f6251['h0041a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0020e] =  If409768b648a33a7ed878a070d4f6251['h0041c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0020f] =  If409768b648a33a7ed878a070d4f6251['h0041e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00210] =  If409768b648a33a7ed878a070d4f6251['h00420] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00211] =  If409768b648a33a7ed878a070d4f6251['h00422] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00212] =  If409768b648a33a7ed878a070d4f6251['h00424] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00213] =  If409768b648a33a7ed878a070d4f6251['h00426] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00214] =  If409768b648a33a7ed878a070d4f6251['h00428] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00215] =  If409768b648a33a7ed878a070d4f6251['h0042a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00216] =  If409768b648a33a7ed878a070d4f6251['h0042c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00217] =  If409768b648a33a7ed878a070d4f6251['h0042e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00218] =  If409768b648a33a7ed878a070d4f6251['h00430] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00219] =  If409768b648a33a7ed878a070d4f6251['h00432] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0021a] =  If409768b648a33a7ed878a070d4f6251['h00434] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0021b] =  If409768b648a33a7ed878a070d4f6251['h00436] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0021c] =  If409768b648a33a7ed878a070d4f6251['h00438] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0021d] =  If409768b648a33a7ed878a070d4f6251['h0043a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0021e] =  If409768b648a33a7ed878a070d4f6251['h0043c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0021f] =  If409768b648a33a7ed878a070d4f6251['h0043e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00220] =  If409768b648a33a7ed878a070d4f6251['h00440] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00221] =  If409768b648a33a7ed878a070d4f6251['h00442] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00222] =  If409768b648a33a7ed878a070d4f6251['h00444] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00223] =  If409768b648a33a7ed878a070d4f6251['h00446] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00224] =  If409768b648a33a7ed878a070d4f6251['h00448] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00225] =  If409768b648a33a7ed878a070d4f6251['h0044a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00226] =  If409768b648a33a7ed878a070d4f6251['h0044c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00227] =  If409768b648a33a7ed878a070d4f6251['h0044e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00228] =  If409768b648a33a7ed878a070d4f6251['h00450] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00229] =  If409768b648a33a7ed878a070d4f6251['h00452] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0022a] =  If409768b648a33a7ed878a070d4f6251['h00454] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0022b] =  If409768b648a33a7ed878a070d4f6251['h00456] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0022c] =  If409768b648a33a7ed878a070d4f6251['h00458] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0022d] =  If409768b648a33a7ed878a070d4f6251['h0045a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0022e] =  If409768b648a33a7ed878a070d4f6251['h0045c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0022f] =  If409768b648a33a7ed878a070d4f6251['h0045e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00230] =  If409768b648a33a7ed878a070d4f6251['h00460] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00231] =  If409768b648a33a7ed878a070d4f6251['h00462] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00232] =  If409768b648a33a7ed878a070d4f6251['h00464] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00233] =  If409768b648a33a7ed878a070d4f6251['h00466] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00234] =  If409768b648a33a7ed878a070d4f6251['h00468] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00235] =  If409768b648a33a7ed878a070d4f6251['h0046a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00236] =  If409768b648a33a7ed878a070d4f6251['h0046c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00237] =  If409768b648a33a7ed878a070d4f6251['h0046e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00238] =  If409768b648a33a7ed878a070d4f6251['h00470] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00239] =  If409768b648a33a7ed878a070d4f6251['h00472] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0023a] =  If409768b648a33a7ed878a070d4f6251['h00474] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0023b] =  If409768b648a33a7ed878a070d4f6251['h00476] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0023c] =  If409768b648a33a7ed878a070d4f6251['h00478] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0023d] =  If409768b648a33a7ed878a070d4f6251['h0047a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0023e] =  If409768b648a33a7ed878a070d4f6251['h0047c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0023f] =  If409768b648a33a7ed878a070d4f6251['h0047e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00240] =  If409768b648a33a7ed878a070d4f6251['h00480] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00241] =  If409768b648a33a7ed878a070d4f6251['h00482] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00242] =  If409768b648a33a7ed878a070d4f6251['h00484] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00243] =  If409768b648a33a7ed878a070d4f6251['h00486] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00244] =  If409768b648a33a7ed878a070d4f6251['h00488] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00245] =  If409768b648a33a7ed878a070d4f6251['h0048a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00246] =  If409768b648a33a7ed878a070d4f6251['h0048c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00247] =  If409768b648a33a7ed878a070d4f6251['h0048e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00248] =  If409768b648a33a7ed878a070d4f6251['h00490] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00249] =  If409768b648a33a7ed878a070d4f6251['h00492] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0024a] =  If409768b648a33a7ed878a070d4f6251['h00494] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0024b] =  If409768b648a33a7ed878a070d4f6251['h00496] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0024c] =  If409768b648a33a7ed878a070d4f6251['h00498] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0024d] =  If409768b648a33a7ed878a070d4f6251['h0049a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0024e] =  If409768b648a33a7ed878a070d4f6251['h0049c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0024f] =  If409768b648a33a7ed878a070d4f6251['h0049e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00250] =  If409768b648a33a7ed878a070d4f6251['h004a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00251] =  If409768b648a33a7ed878a070d4f6251['h004a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00252] =  If409768b648a33a7ed878a070d4f6251['h004a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00253] =  If409768b648a33a7ed878a070d4f6251['h004a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00254] =  If409768b648a33a7ed878a070d4f6251['h004a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00255] =  If409768b648a33a7ed878a070d4f6251['h004aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00256] =  If409768b648a33a7ed878a070d4f6251['h004ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00257] =  If409768b648a33a7ed878a070d4f6251['h004ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00258] =  If409768b648a33a7ed878a070d4f6251['h004b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00259] =  If409768b648a33a7ed878a070d4f6251['h004b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0025a] =  If409768b648a33a7ed878a070d4f6251['h004b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0025b] =  If409768b648a33a7ed878a070d4f6251['h004b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0025c] =  If409768b648a33a7ed878a070d4f6251['h004b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0025d] =  If409768b648a33a7ed878a070d4f6251['h004ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0025e] =  If409768b648a33a7ed878a070d4f6251['h004bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0025f] =  If409768b648a33a7ed878a070d4f6251['h004be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00260] =  If409768b648a33a7ed878a070d4f6251['h004c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00261] =  If409768b648a33a7ed878a070d4f6251['h004c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00262] =  If409768b648a33a7ed878a070d4f6251['h004c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00263] =  If409768b648a33a7ed878a070d4f6251['h004c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00264] =  If409768b648a33a7ed878a070d4f6251['h004c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00265] =  If409768b648a33a7ed878a070d4f6251['h004ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00266] =  If409768b648a33a7ed878a070d4f6251['h004cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00267] =  If409768b648a33a7ed878a070d4f6251['h004ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00268] =  If409768b648a33a7ed878a070d4f6251['h004d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00269] =  If409768b648a33a7ed878a070d4f6251['h004d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0026a] =  If409768b648a33a7ed878a070d4f6251['h004d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0026b] =  If409768b648a33a7ed878a070d4f6251['h004d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0026c] =  If409768b648a33a7ed878a070d4f6251['h004d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0026d] =  If409768b648a33a7ed878a070d4f6251['h004da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0026e] =  If409768b648a33a7ed878a070d4f6251['h004dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0026f] =  If409768b648a33a7ed878a070d4f6251['h004de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00270] =  If409768b648a33a7ed878a070d4f6251['h004e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00271] =  If409768b648a33a7ed878a070d4f6251['h004e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00272] =  If409768b648a33a7ed878a070d4f6251['h004e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00273] =  If409768b648a33a7ed878a070d4f6251['h004e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00274] =  If409768b648a33a7ed878a070d4f6251['h004e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00275] =  If409768b648a33a7ed878a070d4f6251['h004ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00276] =  If409768b648a33a7ed878a070d4f6251['h004ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00277] =  If409768b648a33a7ed878a070d4f6251['h004ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00278] =  If409768b648a33a7ed878a070d4f6251['h004f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00279] =  If409768b648a33a7ed878a070d4f6251['h004f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0027a] =  If409768b648a33a7ed878a070d4f6251['h004f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0027b] =  If409768b648a33a7ed878a070d4f6251['h004f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0027c] =  If409768b648a33a7ed878a070d4f6251['h004f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0027d] =  If409768b648a33a7ed878a070d4f6251['h004fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0027e] =  If409768b648a33a7ed878a070d4f6251['h004fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0027f] =  If409768b648a33a7ed878a070d4f6251['h004fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00280] =  If409768b648a33a7ed878a070d4f6251['h00500] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00281] =  If409768b648a33a7ed878a070d4f6251['h00502] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00282] =  If409768b648a33a7ed878a070d4f6251['h00504] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00283] =  If409768b648a33a7ed878a070d4f6251['h00506] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00284] =  If409768b648a33a7ed878a070d4f6251['h00508] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00285] =  If409768b648a33a7ed878a070d4f6251['h0050a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00286] =  If409768b648a33a7ed878a070d4f6251['h0050c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00287] =  If409768b648a33a7ed878a070d4f6251['h0050e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00288] =  If409768b648a33a7ed878a070d4f6251['h00510] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00289] =  If409768b648a33a7ed878a070d4f6251['h00512] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0028a] =  If409768b648a33a7ed878a070d4f6251['h00514] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0028b] =  If409768b648a33a7ed878a070d4f6251['h00516] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0028c] =  If409768b648a33a7ed878a070d4f6251['h00518] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0028d] =  If409768b648a33a7ed878a070d4f6251['h0051a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0028e] =  If409768b648a33a7ed878a070d4f6251['h0051c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0028f] =  If409768b648a33a7ed878a070d4f6251['h0051e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00290] =  If409768b648a33a7ed878a070d4f6251['h00520] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00291] =  If409768b648a33a7ed878a070d4f6251['h00522] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00292] =  If409768b648a33a7ed878a070d4f6251['h00524] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00293] =  If409768b648a33a7ed878a070d4f6251['h00526] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00294] =  If409768b648a33a7ed878a070d4f6251['h00528] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00295] =  If409768b648a33a7ed878a070d4f6251['h0052a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00296] =  If409768b648a33a7ed878a070d4f6251['h0052c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00297] =  If409768b648a33a7ed878a070d4f6251['h0052e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00298] =  If409768b648a33a7ed878a070d4f6251['h00530] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00299] =  If409768b648a33a7ed878a070d4f6251['h00532] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0029a] =  If409768b648a33a7ed878a070d4f6251['h00534] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0029b] =  If409768b648a33a7ed878a070d4f6251['h00536] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0029c] =  If409768b648a33a7ed878a070d4f6251['h00538] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0029d] =  If409768b648a33a7ed878a070d4f6251['h0053a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0029e] =  If409768b648a33a7ed878a070d4f6251['h0053c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0029f] =  If409768b648a33a7ed878a070d4f6251['h0053e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002a0] =  If409768b648a33a7ed878a070d4f6251['h00540] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002a1] =  If409768b648a33a7ed878a070d4f6251['h00542] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002a2] =  If409768b648a33a7ed878a070d4f6251['h00544] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002a3] =  If409768b648a33a7ed878a070d4f6251['h00546] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002a4] =  If409768b648a33a7ed878a070d4f6251['h00548] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002a5] =  If409768b648a33a7ed878a070d4f6251['h0054a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002a6] =  If409768b648a33a7ed878a070d4f6251['h0054c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002a7] =  If409768b648a33a7ed878a070d4f6251['h0054e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002a8] =  If409768b648a33a7ed878a070d4f6251['h00550] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002a9] =  If409768b648a33a7ed878a070d4f6251['h00552] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002aa] =  If409768b648a33a7ed878a070d4f6251['h00554] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ab] =  If409768b648a33a7ed878a070d4f6251['h00556] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ac] =  If409768b648a33a7ed878a070d4f6251['h00558] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ad] =  If409768b648a33a7ed878a070d4f6251['h0055a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ae] =  If409768b648a33a7ed878a070d4f6251['h0055c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002af] =  If409768b648a33a7ed878a070d4f6251['h0055e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002b0] =  If409768b648a33a7ed878a070d4f6251['h00560] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002b1] =  If409768b648a33a7ed878a070d4f6251['h00562] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002b2] =  If409768b648a33a7ed878a070d4f6251['h00564] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002b3] =  If409768b648a33a7ed878a070d4f6251['h00566] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002b4] =  If409768b648a33a7ed878a070d4f6251['h00568] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002b5] =  If409768b648a33a7ed878a070d4f6251['h0056a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002b6] =  If409768b648a33a7ed878a070d4f6251['h0056c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002b7] =  If409768b648a33a7ed878a070d4f6251['h0056e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002b8] =  If409768b648a33a7ed878a070d4f6251['h00570] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002b9] =  If409768b648a33a7ed878a070d4f6251['h00572] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ba] =  If409768b648a33a7ed878a070d4f6251['h00574] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002bb] =  If409768b648a33a7ed878a070d4f6251['h00576] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002bc] =  If409768b648a33a7ed878a070d4f6251['h00578] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002bd] =  If409768b648a33a7ed878a070d4f6251['h0057a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002be] =  If409768b648a33a7ed878a070d4f6251['h0057c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002bf] =  If409768b648a33a7ed878a070d4f6251['h0057e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002c0] =  If409768b648a33a7ed878a070d4f6251['h00580] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002c1] =  If409768b648a33a7ed878a070d4f6251['h00582] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002c2] =  If409768b648a33a7ed878a070d4f6251['h00584] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002c3] =  If409768b648a33a7ed878a070d4f6251['h00586] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002c4] =  If409768b648a33a7ed878a070d4f6251['h00588] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002c5] =  If409768b648a33a7ed878a070d4f6251['h0058a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002c6] =  If409768b648a33a7ed878a070d4f6251['h0058c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002c7] =  If409768b648a33a7ed878a070d4f6251['h0058e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002c8] =  If409768b648a33a7ed878a070d4f6251['h00590] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002c9] =  If409768b648a33a7ed878a070d4f6251['h00592] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ca] =  If409768b648a33a7ed878a070d4f6251['h00594] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002cb] =  If409768b648a33a7ed878a070d4f6251['h00596] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002cc] =  If409768b648a33a7ed878a070d4f6251['h00598] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002cd] =  If409768b648a33a7ed878a070d4f6251['h0059a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ce] =  If409768b648a33a7ed878a070d4f6251['h0059c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002cf] =  If409768b648a33a7ed878a070d4f6251['h0059e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002d0] =  If409768b648a33a7ed878a070d4f6251['h005a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002d1] =  If409768b648a33a7ed878a070d4f6251['h005a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002d2] =  If409768b648a33a7ed878a070d4f6251['h005a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002d3] =  If409768b648a33a7ed878a070d4f6251['h005a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002d4] =  If409768b648a33a7ed878a070d4f6251['h005a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002d5] =  If409768b648a33a7ed878a070d4f6251['h005aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002d6] =  If409768b648a33a7ed878a070d4f6251['h005ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002d7] =  If409768b648a33a7ed878a070d4f6251['h005ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002d8] =  If409768b648a33a7ed878a070d4f6251['h005b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002d9] =  If409768b648a33a7ed878a070d4f6251['h005b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002da] =  If409768b648a33a7ed878a070d4f6251['h005b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002db] =  If409768b648a33a7ed878a070d4f6251['h005b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002dc] =  If409768b648a33a7ed878a070d4f6251['h005b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002dd] =  If409768b648a33a7ed878a070d4f6251['h005ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002de] =  If409768b648a33a7ed878a070d4f6251['h005bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002df] =  If409768b648a33a7ed878a070d4f6251['h005be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002e0] =  If409768b648a33a7ed878a070d4f6251['h005c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002e1] =  If409768b648a33a7ed878a070d4f6251['h005c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002e2] =  If409768b648a33a7ed878a070d4f6251['h005c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002e3] =  If409768b648a33a7ed878a070d4f6251['h005c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002e4] =  If409768b648a33a7ed878a070d4f6251['h005c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002e5] =  If409768b648a33a7ed878a070d4f6251['h005ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002e6] =  If409768b648a33a7ed878a070d4f6251['h005cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002e7] =  If409768b648a33a7ed878a070d4f6251['h005ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002e8] =  If409768b648a33a7ed878a070d4f6251['h005d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002e9] =  If409768b648a33a7ed878a070d4f6251['h005d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ea] =  If409768b648a33a7ed878a070d4f6251['h005d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002eb] =  If409768b648a33a7ed878a070d4f6251['h005d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ec] =  If409768b648a33a7ed878a070d4f6251['h005d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ed] =  If409768b648a33a7ed878a070d4f6251['h005da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ee] =  If409768b648a33a7ed878a070d4f6251['h005dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ef] =  If409768b648a33a7ed878a070d4f6251['h005de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002f0] =  If409768b648a33a7ed878a070d4f6251['h005e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002f1] =  If409768b648a33a7ed878a070d4f6251['h005e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002f2] =  If409768b648a33a7ed878a070d4f6251['h005e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002f3] =  If409768b648a33a7ed878a070d4f6251['h005e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002f4] =  If409768b648a33a7ed878a070d4f6251['h005e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002f5] =  If409768b648a33a7ed878a070d4f6251['h005ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002f6] =  If409768b648a33a7ed878a070d4f6251['h005ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002f7] =  If409768b648a33a7ed878a070d4f6251['h005ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002f8] =  If409768b648a33a7ed878a070d4f6251['h005f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002f9] =  If409768b648a33a7ed878a070d4f6251['h005f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002fa] =  If409768b648a33a7ed878a070d4f6251['h005f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002fb] =  If409768b648a33a7ed878a070d4f6251['h005f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002fc] =  If409768b648a33a7ed878a070d4f6251['h005f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002fd] =  If409768b648a33a7ed878a070d4f6251['h005fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002fe] =  If409768b648a33a7ed878a070d4f6251['h005fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h002ff] =  If409768b648a33a7ed878a070d4f6251['h005fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00300] =  If409768b648a33a7ed878a070d4f6251['h00600] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00301] =  If409768b648a33a7ed878a070d4f6251['h00602] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00302] =  If409768b648a33a7ed878a070d4f6251['h00604] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00303] =  If409768b648a33a7ed878a070d4f6251['h00606] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00304] =  If409768b648a33a7ed878a070d4f6251['h00608] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00305] =  If409768b648a33a7ed878a070d4f6251['h0060a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00306] =  If409768b648a33a7ed878a070d4f6251['h0060c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00307] =  If409768b648a33a7ed878a070d4f6251['h0060e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00308] =  If409768b648a33a7ed878a070d4f6251['h00610] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00309] =  If409768b648a33a7ed878a070d4f6251['h00612] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0030a] =  If409768b648a33a7ed878a070d4f6251['h00614] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0030b] =  If409768b648a33a7ed878a070d4f6251['h00616] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0030c] =  If409768b648a33a7ed878a070d4f6251['h00618] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0030d] =  If409768b648a33a7ed878a070d4f6251['h0061a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0030e] =  If409768b648a33a7ed878a070d4f6251['h0061c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0030f] =  If409768b648a33a7ed878a070d4f6251['h0061e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00310] =  If409768b648a33a7ed878a070d4f6251['h00620] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00311] =  If409768b648a33a7ed878a070d4f6251['h00622] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00312] =  If409768b648a33a7ed878a070d4f6251['h00624] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00313] =  If409768b648a33a7ed878a070d4f6251['h00626] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00314] =  If409768b648a33a7ed878a070d4f6251['h00628] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00315] =  If409768b648a33a7ed878a070d4f6251['h0062a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00316] =  If409768b648a33a7ed878a070d4f6251['h0062c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00317] =  If409768b648a33a7ed878a070d4f6251['h0062e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00318] =  If409768b648a33a7ed878a070d4f6251['h00630] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00319] =  If409768b648a33a7ed878a070d4f6251['h00632] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0031a] =  If409768b648a33a7ed878a070d4f6251['h00634] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0031b] =  If409768b648a33a7ed878a070d4f6251['h00636] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0031c] =  If409768b648a33a7ed878a070d4f6251['h00638] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0031d] =  If409768b648a33a7ed878a070d4f6251['h0063a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0031e] =  If409768b648a33a7ed878a070d4f6251['h0063c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0031f] =  If409768b648a33a7ed878a070d4f6251['h0063e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00320] =  If409768b648a33a7ed878a070d4f6251['h00640] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00321] =  If409768b648a33a7ed878a070d4f6251['h00642] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00322] =  If409768b648a33a7ed878a070d4f6251['h00644] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00323] =  If409768b648a33a7ed878a070d4f6251['h00646] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00324] =  If409768b648a33a7ed878a070d4f6251['h00648] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00325] =  If409768b648a33a7ed878a070d4f6251['h0064a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00326] =  If409768b648a33a7ed878a070d4f6251['h0064c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00327] =  If409768b648a33a7ed878a070d4f6251['h0064e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00328] =  If409768b648a33a7ed878a070d4f6251['h00650] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00329] =  If409768b648a33a7ed878a070d4f6251['h00652] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0032a] =  If409768b648a33a7ed878a070d4f6251['h00654] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0032b] =  If409768b648a33a7ed878a070d4f6251['h00656] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0032c] =  If409768b648a33a7ed878a070d4f6251['h00658] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0032d] =  If409768b648a33a7ed878a070d4f6251['h0065a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0032e] =  If409768b648a33a7ed878a070d4f6251['h0065c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0032f] =  If409768b648a33a7ed878a070d4f6251['h0065e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00330] =  If409768b648a33a7ed878a070d4f6251['h00660] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00331] =  If409768b648a33a7ed878a070d4f6251['h00662] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00332] =  If409768b648a33a7ed878a070d4f6251['h00664] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00333] =  If409768b648a33a7ed878a070d4f6251['h00666] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00334] =  If409768b648a33a7ed878a070d4f6251['h00668] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00335] =  If409768b648a33a7ed878a070d4f6251['h0066a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00336] =  If409768b648a33a7ed878a070d4f6251['h0066c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00337] =  If409768b648a33a7ed878a070d4f6251['h0066e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00338] =  If409768b648a33a7ed878a070d4f6251['h00670] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00339] =  If409768b648a33a7ed878a070d4f6251['h00672] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0033a] =  If409768b648a33a7ed878a070d4f6251['h00674] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0033b] =  If409768b648a33a7ed878a070d4f6251['h00676] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0033c] =  If409768b648a33a7ed878a070d4f6251['h00678] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0033d] =  If409768b648a33a7ed878a070d4f6251['h0067a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0033e] =  If409768b648a33a7ed878a070d4f6251['h0067c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0033f] =  If409768b648a33a7ed878a070d4f6251['h0067e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00340] =  If409768b648a33a7ed878a070d4f6251['h00680] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00341] =  If409768b648a33a7ed878a070d4f6251['h00682] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00342] =  If409768b648a33a7ed878a070d4f6251['h00684] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00343] =  If409768b648a33a7ed878a070d4f6251['h00686] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00344] =  If409768b648a33a7ed878a070d4f6251['h00688] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00345] =  If409768b648a33a7ed878a070d4f6251['h0068a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00346] =  If409768b648a33a7ed878a070d4f6251['h0068c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00347] =  If409768b648a33a7ed878a070d4f6251['h0068e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00348] =  If409768b648a33a7ed878a070d4f6251['h00690] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00349] =  If409768b648a33a7ed878a070d4f6251['h00692] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0034a] =  If409768b648a33a7ed878a070d4f6251['h00694] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0034b] =  If409768b648a33a7ed878a070d4f6251['h00696] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0034c] =  If409768b648a33a7ed878a070d4f6251['h00698] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0034d] =  If409768b648a33a7ed878a070d4f6251['h0069a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0034e] =  If409768b648a33a7ed878a070d4f6251['h0069c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0034f] =  If409768b648a33a7ed878a070d4f6251['h0069e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00350] =  If409768b648a33a7ed878a070d4f6251['h006a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00351] =  If409768b648a33a7ed878a070d4f6251['h006a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00352] =  If409768b648a33a7ed878a070d4f6251['h006a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00353] =  If409768b648a33a7ed878a070d4f6251['h006a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00354] =  If409768b648a33a7ed878a070d4f6251['h006a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00355] =  If409768b648a33a7ed878a070d4f6251['h006aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00356] =  If409768b648a33a7ed878a070d4f6251['h006ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00357] =  If409768b648a33a7ed878a070d4f6251['h006ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00358] =  If409768b648a33a7ed878a070d4f6251['h006b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00359] =  If409768b648a33a7ed878a070d4f6251['h006b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0035a] =  If409768b648a33a7ed878a070d4f6251['h006b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0035b] =  If409768b648a33a7ed878a070d4f6251['h006b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0035c] =  If409768b648a33a7ed878a070d4f6251['h006b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0035d] =  If409768b648a33a7ed878a070d4f6251['h006ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0035e] =  If409768b648a33a7ed878a070d4f6251['h006bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0035f] =  If409768b648a33a7ed878a070d4f6251['h006be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00360] =  If409768b648a33a7ed878a070d4f6251['h006c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00361] =  If409768b648a33a7ed878a070d4f6251['h006c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00362] =  If409768b648a33a7ed878a070d4f6251['h006c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00363] =  If409768b648a33a7ed878a070d4f6251['h006c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00364] =  If409768b648a33a7ed878a070d4f6251['h006c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00365] =  If409768b648a33a7ed878a070d4f6251['h006ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00366] =  If409768b648a33a7ed878a070d4f6251['h006cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00367] =  If409768b648a33a7ed878a070d4f6251['h006ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00368] =  If409768b648a33a7ed878a070d4f6251['h006d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00369] =  If409768b648a33a7ed878a070d4f6251['h006d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0036a] =  If409768b648a33a7ed878a070d4f6251['h006d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0036b] =  If409768b648a33a7ed878a070d4f6251['h006d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0036c] =  If409768b648a33a7ed878a070d4f6251['h006d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0036d] =  If409768b648a33a7ed878a070d4f6251['h006da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0036e] =  If409768b648a33a7ed878a070d4f6251['h006dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0036f] =  If409768b648a33a7ed878a070d4f6251['h006de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00370] =  If409768b648a33a7ed878a070d4f6251['h006e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00371] =  If409768b648a33a7ed878a070d4f6251['h006e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00372] =  If409768b648a33a7ed878a070d4f6251['h006e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00373] =  If409768b648a33a7ed878a070d4f6251['h006e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00374] =  If409768b648a33a7ed878a070d4f6251['h006e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00375] =  If409768b648a33a7ed878a070d4f6251['h006ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00376] =  If409768b648a33a7ed878a070d4f6251['h006ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00377] =  If409768b648a33a7ed878a070d4f6251['h006ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00378] =  If409768b648a33a7ed878a070d4f6251['h006f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00379] =  If409768b648a33a7ed878a070d4f6251['h006f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0037a] =  If409768b648a33a7ed878a070d4f6251['h006f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0037b] =  If409768b648a33a7ed878a070d4f6251['h006f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0037c] =  If409768b648a33a7ed878a070d4f6251['h006f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0037d] =  If409768b648a33a7ed878a070d4f6251['h006fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0037e] =  If409768b648a33a7ed878a070d4f6251['h006fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0037f] =  If409768b648a33a7ed878a070d4f6251['h006fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00380] =  If409768b648a33a7ed878a070d4f6251['h00700] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00381] =  If409768b648a33a7ed878a070d4f6251['h00702] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00382] =  If409768b648a33a7ed878a070d4f6251['h00704] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00383] =  If409768b648a33a7ed878a070d4f6251['h00706] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00384] =  If409768b648a33a7ed878a070d4f6251['h00708] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00385] =  If409768b648a33a7ed878a070d4f6251['h0070a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00386] =  If409768b648a33a7ed878a070d4f6251['h0070c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00387] =  If409768b648a33a7ed878a070d4f6251['h0070e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00388] =  If409768b648a33a7ed878a070d4f6251['h00710] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00389] =  If409768b648a33a7ed878a070d4f6251['h00712] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0038a] =  If409768b648a33a7ed878a070d4f6251['h00714] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0038b] =  If409768b648a33a7ed878a070d4f6251['h00716] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0038c] =  If409768b648a33a7ed878a070d4f6251['h00718] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0038d] =  If409768b648a33a7ed878a070d4f6251['h0071a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0038e] =  If409768b648a33a7ed878a070d4f6251['h0071c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0038f] =  If409768b648a33a7ed878a070d4f6251['h0071e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00390] =  If409768b648a33a7ed878a070d4f6251['h00720] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00391] =  If409768b648a33a7ed878a070d4f6251['h00722] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00392] =  If409768b648a33a7ed878a070d4f6251['h00724] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00393] =  If409768b648a33a7ed878a070d4f6251['h00726] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00394] =  If409768b648a33a7ed878a070d4f6251['h00728] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00395] =  If409768b648a33a7ed878a070d4f6251['h0072a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00396] =  If409768b648a33a7ed878a070d4f6251['h0072c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00397] =  If409768b648a33a7ed878a070d4f6251['h0072e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00398] =  If409768b648a33a7ed878a070d4f6251['h00730] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00399] =  If409768b648a33a7ed878a070d4f6251['h00732] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0039a] =  If409768b648a33a7ed878a070d4f6251['h00734] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0039b] =  If409768b648a33a7ed878a070d4f6251['h00736] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0039c] =  If409768b648a33a7ed878a070d4f6251['h00738] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0039d] =  If409768b648a33a7ed878a070d4f6251['h0073a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0039e] =  If409768b648a33a7ed878a070d4f6251['h0073c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0039f] =  If409768b648a33a7ed878a070d4f6251['h0073e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003a0] =  If409768b648a33a7ed878a070d4f6251['h00740] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003a1] =  If409768b648a33a7ed878a070d4f6251['h00742] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003a2] =  If409768b648a33a7ed878a070d4f6251['h00744] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003a3] =  If409768b648a33a7ed878a070d4f6251['h00746] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003a4] =  If409768b648a33a7ed878a070d4f6251['h00748] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003a5] =  If409768b648a33a7ed878a070d4f6251['h0074a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003a6] =  If409768b648a33a7ed878a070d4f6251['h0074c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003a7] =  If409768b648a33a7ed878a070d4f6251['h0074e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003a8] =  If409768b648a33a7ed878a070d4f6251['h00750] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003a9] =  If409768b648a33a7ed878a070d4f6251['h00752] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003aa] =  If409768b648a33a7ed878a070d4f6251['h00754] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ab] =  If409768b648a33a7ed878a070d4f6251['h00756] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ac] =  If409768b648a33a7ed878a070d4f6251['h00758] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ad] =  If409768b648a33a7ed878a070d4f6251['h0075a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ae] =  If409768b648a33a7ed878a070d4f6251['h0075c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003af] =  If409768b648a33a7ed878a070d4f6251['h0075e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003b0] =  If409768b648a33a7ed878a070d4f6251['h00760] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003b1] =  If409768b648a33a7ed878a070d4f6251['h00762] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003b2] =  If409768b648a33a7ed878a070d4f6251['h00764] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003b3] =  If409768b648a33a7ed878a070d4f6251['h00766] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003b4] =  If409768b648a33a7ed878a070d4f6251['h00768] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003b5] =  If409768b648a33a7ed878a070d4f6251['h0076a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003b6] =  If409768b648a33a7ed878a070d4f6251['h0076c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003b7] =  If409768b648a33a7ed878a070d4f6251['h0076e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003b8] =  If409768b648a33a7ed878a070d4f6251['h00770] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003b9] =  If409768b648a33a7ed878a070d4f6251['h00772] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ba] =  If409768b648a33a7ed878a070d4f6251['h00774] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003bb] =  If409768b648a33a7ed878a070d4f6251['h00776] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003bc] =  If409768b648a33a7ed878a070d4f6251['h00778] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003bd] =  If409768b648a33a7ed878a070d4f6251['h0077a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003be] =  If409768b648a33a7ed878a070d4f6251['h0077c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003bf] =  If409768b648a33a7ed878a070d4f6251['h0077e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003c0] =  If409768b648a33a7ed878a070d4f6251['h00780] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003c1] =  If409768b648a33a7ed878a070d4f6251['h00782] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003c2] =  If409768b648a33a7ed878a070d4f6251['h00784] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003c3] =  If409768b648a33a7ed878a070d4f6251['h00786] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003c4] =  If409768b648a33a7ed878a070d4f6251['h00788] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003c5] =  If409768b648a33a7ed878a070d4f6251['h0078a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003c6] =  If409768b648a33a7ed878a070d4f6251['h0078c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003c7] =  If409768b648a33a7ed878a070d4f6251['h0078e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003c8] =  If409768b648a33a7ed878a070d4f6251['h00790] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003c9] =  If409768b648a33a7ed878a070d4f6251['h00792] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ca] =  If409768b648a33a7ed878a070d4f6251['h00794] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003cb] =  If409768b648a33a7ed878a070d4f6251['h00796] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003cc] =  If409768b648a33a7ed878a070d4f6251['h00798] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003cd] =  If409768b648a33a7ed878a070d4f6251['h0079a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ce] =  If409768b648a33a7ed878a070d4f6251['h0079c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003cf] =  If409768b648a33a7ed878a070d4f6251['h0079e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003d0] =  If409768b648a33a7ed878a070d4f6251['h007a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003d1] =  If409768b648a33a7ed878a070d4f6251['h007a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003d2] =  If409768b648a33a7ed878a070d4f6251['h007a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003d3] =  If409768b648a33a7ed878a070d4f6251['h007a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003d4] =  If409768b648a33a7ed878a070d4f6251['h007a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003d5] =  If409768b648a33a7ed878a070d4f6251['h007aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003d6] =  If409768b648a33a7ed878a070d4f6251['h007ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003d7] =  If409768b648a33a7ed878a070d4f6251['h007ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003d8] =  If409768b648a33a7ed878a070d4f6251['h007b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003d9] =  If409768b648a33a7ed878a070d4f6251['h007b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003da] =  If409768b648a33a7ed878a070d4f6251['h007b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003db] =  If409768b648a33a7ed878a070d4f6251['h007b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003dc] =  If409768b648a33a7ed878a070d4f6251['h007b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003dd] =  If409768b648a33a7ed878a070d4f6251['h007ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003de] =  If409768b648a33a7ed878a070d4f6251['h007bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003df] =  If409768b648a33a7ed878a070d4f6251['h007be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003e0] =  If409768b648a33a7ed878a070d4f6251['h007c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003e1] =  If409768b648a33a7ed878a070d4f6251['h007c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003e2] =  If409768b648a33a7ed878a070d4f6251['h007c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003e3] =  If409768b648a33a7ed878a070d4f6251['h007c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003e4] =  If409768b648a33a7ed878a070d4f6251['h007c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003e5] =  If409768b648a33a7ed878a070d4f6251['h007ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003e6] =  If409768b648a33a7ed878a070d4f6251['h007cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003e7] =  If409768b648a33a7ed878a070d4f6251['h007ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003e8] =  If409768b648a33a7ed878a070d4f6251['h007d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003e9] =  If409768b648a33a7ed878a070d4f6251['h007d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ea] =  If409768b648a33a7ed878a070d4f6251['h007d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003eb] =  If409768b648a33a7ed878a070d4f6251['h007d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ec] =  If409768b648a33a7ed878a070d4f6251['h007d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ed] =  If409768b648a33a7ed878a070d4f6251['h007da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ee] =  If409768b648a33a7ed878a070d4f6251['h007dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ef] =  If409768b648a33a7ed878a070d4f6251['h007de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003f0] =  If409768b648a33a7ed878a070d4f6251['h007e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003f1] =  If409768b648a33a7ed878a070d4f6251['h007e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003f2] =  If409768b648a33a7ed878a070d4f6251['h007e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003f3] =  If409768b648a33a7ed878a070d4f6251['h007e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003f4] =  If409768b648a33a7ed878a070d4f6251['h007e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003f5] =  If409768b648a33a7ed878a070d4f6251['h007ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003f6] =  If409768b648a33a7ed878a070d4f6251['h007ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003f7] =  If409768b648a33a7ed878a070d4f6251['h007ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003f8] =  If409768b648a33a7ed878a070d4f6251['h007f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003f9] =  If409768b648a33a7ed878a070d4f6251['h007f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003fa] =  If409768b648a33a7ed878a070d4f6251['h007f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003fb] =  If409768b648a33a7ed878a070d4f6251['h007f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003fc] =  If409768b648a33a7ed878a070d4f6251['h007f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003fd] =  If409768b648a33a7ed878a070d4f6251['h007fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003fe] =  If409768b648a33a7ed878a070d4f6251['h007fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h003ff] =  If409768b648a33a7ed878a070d4f6251['h007fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00400] =  If409768b648a33a7ed878a070d4f6251['h00800] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00401] =  If409768b648a33a7ed878a070d4f6251['h00802] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00402] =  If409768b648a33a7ed878a070d4f6251['h00804] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00403] =  If409768b648a33a7ed878a070d4f6251['h00806] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00404] =  If409768b648a33a7ed878a070d4f6251['h00808] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00405] =  If409768b648a33a7ed878a070d4f6251['h0080a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00406] =  If409768b648a33a7ed878a070d4f6251['h0080c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00407] =  If409768b648a33a7ed878a070d4f6251['h0080e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00408] =  If409768b648a33a7ed878a070d4f6251['h00810] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00409] =  If409768b648a33a7ed878a070d4f6251['h00812] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0040a] =  If409768b648a33a7ed878a070d4f6251['h00814] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0040b] =  If409768b648a33a7ed878a070d4f6251['h00816] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0040c] =  If409768b648a33a7ed878a070d4f6251['h00818] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0040d] =  If409768b648a33a7ed878a070d4f6251['h0081a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0040e] =  If409768b648a33a7ed878a070d4f6251['h0081c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0040f] =  If409768b648a33a7ed878a070d4f6251['h0081e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00410] =  If409768b648a33a7ed878a070d4f6251['h00820] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00411] =  If409768b648a33a7ed878a070d4f6251['h00822] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00412] =  If409768b648a33a7ed878a070d4f6251['h00824] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00413] =  If409768b648a33a7ed878a070d4f6251['h00826] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00414] =  If409768b648a33a7ed878a070d4f6251['h00828] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00415] =  If409768b648a33a7ed878a070d4f6251['h0082a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00416] =  If409768b648a33a7ed878a070d4f6251['h0082c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00417] =  If409768b648a33a7ed878a070d4f6251['h0082e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00418] =  If409768b648a33a7ed878a070d4f6251['h00830] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00419] =  If409768b648a33a7ed878a070d4f6251['h00832] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0041a] =  If409768b648a33a7ed878a070d4f6251['h00834] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0041b] =  If409768b648a33a7ed878a070d4f6251['h00836] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0041c] =  If409768b648a33a7ed878a070d4f6251['h00838] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0041d] =  If409768b648a33a7ed878a070d4f6251['h0083a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0041e] =  If409768b648a33a7ed878a070d4f6251['h0083c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0041f] =  If409768b648a33a7ed878a070d4f6251['h0083e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00420] =  If409768b648a33a7ed878a070d4f6251['h00840] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00421] =  If409768b648a33a7ed878a070d4f6251['h00842] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00422] =  If409768b648a33a7ed878a070d4f6251['h00844] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00423] =  If409768b648a33a7ed878a070d4f6251['h00846] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00424] =  If409768b648a33a7ed878a070d4f6251['h00848] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00425] =  If409768b648a33a7ed878a070d4f6251['h0084a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00426] =  If409768b648a33a7ed878a070d4f6251['h0084c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00427] =  If409768b648a33a7ed878a070d4f6251['h0084e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00428] =  If409768b648a33a7ed878a070d4f6251['h00850] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00429] =  If409768b648a33a7ed878a070d4f6251['h00852] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0042a] =  If409768b648a33a7ed878a070d4f6251['h00854] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0042b] =  If409768b648a33a7ed878a070d4f6251['h00856] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0042c] =  If409768b648a33a7ed878a070d4f6251['h00858] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0042d] =  If409768b648a33a7ed878a070d4f6251['h0085a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0042e] =  If409768b648a33a7ed878a070d4f6251['h0085c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0042f] =  If409768b648a33a7ed878a070d4f6251['h0085e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00430] =  If409768b648a33a7ed878a070d4f6251['h00860] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00431] =  If409768b648a33a7ed878a070d4f6251['h00862] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00432] =  If409768b648a33a7ed878a070d4f6251['h00864] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00433] =  If409768b648a33a7ed878a070d4f6251['h00866] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00434] =  If409768b648a33a7ed878a070d4f6251['h00868] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00435] =  If409768b648a33a7ed878a070d4f6251['h0086a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00436] =  If409768b648a33a7ed878a070d4f6251['h0086c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00437] =  If409768b648a33a7ed878a070d4f6251['h0086e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00438] =  If409768b648a33a7ed878a070d4f6251['h00870] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00439] =  If409768b648a33a7ed878a070d4f6251['h00872] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0043a] =  If409768b648a33a7ed878a070d4f6251['h00874] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0043b] =  If409768b648a33a7ed878a070d4f6251['h00876] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0043c] =  If409768b648a33a7ed878a070d4f6251['h00878] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0043d] =  If409768b648a33a7ed878a070d4f6251['h0087a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0043e] =  If409768b648a33a7ed878a070d4f6251['h0087c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0043f] =  If409768b648a33a7ed878a070d4f6251['h0087e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00440] =  If409768b648a33a7ed878a070d4f6251['h00880] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00441] =  If409768b648a33a7ed878a070d4f6251['h00882] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00442] =  If409768b648a33a7ed878a070d4f6251['h00884] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00443] =  If409768b648a33a7ed878a070d4f6251['h00886] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00444] =  If409768b648a33a7ed878a070d4f6251['h00888] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00445] =  If409768b648a33a7ed878a070d4f6251['h0088a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00446] =  If409768b648a33a7ed878a070d4f6251['h0088c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00447] =  If409768b648a33a7ed878a070d4f6251['h0088e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00448] =  If409768b648a33a7ed878a070d4f6251['h00890] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00449] =  If409768b648a33a7ed878a070d4f6251['h00892] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0044a] =  If409768b648a33a7ed878a070d4f6251['h00894] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0044b] =  If409768b648a33a7ed878a070d4f6251['h00896] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0044c] =  If409768b648a33a7ed878a070d4f6251['h00898] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0044d] =  If409768b648a33a7ed878a070d4f6251['h0089a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0044e] =  If409768b648a33a7ed878a070d4f6251['h0089c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0044f] =  If409768b648a33a7ed878a070d4f6251['h0089e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00450] =  If409768b648a33a7ed878a070d4f6251['h008a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00451] =  If409768b648a33a7ed878a070d4f6251['h008a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00452] =  If409768b648a33a7ed878a070d4f6251['h008a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00453] =  If409768b648a33a7ed878a070d4f6251['h008a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00454] =  If409768b648a33a7ed878a070d4f6251['h008a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00455] =  If409768b648a33a7ed878a070d4f6251['h008aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00456] =  If409768b648a33a7ed878a070d4f6251['h008ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00457] =  If409768b648a33a7ed878a070d4f6251['h008ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00458] =  If409768b648a33a7ed878a070d4f6251['h008b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00459] =  If409768b648a33a7ed878a070d4f6251['h008b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0045a] =  If409768b648a33a7ed878a070d4f6251['h008b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0045b] =  If409768b648a33a7ed878a070d4f6251['h008b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0045c] =  If409768b648a33a7ed878a070d4f6251['h008b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0045d] =  If409768b648a33a7ed878a070d4f6251['h008ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0045e] =  If409768b648a33a7ed878a070d4f6251['h008bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0045f] =  If409768b648a33a7ed878a070d4f6251['h008be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00460] =  If409768b648a33a7ed878a070d4f6251['h008c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00461] =  If409768b648a33a7ed878a070d4f6251['h008c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00462] =  If409768b648a33a7ed878a070d4f6251['h008c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00463] =  If409768b648a33a7ed878a070d4f6251['h008c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00464] =  If409768b648a33a7ed878a070d4f6251['h008c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00465] =  If409768b648a33a7ed878a070d4f6251['h008ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00466] =  If409768b648a33a7ed878a070d4f6251['h008cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00467] =  If409768b648a33a7ed878a070d4f6251['h008ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00468] =  If409768b648a33a7ed878a070d4f6251['h008d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00469] =  If409768b648a33a7ed878a070d4f6251['h008d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0046a] =  If409768b648a33a7ed878a070d4f6251['h008d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0046b] =  If409768b648a33a7ed878a070d4f6251['h008d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0046c] =  If409768b648a33a7ed878a070d4f6251['h008d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0046d] =  If409768b648a33a7ed878a070d4f6251['h008da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0046e] =  If409768b648a33a7ed878a070d4f6251['h008dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0046f] =  If409768b648a33a7ed878a070d4f6251['h008de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00470] =  If409768b648a33a7ed878a070d4f6251['h008e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00471] =  If409768b648a33a7ed878a070d4f6251['h008e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00472] =  If409768b648a33a7ed878a070d4f6251['h008e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00473] =  If409768b648a33a7ed878a070d4f6251['h008e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00474] =  If409768b648a33a7ed878a070d4f6251['h008e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00475] =  If409768b648a33a7ed878a070d4f6251['h008ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00476] =  If409768b648a33a7ed878a070d4f6251['h008ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00477] =  If409768b648a33a7ed878a070d4f6251['h008ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00478] =  If409768b648a33a7ed878a070d4f6251['h008f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00479] =  If409768b648a33a7ed878a070d4f6251['h008f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0047a] =  If409768b648a33a7ed878a070d4f6251['h008f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0047b] =  If409768b648a33a7ed878a070d4f6251['h008f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0047c] =  If409768b648a33a7ed878a070d4f6251['h008f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0047d] =  If409768b648a33a7ed878a070d4f6251['h008fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0047e] =  If409768b648a33a7ed878a070d4f6251['h008fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0047f] =  If409768b648a33a7ed878a070d4f6251['h008fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00480] =  If409768b648a33a7ed878a070d4f6251['h00900] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00481] =  If409768b648a33a7ed878a070d4f6251['h00902] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00482] =  If409768b648a33a7ed878a070d4f6251['h00904] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00483] =  If409768b648a33a7ed878a070d4f6251['h00906] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00484] =  If409768b648a33a7ed878a070d4f6251['h00908] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00485] =  If409768b648a33a7ed878a070d4f6251['h0090a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00486] =  If409768b648a33a7ed878a070d4f6251['h0090c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00487] =  If409768b648a33a7ed878a070d4f6251['h0090e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00488] =  If409768b648a33a7ed878a070d4f6251['h00910] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00489] =  If409768b648a33a7ed878a070d4f6251['h00912] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0048a] =  If409768b648a33a7ed878a070d4f6251['h00914] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0048b] =  If409768b648a33a7ed878a070d4f6251['h00916] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0048c] =  If409768b648a33a7ed878a070d4f6251['h00918] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0048d] =  If409768b648a33a7ed878a070d4f6251['h0091a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0048e] =  If409768b648a33a7ed878a070d4f6251['h0091c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0048f] =  If409768b648a33a7ed878a070d4f6251['h0091e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00490] =  If409768b648a33a7ed878a070d4f6251['h00920] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00491] =  If409768b648a33a7ed878a070d4f6251['h00922] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00492] =  If409768b648a33a7ed878a070d4f6251['h00924] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00493] =  If409768b648a33a7ed878a070d4f6251['h00926] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00494] =  If409768b648a33a7ed878a070d4f6251['h00928] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00495] =  If409768b648a33a7ed878a070d4f6251['h0092a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00496] =  If409768b648a33a7ed878a070d4f6251['h0092c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00497] =  If409768b648a33a7ed878a070d4f6251['h0092e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00498] =  If409768b648a33a7ed878a070d4f6251['h00930] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00499] =  If409768b648a33a7ed878a070d4f6251['h00932] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0049a] =  If409768b648a33a7ed878a070d4f6251['h00934] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0049b] =  If409768b648a33a7ed878a070d4f6251['h00936] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0049c] =  If409768b648a33a7ed878a070d4f6251['h00938] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0049d] =  If409768b648a33a7ed878a070d4f6251['h0093a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0049e] =  If409768b648a33a7ed878a070d4f6251['h0093c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0049f] =  If409768b648a33a7ed878a070d4f6251['h0093e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004a0] =  If409768b648a33a7ed878a070d4f6251['h00940] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004a1] =  If409768b648a33a7ed878a070d4f6251['h00942] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004a2] =  If409768b648a33a7ed878a070d4f6251['h00944] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004a3] =  If409768b648a33a7ed878a070d4f6251['h00946] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004a4] =  If409768b648a33a7ed878a070d4f6251['h00948] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004a5] =  If409768b648a33a7ed878a070d4f6251['h0094a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004a6] =  If409768b648a33a7ed878a070d4f6251['h0094c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004a7] =  If409768b648a33a7ed878a070d4f6251['h0094e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004a8] =  If409768b648a33a7ed878a070d4f6251['h00950] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004a9] =  If409768b648a33a7ed878a070d4f6251['h00952] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004aa] =  If409768b648a33a7ed878a070d4f6251['h00954] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ab] =  If409768b648a33a7ed878a070d4f6251['h00956] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ac] =  If409768b648a33a7ed878a070d4f6251['h00958] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ad] =  If409768b648a33a7ed878a070d4f6251['h0095a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ae] =  If409768b648a33a7ed878a070d4f6251['h0095c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004af] =  If409768b648a33a7ed878a070d4f6251['h0095e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004b0] =  If409768b648a33a7ed878a070d4f6251['h00960] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004b1] =  If409768b648a33a7ed878a070d4f6251['h00962] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004b2] =  If409768b648a33a7ed878a070d4f6251['h00964] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004b3] =  If409768b648a33a7ed878a070d4f6251['h00966] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004b4] =  If409768b648a33a7ed878a070d4f6251['h00968] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004b5] =  If409768b648a33a7ed878a070d4f6251['h0096a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004b6] =  If409768b648a33a7ed878a070d4f6251['h0096c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004b7] =  If409768b648a33a7ed878a070d4f6251['h0096e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004b8] =  If409768b648a33a7ed878a070d4f6251['h00970] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004b9] =  If409768b648a33a7ed878a070d4f6251['h00972] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ba] =  If409768b648a33a7ed878a070d4f6251['h00974] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004bb] =  If409768b648a33a7ed878a070d4f6251['h00976] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004bc] =  If409768b648a33a7ed878a070d4f6251['h00978] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004bd] =  If409768b648a33a7ed878a070d4f6251['h0097a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004be] =  If409768b648a33a7ed878a070d4f6251['h0097c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004bf] =  If409768b648a33a7ed878a070d4f6251['h0097e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004c0] =  If409768b648a33a7ed878a070d4f6251['h00980] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004c1] =  If409768b648a33a7ed878a070d4f6251['h00982] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004c2] =  If409768b648a33a7ed878a070d4f6251['h00984] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004c3] =  If409768b648a33a7ed878a070d4f6251['h00986] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004c4] =  If409768b648a33a7ed878a070d4f6251['h00988] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004c5] =  If409768b648a33a7ed878a070d4f6251['h0098a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004c6] =  If409768b648a33a7ed878a070d4f6251['h0098c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004c7] =  If409768b648a33a7ed878a070d4f6251['h0098e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004c8] =  If409768b648a33a7ed878a070d4f6251['h00990] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004c9] =  If409768b648a33a7ed878a070d4f6251['h00992] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ca] =  If409768b648a33a7ed878a070d4f6251['h00994] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004cb] =  If409768b648a33a7ed878a070d4f6251['h00996] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004cc] =  If409768b648a33a7ed878a070d4f6251['h00998] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004cd] =  If409768b648a33a7ed878a070d4f6251['h0099a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ce] =  If409768b648a33a7ed878a070d4f6251['h0099c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004cf] =  If409768b648a33a7ed878a070d4f6251['h0099e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004d0] =  If409768b648a33a7ed878a070d4f6251['h009a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004d1] =  If409768b648a33a7ed878a070d4f6251['h009a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004d2] =  If409768b648a33a7ed878a070d4f6251['h009a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004d3] =  If409768b648a33a7ed878a070d4f6251['h009a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004d4] =  If409768b648a33a7ed878a070d4f6251['h009a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004d5] =  If409768b648a33a7ed878a070d4f6251['h009aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004d6] =  If409768b648a33a7ed878a070d4f6251['h009ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004d7] =  If409768b648a33a7ed878a070d4f6251['h009ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004d8] =  If409768b648a33a7ed878a070d4f6251['h009b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004d9] =  If409768b648a33a7ed878a070d4f6251['h009b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004da] =  If409768b648a33a7ed878a070d4f6251['h009b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004db] =  If409768b648a33a7ed878a070d4f6251['h009b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004dc] =  If409768b648a33a7ed878a070d4f6251['h009b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004dd] =  If409768b648a33a7ed878a070d4f6251['h009ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004de] =  If409768b648a33a7ed878a070d4f6251['h009bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004df] =  If409768b648a33a7ed878a070d4f6251['h009be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004e0] =  If409768b648a33a7ed878a070d4f6251['h009c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004e1] =  If409768b648a33a7ed878a070d4f6251['h009c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004e2] =  If409768b648a33a7ed878a070d4f6251['h009c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004e3] =  If409768b648a33a7ed878a070d4f6251['h009c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004e4] =  If409768b648a33a7ed878a070d4f6251['h009c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004e5] =  If409768b648a33a7ed878a070d4f6251['h009ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004e6] =  If409768b648a33a7ed878a070d4f6251['h009cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004e7] =  If409768b648a33a7ed878a070d4f6251['h009ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004e8] =  If409768b648a33a7ed878a070d4f6251['h009d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004e9] =  If409768b648a33a7ed878a070d4f6251['h009d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ea] =  If409768b648a33a7ed878a070d4f6251['h009d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004eb] =  If409768b648a33a7ed878a070d4f6251['h009d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ec] =  If409768b648a33a7ed878a070d4f6251['h009d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ed] =  If409768b648a33a7ed878a070d4f6251['h009da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ee] =  If409768b648a33a7ed878a070d4f6251['h009dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ef] =  If409768b648a33a7ed878a070d4f6251['h009de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004f0] =  If409768b648a33a7ed878a070d4f6251['h009e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004f1] =  If409768b648a33a7ed878a070d4f6251['h009e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004f2] =  If409768b648a33a7ed878a070d4f6251['h009e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004f3] =  If409768b648a33a7ed878a070d4f6251['h009e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004f4] =  If409768b648a33a7ed878a070d4f6251['h009e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004f5] =  If409768b648a33a7ed878a070d4f6251['h009ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004f6] =  If409768b648a33a7ed878a070d4f6251['h009ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004f7] =  If409768b648a33a7ed878a070d4f6251['h009ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004f8] =  If409768b648a33a7ed878a070d4f6251['h009f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004f9] =  If409768b648a33a7ed878a070d4f6251['h009f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004fa] =  If409768b648a33a7ed878a070d4f6251['h009f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004fb] =  If409768b648a33a7ed878a070d4f6251['h009f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004fc] =  If409768b648a33a7ed878a070d4f6251['h009f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004fd] =  If409768b648a33a7ed878a070d4f6251['h009fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004fe] =  If409768b648a33a7ed878a070d4f6251['h009fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h004ff] =  If409768b648a33a7ed878a070d4f6251['h009fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00500] =  If409768b648a33a7ed878a070d4f6251['h00a00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00501] =  If409768b648a33a7ed878a070d4f6251['h00a02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00502] =  If409768b648a33a7ed878a070d4f6251['h00a04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00503] =  If409768b648a33a7ed878a070d4f6251['h00a06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00504] =  If409768b648a33a7ed878a070d4f6251['h00a08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00505] =  If409768b648a33a7ed878a070d4f6251['h00a0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00506] =  If409768b648a33a7ed878a070d4f6251['h00a0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00507] =  If409768b648a33a7ed878a070d4f6251['h00a0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00508] =  If409768b648a33a7ed878a070d4f6251['h00a10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00509] =  If409768b648a33a7ed878a070d4f6251['h00a12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0050a] =  If409768b648a33a7ed878a070d4f6251['h00a14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0050b] =  If409768b648a33a7ed878a070d4f6251['h00a16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0050c] =  If409768b648a33a7ed878a070d4f6251['h00a18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0050d] =  If409768b648a33a7ed878a070d4f6251['h00a1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0050e] =  If409768b648a33a7ed878a070d4f6251['h00a1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0050f] =  If409768b648a33a7ed878a070d4f6251['h00a1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00510] =  If409768b648a33a7ed878a070d4f6251['h00a20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00511] =  If409768b648a33a7ed878a070d4f6251['h00a22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00512] =  If409768b648a33a7ed878a070d4f6251['h00a24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00513] =  If409768b648a33a7ed878a070d4f6251['h00a26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00514] =  If409768b648a33a7ed878a070d4f6251['h00a28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00515] =  If409768b648a33a7ed878a070d4f6251['h00a2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00516] =  If409768b648a33a7ed878a070d4f6251['h00a2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00517] =  If409768b648a33a7ed878a070d4f6251['h00a2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00518] =  If409768b648a33a7ed878a070d4f6251['h00a30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00519] =  If409768b648a33a7ed878a070d4f6251['h00a32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0051a] =  If409768b648a33a7ed878a070d4f6251['h00a34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0051b] =  If409768b648a33a7ed878a070d4f6251['h00a36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0051c] =  If409768b648a33a7ed878a070d4f6251['h00a38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0051d] =  If409768b648a33a7ed878a070d4f6251['h00a3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0051e] =  If409768b648a33a7ed878a070d4f6251['h00a3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0051f] =  If409768b648a33a7ed878a070d4f6251['h00a3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00520] =  If409768b648a33a7ed878a070d4f6251['h00a40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00521] =  If409768b648a33a7ed878a070d4f6251['h00a42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00522] =  If409768b648a33a7ed878a070d4f6251['h00a44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00523] =  If409768b648a33a7ed878a070d4f6251['h00a46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00524] =  If409768b648a33a7ed878a070d4f6251['h00a48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00525] =  If409768b648a33a7ed878a070d4f6251['h00a4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00526] =  If409768b648a33a7ed878a070d4f6251['h00a4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00527] =  If409768b648a33a7ed878a070d4f6251['h00a4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00528] =  If409768b648a33a7ed878a070d4f6251['h00a50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00529] =  If409768b648a33a7ed878a070d4f6251['h00a52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0052a] =  If409768b648a33a7ed878a070d4f6251['h00a54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0052b] =  If409768b648a33a7ed878a070d4f6251['h00a56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0052c] =  If409768b648a33a7ed878a070d4f6251['h00a58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0052d] =  If409768b648a33a7ed878a070d4f6251['h00a5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0052e] =  If409768b648a33a7ed878a070d4f6251['h00a5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0052f] =  If409768b648a33a7ed878a070d4f6251['h00a5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00530] =  If409768b648a33a7ed878a070d4f6251['h00a60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00531] =  If409768b648a33a7ed878a070d4f6251['h00a62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00532] =  If409768b648a33a7ed878a070d4f6251['h00a64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00533] =  If409768b648a33a7ed878a070d4f6251['h00a66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00534] =  If409768b648a33a7ed878a070d4f6251['h00a68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00535] =  If409768b648a33a7ed878a070d4f6251['h00a6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00536] =  If409768b648a33a7ed878a070d4f6251['h00a6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00537] =  If409768b648a33a7ed878a070d4f6251['h00a6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00538] =  If409768b648a33a7ed878a070d4f6251['h00a70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00539] =  If409768b648a33a7ed878a070d4f6251['h00a72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0053a] =  If409768b648a33a7ed878a070d4f6251['h00a74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0053b] =  If409768b648a33a7ed878a070d4f6251['h00a76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0053c] =  If409768b648a33a7ed878a070d4f6251['h00a78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0053d] =  If409768b648a33a7ed878a070d4f6251['h00a7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0053e] =  If409768b648a33a7ed878a070d4f6251['h00a7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0053f] =  If409768b648a33a7ed878a070d4f6251['h00a7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00540] =  If409768b648a33a7ed878a070d4f6251['h00a80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00541] =  If409768b648a33a7ed878a070d4f6251['h00a82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00542] =  If409768b648a33a7ed878a070d4f6251['h00a84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00543] =  If409768b648a33a7ed878a070d4f6251['h00a86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00544] =  If409768b648a33a7ed878a070d4f6251['h00a88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00545] =  If409768b648a33a7ed878a070d4f6251['h00a8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00546] =  If409768b648a33a7ed878a070d4f6251['h00a8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00547] =  If409768b648a33a7ed878a070d4f6251['h00a8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00548] =  If409768b648a33a7ed878a070d4f6251['h00a90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00549] =  If409768b648a33a7ed878a070d4f6251['h00a92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0054a] =  If409768b648a33a7ed878a070d4f6251['h00a94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0054b] =  If409768b648a33a7ed878a070d4f6251['h00a96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0054c] =  If409768b648a33a7ed878a070d4f6251['h00a98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0054d] =  If409768b648a33a7ed878a070d4f6251['h00a9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0054e] =  If409768b648a33a7ed878a070d4f6251['h00a9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0054f] =  If409768b648a33a7ed878a070d4f6251['h00a9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00550] =  If409768b648a33a7ed878a070d4f6251['h00aa0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00551] =  If409768b648a33a7ed878a070d4f6251['h00aa2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00552] =  If409768b648a33a7ed878a070d4f6251['h00aa4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00553] =  If409768b648a33a7ed878a070d4f6251['h00aa6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00554] =  If409768b648a33a7ed878a070d4f6251['h00aa8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00555] =  If409768b648a33a7ed878a070d4f6251['h00aaa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00556] =  If409768b648a33a7ed878a070d4f6251['h00aac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00557] =  If409768b648a33a7ed878a070d4f6251['h00aae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00558] =  If409768b648a33a7ed878a070d4f6251['h00ab0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00559] =  If409768b648a33a7ed878a070d4f6251['h00ab2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0055a] =  If409768b648a33a7ed878a070d4f6251['h00ab4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0055b] =  If409768b648a33a7ed878a070d4f6251['h00ab6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0055c] =  If409768b648a33a7ed878a070d4f6251['h00ab8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0055d] =  If409768b648a33a7ed878a070d4f6251['h00aba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0055e] =  If409768b648a33a7ed878a070d4f6251['h00abc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0055f] =  If409768b648a33a7ed878a070d4f6251['h00abe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00560] =  If409768b648a33a7ed878a070d4f6251['h00ac0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00561] =  If409768b648a33a7ed878a070d4f6251['h00ac2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00562] =  If409768b648a33a7ed878a070d4f6251['h00ac4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00563] =  If409768b648a33a7ed878a070d4f6251['h00ac6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00564] =  If409768b648a33a7ed878a070d4f6251['h00ac8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00565] =  If409768b648a33a7ed878a070d4f6251['h00aca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00566] =  If409768b648a33a7ed878a070d4f6251['h00acc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00567] =  If409768b648a33a7ed878a070d4f6251['h00ace] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00568] =  If409768b648a33a7ed878a070d4f6251['h00ad0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00569] =  If409768b648a33a7ed878a070d4f6251['h00ad2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0056a] =  If409768b648a33a7ed878a070d4f6251['h00ad4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0056b] =  If409768b648a33a7ed878a070d4f6251['h00ad6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0056c] =  If409768b648a33a7ed878a070d4f6251['h00ad8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0056d] =  If409768b648a33a7ed878a070d4f6251['h00ada] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0056e] =  If409768b648a33a7ed878a070d4f6251['h00adc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0056f] =  If409768b648a33a7ed878a070d4f6251['h00ade] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00570] =  If409768b648a33a7ed878a070d4f6251['h00ae0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00571] =  If409768b648a33a7ed878a070d4f6251['h00ae2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00572] =  If409768b648a33a7ed878a070d4f6251['h00ae4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00573] =  If409768b648a33a7ed878a070d4f6251['h00ae6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00574] =  If409768b648a33a7ed878a070d4f6251['h00ae8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00575] =  If409768b648a33a7ed878a070d4f6251['h00aea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00576] =  If409768b648a33a7ed878a070d4f6251['h00aec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00577] =  If409768b648a33a7ed878a070d4f6251['h00aee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00578] =  If409768b648a33a7ed878a070d4f6251['h00af0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00579] =  If409768b648a33a7ed878a070d4f6251['h00af2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0057a] =  If409768b648a33a7ed878a070d4f6251['h00af4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0057b] =  If409768b648a33a7ed878a070d4f6251['h00af6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0057c] =  If409768b648a33a7ed878a070d4f6251['h00af8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0057d] =  If409768b648a33a7ed878a070d4f6251['h00afa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0057e] =  If409768b648a33a7ed878a070d4f6251['h00afc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0057f] =  If409768b648a33a7ed878a070d4f6251['h00afe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00580] =  If409768b648a33a7ed878a070d4f6251['h00b00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00581] =  If409768b648a33a7ed878a070d4f6251['h00b02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00582] =  If409768b648a33a7ed878a070d4f6251['h00b04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00583] =  If409768b648a33a7ed878a070d4f6251['h00b06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00584] =  If409768b648a33a7ed878a070d4f6251['h00b08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00585] =  If409768b648a33a7ed878a070d4f6251['h00b0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00586] =  If409768b648a33a7ed878a070d4f6251['h00b0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00587] =  If409768b648a33a7ed878a070d4f6251['h00b0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00588] =  If409768b648a33a7ed878a070d4f6251['h00b10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00589] =  If409768b648a33a7ed878a070d4f6251['h00b12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0058a] =  If409768b648a33a7ed878a070d4f6251['h00b14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0058b] =  If409768b648a33a7ed878a070d4f6251['h00b16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0058c] =  If409768b648a33a7ed878a070d4f6251['h00b18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0058d] =  If409768b648a33a7ed878a070d4f6251['h00b1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0058e] =  If409768b648a33a7ed878a070d4f6251['h00b1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0058f] =  If409768b648a33a7ed878a070d4f6251['h00b1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00590] =  If409768b648a33a7ed878a070d4f6251['h00b20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00591] =  If409768b648a33a7ed878a070d4f6251['h00b22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00592] =  If409768b648a33a7ed878a070d4f6251['h00b24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00593] =  If409768b648a33a7ed878a070d4f6251['h00b26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00594] =  If409768b648a33a7ed878a070d4f6251['h00b28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00595] =  If409768b648a33a7ed878a070d4f6251['h00b2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00596] =  If409768b648a33a7ed878a070d4f6251['h00b2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00597] =  If409768b648a33a7ed878a070d4f6251['h00b2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00598] =  If409768b648a33a7ed878a070d4f6251['h00b30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00599] =  If409768b648a33a7ed878a070d4f6251['h00b32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0059a] =  If409768b648a33a7ed878a070d4f6251['h00b34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0059b] =  If409768b648a33a7ed878a070d4f6251['h00b36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0059c] =  If409768b648a33a7ed878a070d4f6251['h00b38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0059d] =  If409768b648a33a7ed878a070d4f6251['h00b3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0059e] =  If409768b648a33a7ed878a070d4f6251['h00b3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0059f] =  If409768b648a33a7ed878a070d4f6251['h00b3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005a0] =  If409768b648a33a7ed878a070d4f6251['h00b40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005a1] =  If409768b648a33a7ed878a070d4f6251['h00b42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005a2] =  If409768b648a33a7ed878a070d4f6251['h00b44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005a3] =  If409768b648a33a7ed878a070d4f6251['h00b46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005a4] =  If409768b648a33a7ed878a070d4f6251['h00b48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005a5] =  If409768b648a33a7ed878a070d4f6251['h00b4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005a6] =  If409768b648a33a7ed878a070d4f6251['h00b4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005a7] =  If409768b648a33a7ed878a070d4f6251['h00b4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005a8] =  If409768b648a33a7ed878a070d4f6251['h00b50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005a9] =  If409768b648a33a7ed878a070d4f6251['h00b52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005aa] =  If409768b648a33a7ed878a070d4f6251['h00b54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ab] =  If409768b648a33a7ed878a070d4f6251['h00b56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ac] =  If409768b648a33a7ed878a070d4f6251['h00b58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ad] =  If409768b648a33a7ed878a070d4f6251['h00b5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ae] =  If409768b648a33a7ed878a070d4f6251['h00b5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005af] =  If409768b648a33a7ed878a070d4f6251['h00b5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005b0] =  If409768b648a33a7ed878a070d4f6251['h00b60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005b1] =  If409768b648a33a7ed878a070d4f6251['h00b62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005b2] =  If409768b648a33a7ed878a070d4f6251['h00b64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005b3] =  If409768b648a33a7ed878a070d4f6251['h00b66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005b4] =  If409768b648a33a7ed878a070d4f6251['h00b68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005b5] =  If409768b648a33a7ed878a070d4f6251['h00b6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005b6] =  If409768b648a33a7ed878a070d4f6251['h00b6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005b7] =  If409768b648a33a7ed878a070d4f6251['h00b6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005b8] =  If409768b648a33a7ed878a070d4f6251['h00b70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005b9] =  If409768b648a33a7ed878a070d4f6251['h00b72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ba] =  If409768b648a33a7ed878a070d4f6251['h00b74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005bb] =  If409768b648a33a7ed878a070d4f6251['h00b76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005bc] =  If409768b648a33a7ed878a070d4f6251['h00b78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005bd] =  If409768b648a33a7ed878a070d4f6251['h00b7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005be] =  If409768b648a33a7ed878a070d4f6251['h00b7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005bf] =  If409768b648a33a7ed878a070d4f6251['h00b7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005c0] =  If409768b648a33a7ed878a070d4f6251['h00b80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005c1] =  If409768b648a33a7ed878a070d4f6251['h00b82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005c2] =  If409768b648a33a7ed878a070d4f6251['h00b84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005c3] =  If409768b648a33a7ed878a070d4f6251['h00b86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005c4] =  If409768b648a33a7ed878a070d4f6251['h00b88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005c5] =  If409768b648a33a7ed878a070d4f6251['h00b8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005c6] =  If409768b648a33a7ed878a070d4f6251['h00b8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005c7] =  If409768b648a33a7ed878a070d4f6251['h00b8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005c8] =  If409768b648a33a7ed878a070d4f6251['h00b90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005c9] =  If409768b648a33a7ed878a070d4f6251['h00b92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ca] =  If409768b648a33a7ed878a070d4f6251['h00b94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005cb] =  If409768b648a33a7ed878a070d4f6251['h00b96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005cc] =  If409768b648a33a7ed878a070d4f6251['h00b98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005cd] =  If409768b648a33a7ed878a070d4f6251['h00b9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ce] =  If409768b648a33a7ed878a070d4f6251['h00b9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005cf] =  If409768b648a33a7ed878a070d4f6251['h00b9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005d0] =  If409768b648a33a7ed878a070d4f6251['h00ba0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005d1] =  If409768b648a33a7ed878a070d4f6251['h00ba2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005d2] =  If409768b648a33a7ed878a070d4f6251['h00ba4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005d3] =  If409768b648a33a7ed878a070d4f6251['h00ba6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005d4] =  If409768b648a33a7ed878a070d4f6251['h00ba8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005d5] =  If409768b648a33a7ed878a070d4f6251['h00baa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005d6] =  If409768b648a33a7ed878a070d4f6251['h00bac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005d7] =  If409768b648a33a7ed878a070d4f6251['h00bae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005d8] =  If409768b648a33a7ed878a070d4f6251['h00bb0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005d9] =  If409768b648a33a7ed878a070d4f6251['h00bb2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005da] =  If409768b648a33a7ed878a070d4f6251['h00bb4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005db] =  If409768b648a33a7ed878a070d4f6251['h00bb6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005dc] =  If409768b648a33a7ed878a070d4f6251['h00bb8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005dd] =  If409768b648a33a7ed878a070d4f6251['h00bba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005de] =  If409768b648a33a7ed878a070d4f6251['h00bbc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005df] =  If409768b648a33a7ed878a070d4f6251['h00bbe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005e0] =  If409768b648a33a7ed878a070d4f6251['h00bc0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005e1] =  If409768b648a33a7ed878a070d4f6251['h00bc2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005e2] =  If409768b648a33a7ed878a070d4f6251['h00bc4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005e3] =  If409768b648a33a7ed878a070d4f6251['h00bc6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005e4] =  If409768b648a33a7ed878a070d4f6251['h00bc8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005e5] =  If409768b648a33a7ed878a070d4f6251['h00bca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005e6] =  If409768b648a33a7ed878a070d4f6251['h00bcc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005e7] =  If409768b648a33a7ed878a070d4f6251['h00bce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005e8] =  If409768b648a33a7ed878a070d4f6251['h00bd0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005e9] =  If409768b648a33a7ed878a070d4f6251['h00bd2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ea] =  If409768b648a33a7ed878a070d4f6251['h00bd4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005eb] =  If409768b648a33a7ed878a070d4f6251['h00bd6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ec] =  If409768b648a33a7ed878a070d4f6251['h00bd8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ed] =  If409768b648a33a7ed878a070d4f6251['h00bda] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ee] =  If409768b648a33a7ed878a070d4f6251['h00bdc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ef] =  If409768b648a33a7ed878a070d4f6251['h00bde] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005f0] =  If409768b648a33a7ed878a070d4f6251['h00be0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005f1] =  If409768b648a33a7ed878a070d4f6251['h00be2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005f2] =  If409768b648a33a7ed878a070d4f6251['h00be4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005f3] =  If409768b648a33a7ed878a070d4f6251['h00be6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005f4] =  If409768b648a33a7ed878a070d4f6251['h00be8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005f5] =  If409768b648a33a7ed878a070d4f6251['h00bea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005f6] =  If409768b648a33a7ed878a070d4f6251['h00bec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005f7] =  If409768b648a33a7ed878a070d4f6251['h00bee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005f8] =  If409768b648a33a7ed878a070d4f6251['h00bf0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005f9] =  If409768b648a33a7ed878a070d4f6251['h00bf2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005fa] =  If409768b648a33a7ed878a070d4f6251['h00bf4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005fb] =  If409768b648a33a7ed878a070d4f6251['h00bf6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005fc] =  If409768b648a33a7ed878a070d4f6251['h00bf8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005fd] =  If409768b648a33a7ed878a070d4f6251['h00bfa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005fe] =  If409768b648a33a7ed878a070d4f6251['h00bfc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h005ff] =  If409768b648a33a7ed878a070d4f6251['h00bfe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00600] =  If409768b648a33a7ed878a070d4f6251['h00c00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00601] =  If409768b648a33a7ed878a070d4f6251['h00c02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00602] =  If409768b648a33a7ed878a070d4f6251['h00c04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00603] =  If409768b648a33a7ed878a070d4f6251['h00c06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00604] =  If409768b648a33a7ed878a070d4f6251['h00c08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00605] =  If409768b648a33a7ed878a070d4f6251['h00c0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00606] =  If409768b648a33a7ed878a070d4f6251['h00c0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00607] =  If409768b648a33a7ed878a070d4f6251['h00c0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00608] =  If409768b648a33a7ed878a070d4f6251['h00c10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00609] =  If409768b648a33a7ed878a070d4f6251['h00c12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0060a] =  If409768b648a33a7ed878a070d4f6251['h00c14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0060b] =  If409768b648a33a7ed878a070d4f6251['h00c16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0060c] =  If409768b648a33a7ed878a070d4f6251['h00c18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0060d] =  If409768b648a33a7ed878a070d4f6251['h00c1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0060e] =  If409768b648a33a7ed878a070d4f6251['h00c1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0060f] =  If409768b648a33a7ed878a070d4f6251['h00c1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00610] =  If409768b648a33a7ed878a070d4f6251['h00c20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00611] =  If409768b648a33a7ed878a070d4f6251['h00c22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00612] =  If409768b648a33a7ed878a070d4f6251['h00c24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00613] =  If409768b648a33a7ed878a070d4f6251['h00c26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00614] =  If409768b648a33a7ed878a070d4f6251['h00c28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00615] =  If409768b648a33a7ed878a070d4f6251['h00c2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00616] =  If409768b648a33a7ed878a070d4f6251['h00c2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00617] =  If409768b648a33a7ed878a070d4f6251['h00c2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00618] =  If409768b648a33a7ed878a070d4f6251['h00c30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00619] =  If409768b648a33a7ed878a070d4f6251['h00c32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0061a] =  If409768b648a33a7ed878a070d4f6251['h00c34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0061b] =  If409768b648a33a7ed878a070d4f6251['h00c36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0061c] =  If409768b648a33a7ed878a070d4f6251['h00c38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0061d] =  If409768b648a33a7ed878a070d4f6251['h00c3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0061e] =  If409768b648a33a7ed878a070d4f6251['h00c3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0061f] =  If409768b648a33a7ed878a070d4f6251['h00c3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00620] =  If409768b648a33a7ed878a070d4f6251['h00c40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00621] =  If409768b648a33a7ed878a070d4f6251['h00c42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00622] =  If409768b648a33a7ed878a070d4f6251['h00c44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00623] =  If409768b648a33a7ed878a070d4f6251['h00c46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00624] =  If409768b648a33a7ed878a070d4f6251['h00c48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00625] =  If409768b648a33a7ed878a070d4f6251['h00c4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00626] =  If409768b648a33a7ed878a070d4f6251['h00c4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00627] =  If409768b648a33a7ed878a070d4f6251['h00c4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00628] =  If409768b648a33a7ed878a070d4f6251['h00c50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00629] =  If409768b648a33a7ed878a070d4f6251['h00c52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0062a] =  If409768b648a33a7ed878a070d4f6251['h00c54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0062b] =  If409768b648a33a7ed878a070d4f6251['h00c56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0062c] =  If409768b648a33a7ed878a070d4f6251['h00c58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0062d] =  If409768b648a33a7ed878a070d4f6251['h00c5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0062e] =  If409768b648a33a7ed878a070d4f6251['h00c5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0062f] =  If409768b648a33a7ed878a070d4f6251['h00c5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00630] =  If409768b648a33a7ed878a070d4f6251['h00c60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00631] =  If409768b648a33a7ed878a070d4f6251['h00c62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00632] =  If409768b648a33a7ed878a070d4f6251['h00c64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00633] =  If409768b648a33a7ed878a070d4f6251['h00c66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00634] =  If409768b648a33a7ed878a070d4f6251['h00c68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00635] =  If409768b648a33a7ed878a070d4f6251['h00c6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00636] =  If409768b648a33a7ed878a070d4f6251['h00c6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00637] =  If409768b648a33a7ed878a070d4f6251['h00c6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00638] =  If409768b648a33a7ed878a070d4f6251['h00c70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00639] =  If409768b648a33a7ed878a070d4f6251['h00c72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0063a] =  If409768b648a33a7ed878a070d4f6251['h00c74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0063b] =  If409768b648a33a7ed878a070d4f6251['h00c76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0063c] =  If409768b648a33a7ed878a070d4f6251['h00c78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0063d] =  If409768b648a33a7ed878a070d4f6251['h00c7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0063e] =  If409768b648a33a7ed878a070d4f6251['h00c7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0063f] =  If409768b648a33a7ed878a070d4f6251['h00c7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00640] =  If409768b648a33a7ed878a070d4f6251['h00c80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00641] =  If409768b648a33a7ed878a070d4f6251['h00c82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00642] =  If409768b648a33a7ed878a070d4f6251['h00c84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00643] =  If409768b648a33a7ed878a070d4f6251['h00c86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00644] =  If409768b648a33a7ed878a070d4f6251['h00c88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00645] =  If409768b648a33a7ed878a070d4f6251['h00c8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00646] =  If409768b648a33a7ed878a070d4f6251['h00c8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00647] =  If409768b648a33a7ed878a070d4f6251['h00c8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00648] =  If409768b648a33a7ed878a070d4f6251['h00c90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00649] =  If409768b648a33a7ed878a070d4f6251['h00c92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0064a] =  If409768b648a33a7ed878a070d4f6251['h00c94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0064b] =  If409768b648a33a7ed878a070d4f6251['h00c96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0064c] =  If409768b648a33a7ed878a070d4f6251['h00c98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0064d] =  If409768b648a33a7ed878a070d4f6251['h00c9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0064e] =  If409768b648a33a7ed878a070d4f6251['h00c9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0064f] =  If409768b648a33a7ed878a070d4f6251['h00c9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00650] =  If409768b648a33a7ed878a070d4f6251['h00ca0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00651] =  If409768b648a33a7ed878a070d4f6251['h00ca2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00652] =  If409768b648a33a7ed878a070d4f6251['h00ca4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00653] =  If409768b648a33a7ed878a070d4f6251['h00ca6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00654] =  If409768b648a33a7ed878a070d4f6251['h00ca8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00655] =  If409768b648a33a7ed878a070d4f6251['h00caa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00656] =  If409768b648a33a7ed878a070d4f6251['h00cac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00657] =  If409768b648a33a7ed878a070d4f6251['h00cae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00658] =  If409768b648a33a7ed878a070d4f6251['h00cb0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00659] =  If409768b648a33a7ed878a070d4f6251['h00cb2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0065a] =  If409768b648a33a7ed878a070d4f6251['h00cb4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0065b] =  If409768b648a33a7ed878a070d4f6251['h00cb6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0065c] =  If409768b648a33a7ed878a070d4f6251['h00cb8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0065d] =  If409768b648a33a7ed878a070d4f6251['h00cba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0065e] =  If409768b648a33a7ed878a070d4f6251['h00cbc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0065f] =  If409768b648a33a7ed878a070d4f6251['h00cbe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00660] =  If409768b648a33a7ed878a070d4f6251['h00cc0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00661] =  If409768b648a33a7ed878a070d4f6251['h00cc2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00662] =  If409768b648a33a7ed878a070d4f6251['h00cc4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00663] =  If409768b648a33a7ed878a070d4f6251['h00cc6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00664] =  If409768b648a33a7ed878a070d4f6251['h00cc8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00665] =  If409768b648a33a7ed878a070d4f6251['h00cca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00666] =  If409768b648a33a7ed878a070d4f6251['h00ccc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00667] =  If409768b648a33a7ed878a070d4f6251['h00cce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00668] =  If409768b648a33a7ed878a070d4f6251['h00cd0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00669] =  If409768b648a33a7ed878a070d4f6251['h00cd2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0066a] =  If409768b648a33a7ed878a070d4f6251['h00cd4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0066b] =  If409768b648a33a7ed878a070d4f6251['h00cd6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0066c] =  If409768b648a33a7ed878a070d4f6251['h00cd8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0066d] =  If409768b648a33a7ed878a070d4f6251['h00cda] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0066e] =  If409768b648a33a7ed878a070d4f6251['h00cdc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0066f] =  If409768b648a33a7ed878a070d4f6251['h00cde] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00670] =  If409768b648a33a7ed878a070d4f6251['h00ce0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00671] =  If409768b648a33a7ed878a070d4f6251['h00ce2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00672] =  If409768b648a33a7ed878a070d4f6251['h00ce4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00673] =  If409768b648a33a7ed878a070d4f6251['h00ce6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00674] =  If409768b648a33a7ed878a070d4f6251['h00ce8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00675] =  If409768b648a33a7ed878a070d4f6251['h00cea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00676] =  If409768b648a33a7ed878a070d4f6251['h00cec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00677] =  If409768b648a33a7ed878a070d4f6251['h00cee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00678] =  If409768b648a33a7ed878a070d4f6251['h00cf0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00679] =  If409768b648a33a7ed878a070d4f6251['h00cf2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0067a] =  If409768b648a33a7ed878a070d4f6251['h00cf4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0067b] =  If409768b648a33a7ed878a070d4f6251['h00cf6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0067c] =  If409768b648a33a7ed878a070d4f6251['h00cf8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0067d] =  If409768b648a33a7ed878a070d4f6251['h00cfa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0067e] =  If409768b648a33a7ed878a070d4f6251['h00cfc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0067f] =  If409768b648a33a7ed878a070d4f6251['h00cfe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00680] =  If409768b648a33a7ed878a070d4f6251['h00d00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00681] =  If409768b648a33a7ed878a070d4f6251['h00d02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00682] =  If409768b648a33a7ed878a070d4f6251['h00d04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00683] =  If409768b648a33a7ed878a070d4f6251['h00d06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00684] =  If409768b648a33a7ed878a070d4f6251['h00d08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00685] =  If409768b648a33a7ed878a070d4f6251['h00d0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00686] =  If409768b648a33a7ed878a070d4f6251['h00d0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00687] =  If409768b648a33a7ed878a070d4f6251['h00d0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00688] =  If409768b648a33a7ed878a070d4f6251['h00d10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00689] =  If409768b648a33a7ed878a070d4f6251['h00d12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0068a] =  If409768b648a33a7ed878a070d4f6251['h00d14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0068b] =  If409768b648a33a7ed878a070d4f6251['h00d16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0068c] =  If409768b648a33a7ed878a070d4f6251['h00d18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0068d] =  If409768b648a33a7ed878a070d4f6251['h00d1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0068e] =  If409768b648a33a7ed878a070d4f6251['h00d1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0068f] =  If409768b648a33a7ed878a070d4f6251['h00d1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00690] =  If409768b648a33a7ed878a070d4f6251['h00d20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00691] =  If409768b648a33a7ed878a070d4f6251['h00d22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00692] =  If409768b648a33a7ed878a070d4f6251['h00d24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00693] =  If409768b648a33a7ed878a070d4f6251['h00d26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00694] =  If409768b648a33a7ed878a070d4f6251['h00d28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00695] =  If409768b648a33a7ed878a070d4f6251['h00d2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00696] =  If409768b648a33a7ed878a070d4f6251['h00d2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00697] =  If409768b648a33a7ed878a070d4f6251['h00d2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00698] =  If409768b648a33a7ed878a070d4f6251['h00d30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00699] =  If409768b648a33a7ed878a070d4f6251['h00d32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0069a] =  If409768b648a33a7ed878a070d4f6251['h00d34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0069b] =  If409768b648a33a7ed878a070d4f6251['h00d36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0069c] =  If409768b648a33a7ed878a070d4f6251['h00d38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0069d] =  If409768b648a33a7ed878a070d4f6251['h00d3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0069e] =  If409768b648a33a7ed878a070d4f6251['h00d3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0069f] =  If409768b648a33a7ed878a070d4f6251['h00d3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006a0] =  If409768b648a33a7ed878a070d4f6251['h00d40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006a1] =  If409768b648a33a7ed878a070d4f6251['h00d42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006a2] =  If409768b648a33a7ed878a070d4f6251['h00d44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006a3] =  If409768b648a33a7ed878a070d4f6251['h00d46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006a4] =  If409768b648a33a7ed878a070d4f6251['h00d48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006a5] =  If409768b648a33a7ed878a070d4f6251['h00d4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006a6] =  If409768b648a33a7ed878a070d4f6251['h00d4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006a7] =  If409768b648a33a7ed878a070d4f6251['h00d4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006a8] =  If409768b648a33a7ed878a070d4f6251['h00d50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006a9] =  If409768b648a33a7ed878a070d4f6251['h00d52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006aa] =  If409768b648a33a7ed878a070d4f6251['h00d54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ab] =  If409768b648a33a7ed878a070d4f6251['h00d56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ac] =  If409768b648a33a7ed878a070d4f6251['h00d58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ad] =  If409768b648a33a7ed878a070d4f6251['h00d5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ae] =  If409768b648a33a7ed878a070d4f6251['h00d5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006af] =  If409768b648a33a7ed878a070d4f6251['h00d5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006b0] =  If409768b648a33a7ed878a070d4f6251['h00d60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006b1] =  If409768b648a33a7ed878a070d4f6251['h00d62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006b2] =  If409768b648a33a7ed878a070d4f6251['h00d64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006b3] =  If409768b648a33a7ed878a070d4f6251['h00d66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006b4] =  If409768b648a33a7ed878a070d4f6251['h00d68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006b5] =  If409768b648a33a7ed878a070d4f6251['h00d6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006b6] =  If409768b648a33a7ed878a070d4f6251['h00d6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006b7] =  If409768b648a33a7ed878a070d4f6251['h00d6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006b8] =  If409768b648a33a7ed878a070d4f6251['h00d70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006b9] =  If409768b648a33a7ed878a070d4f6251['h00d72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ba] =  If409768b648a33a7ed878a070d4f6251['h00d74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006bb] =  If409768b648a33a7ed878a070d4f6251['h00d76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006bc] =  If409768b648a33a7ed878a070d4f6251['h00d78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006bd] =  If409768b648a33a7ed878a070d4f6251['h00d7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006be] =  If409768b648a33a7ed878a070d4f6251['h00d7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006bf] =  If409768b648a33a7ed878a070d4f6251['h00d7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006c0] =  If409768b648a33a7ed878a070d4f6251['h00d80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006c1] =  If409768b648a33a7ed878a070d4f6251['h00d82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006c2] =  If409768b648a33a7ed878a070d4f6251['h00d84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006c3] =  If409768b648a33a7ed878a070d4f6251['h00d86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006c4] =  If409768b648a33a7ed878a070d4f6251['h00d88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006c5] =  If409768b648a33a7ed878a070d4f6251['h00d8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006c6] =  If409768b648a33a7ed878a070d4f6251['h00d8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006c7] =  If409768b648a33a7ed878a070d4f6251['h00d8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006c8] =  If409768b648a33a7ed878a070d4f6251['h00d90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006c9] =  If409768b648a33a7ed878a070d4f6251['h00d92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ca] =  If409768b648a33a7ed878a070d4f6251['h00d94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006cb] =  If409768b648a33a7ed878a070d4f6251['h00d96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006cc] =  If409768b648a33a7ed878a070d4f6251['h00d98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006cd] =  If409768b648a33a7ed878a070d4f6251['h00d9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ce] =  If409768b648a33a7ed878a070d4f6251['h00d9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006cf] =  If409768b648a33a7ed878a070d4f6251['h00d9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006d0] =  If409768b648a33a7ed878a070d4f6251['h00da0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006d1] =  If409768b648a33a7ed878a070d4f6251['h00da2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006d2] =  If409768b648a33a7ed878a070d4f6251['h00da4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006d3] =  If409768b648a33a7ed878a070d4f6251['h00da6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006d4] =  If409768b648a33a7ed878a070d4f6251['h00da8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006d5] =  If409768b648a33a7ed878a070d4f6251['h00daa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006d6] =  If409768b648a33a7ed878a070d4f6251['h00dac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006d7] =  If409768b648a33a7ed878a070d4f6251['h00dae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006d8] =  If409768b648a33a7ed878a070d4f6251['h00db0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006d9] =  If409768b648a33a7ed878a070d4f6251['h00db2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006da] =  If409768b648a33a7ed878a070d4f6251['h00db4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006db] =  If409768b648a33a7ed878a070d4f6251['h00db6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006dc] =  If409768b648a33a7ed878a070d4f6251['h00db8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006dd] =  If409768b648a33a7ed878a070d4f6251['h00dba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006de] =  If409768b648a33a7ed878a070d4f6251['h00dbc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006df] =  If409768b648a33a7ed878a070d4f6251['h00dbe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006e0] =  If409768b648a33a7ed878a070d4f6251['h00dc0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006e1] =  If409768b648a33a7ed878a070d4f6251['h00dc2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006e2] =  If409768b648a33a7ed878a070d4f6251['h00dc4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006e3] =  If409768b648a33a7ed878a070d4f6251['h00dc6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006e4] =  If409768b648a33a7ed878a070d4f6251['h00dc8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006e5] =  If409768b648a33a7ed878a070d4f6251['h00dca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006e6] =  If409768b648a33a7ed878a070d4f6251['h00dcc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006e7] =  If409768b648a33a7ed878a070d4f6251['h00dce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006e8] =  If409768b648a33a7ed878a070d4f6251['h00dd0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006e9] =  If409768b648a33a7ed878a070d4f6251['h00dd2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ea] =  If409768b648a33a7ed878a070d4f6251['h00dd4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006eb] =  If409768b648a33a7ed878a070d4f6251['h00dd6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ec] =  If409768b648a33a7ed878a070d4f6251['h00dd8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ed] =  If409768b648a33a7ed878a070d4f6251['h00dda] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ee] =  If409768b648a33a7ed878a070d4f6251['h00ddc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ef] =  If409768b648a33a7ed878a070d4f6251['h00dde] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006f0] =  If409768b648a33a7ed878a070d4f6251['h00de0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006f1] =  If409768b648a33a7ed878a070d4f6251['h00de2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006f2] =  If409768b648a33a7ed878a070d4f6251['h00de4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006f3] =  If409768b648a33a7ed878a070d4f6251['h00de6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006f4] =  If409768b648a33a7ed878a070d4f6251['h00de8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006f5] =  If409768b648a33a7ed878a070d4f6251['h00dea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006f6] =  If409768b648a33a7ed878a070d4f6251['h00dec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006f7] =  If409768b648a33a7ed878a070d4f6251['h00dee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006f8] =  If409768b648a33a7ed878a070d4f6251['h00df0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006f9] =  If409768b648a33a7ed878a070d4f6251['h00df2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006fa] =  If409768b648a33a7ed878a070d4f6251['h00df4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006fb] =  If409768b648a33a7ed878a070d4f6251['h00df6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006fc] =  If409768b648a33a7ed878a070d4f6251['h00df8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006fd] =  If409768b648a33a7ed878a070d4f6251['h00dfa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006fe] =  If409768b648a33a7ed878a070d4f6251['h00dfc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h006ff] =  If409768b648a33a7ed878a070d4f6251['h00dfe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00700] =  If409768b648a33a7ed878a070d4f6251['h00e00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00701] =  If409768b648a33a7ed878a070d4f6251['h00e02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00702] =  If409768b648a33a7ed878a070d4f6251['h00e04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00703] =  If409768b648a33a7ed878a070d4f6251['h00e06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00704] =  If409768b648a33a7ed878a070d4f6251['h00e08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00705] =  If409768b648a33a7ed878a070d4f6251['h00e0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00706] =  If409768b648a33a7ed878a070d4f6251['h00e0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00707] =  If409768b648a33a7ed878a070d4f6251['h00e0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00708] =  If409768b648a33a7ed878a070d4f6251['h00e10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00709] =  If409768b648a33a7ed878a070d4f6251['h00e12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0070a] =  If409768b648a33a7ed878a070d4f6251['h00e14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0070b] =  If409768b648a33a7ed878a070d4f6251['h00e16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0070c] =  If409768b648a33a7ed878a070d4f6251['h00e18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0070d] =  If409768b648a33a7ed878a070d4f6251['h00e1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0070e] =  If409768b648a33a7ed878a070d4f6251['h00e1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0070f] =  If409768b648a33a7ed878a070d4f6251['h00e1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00710] =  If409768b648a33a7ed878a070d4f6251['h00e20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00711] =  If409768b648a33a7ed878a070d4f6251['h00e22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00712] =  If409768b648a33a7ed878a070d4f6251['h00e24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00713] =  If409768b648a33a7ed878a070d4f6251['h00e26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00714] =  If409768b648a33a7ed878a070d4f6251['h00e28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00715] =  If409768b648a33a7ed878a070d4f6251['h00e2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00716] =  If409768b648a33a7ed878a070d4f6251['h00e2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00717] =  If409768b648a33a7ed878a070d4f6251['h00e2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00718] =  If409768b648a33a7ed878a070d4f6251['h00e30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00719] =  If409768b648a33a7ed878a070d4f6251['h00e32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0071a] =  If409768b648a33a7ed878a070d4f6251['h00e34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0071b] =  If409768b648a33a7ed878a070d4f6251['h00e36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0071c] =  If409768b648a33a7ed878a070d4f6251['h00e38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0071d] =  If409768b648a33a7ed878a070d4f6251['h00e3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0071e] =  If409768b648a33a7ed878a070d4f6251['h00e3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0071f] =  If409768b648a33a7ed878a070d4f6251['h00e3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00720] =  If409768b648a33a7ed878a070d4f6251['h00e40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00721] =  If409768b648a33a7ed878a070d4f6251['h00e42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00722] =  If409768b648a33a7ed878a070d4f6251['h00e44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00723] =  If409768b648a33a7ed878a070d4f6251['h00e46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00724] =  If409768b648a33a7ed878a070d4f6251['h00e48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00725] =  If409768b648a33a7ed878a070d4f6251['h00e4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00726] =  If409768b648a33a7ed878a070d4f6251['h00e4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00727] =  If409768b648a33a7ed878a070d4f6251['h00e4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00728] =  If409768b648a33a7ed878a070d4f6251['h00e50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00729] =  If409768b648a33a7ed878a070d4f6251['h00e52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0072a] =  If409768b648a33a7ed878a070d4f6251['h00e54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0072b] =  If409768b648a33a7ed878a070d4f6251['h00e56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0072c] =  If409768b648a33a7ed878a070d4f6251['h00e58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0072d] =  If409768b648a33a7ed878a070d4f6251['h00e5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0072e] =  If409768b648a33a7ed878a070d4f6251['h00e5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0072f] =  If409768b648a33a7ed878a070d4f6251['h00e5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00730] =  If409768b648a33a7ed878a070d4f6251['h00e60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00731] =  If409768b648a33a7ed878a070d4f6251['h00e62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00732] =  If409768b648a33a7ed878a070d4f6251['h00e64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00733] =  If409768b648a33a7ed878a070d4f6251['h00e66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00734] =  If409768b648a33a7ed878a070d4f6251['h00e68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00735] =  If409768b648a33a7ed878a070d4f6251['h00e6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00736] =  If409768b648a33a7ed878a070d4f6251['h00e6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00737] =  If409768b648a33a7ed878a070d4f6251['h00e6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00738] =  If409768b648a33a7ed878a070d4f6251['h00e70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00739] =  If409768b648a33a7ed878a070d4f6251['h00e72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0073a] =  If409768b648a33a7ed878a070d4f6251['h00e74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0073b] =  If409768b648a33a7ed878a070d4f6251['h00e76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0073c] =  If409768b648a33a7ed878a070d4f6251['h00e78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0073d] =  If409768b648a33a7ed878a070d4f6251['h00e7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0073e] =  If409768b648a33a7ed878a070d4f6251['h00e7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0073f] =  If409768b648a33a7ed878a070d4f6251['h00e7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00740] =  If409768b648a33a7ed878a070d4f6251['h00e80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00741] =  If409768b648a33a7ed878a070d4f6251['h00e82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00742] =  If409768b648a33a7ed878a070d4f6251['h00e84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00743] =  If409768b648a33a7ed878a070d4f6251['h00e86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00744] =  If409768b648a33a7ed878a070d4f6251['h00e88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00745] =  If409768b648a33a7ed878a070d4f6251['h00e8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00746] =  If409768b648a33a7ed878a070d4f6251['h00e8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00747] =  If409768b648a33a7ed878a070d4f6251['h00e8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00748] =  If409768b648a33a7ed878a070d4f6251['h00e90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00749] =  If409768b648a33a7ed878a070d4f6251['h00e92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0074a] =  If409768b648a33a7ed878a070d4f6251['h00e94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0074b] =  If409768b648a33a7ed878a070d4f6251['h00e96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0074c] =  If409768b648a33a7ed878a070d4f6251['h00e98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0074d] =  If409768b648a33a7ed878a070d4f6251['h00e9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0074e] =  If409768b648a33a7ed878a070d4f6251['h00e9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0074f] =  If409768b648a33a7ed878a070d4f6251['h00e9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00750] =  If409768b648a33a7ed878a070d4f6251['h00ea0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00751] =  If409768b648a33a7ed878a070d4f6251['h00ea2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00752] =  If409768b648a33a7ed878a070d4f6251['h00ea4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00753] =  If409768b648a33a7ed878a070d4f6251['h00ea6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00754] =  If409768b648a33a7ed878a070d4f6251['h00ea8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00755] =  If409768b648a33a7ed878a070d4f6251['h00eaa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00756] =  If409768b648a33a7ed878a070d4f6251['h00eac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00757] =  If409768b648a33a7ed878a070d4f6251['h00eae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00758] =  If409768b648a33a7ed878a070d4f6251['h00eb0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00759] =  If409768b648a33a7ed878a070d4f6251['h00eb2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0075a] =  If409768b648a33a7ed878a070d4f6251['h00eb4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0075b] =  If409768b648a33a7ed878a070d4f6251['h00eb6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0075c] =  If409768b648a33a7ed878a070d4f6251['h00eb8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0075d] =  If409768b648a33a7ed878a070d4f6251['h00eba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0075e] =  If409768b648a33a7ed878a070d4f6251['h00ebc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0075f] =  If409768b648a33a7ed878a070d4f6251['h00ebe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00760] =  If409768b648a33a7ed878a070d4f6251['h00ec0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00761] =  If409768b648a33a7ed878a070d4f6251['h00ec2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00762] =  If409768b648a33a7ed878a070d4f6251['h00ec4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00763] =  If409768b648a33a7ed878a070d4f6251['h00ec6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00764] =  If409768b648a33a7ed878a070d4f6251['h00ec8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00765] =  If409768b648a33a7ed878a070d4f6251['h00eca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00766] =  If409768b648a33a7ed878a070d4f6251['h00ecc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00767] =  If409768b648a33a7ed878a070d4f6251['h00ece] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00768] =  If409768b648a33a7ed878a070d4f6251['h00ed0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00769] =  If409768b648a33a7ed878a070d4f6251['h00ed2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0076a] =  If409768b648a33a7ed878a070d4f6251['h00ed4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0076b] =  If409768b648a33a7ed878a070d4f6251['h00ed6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0076c] =  If409768b648a33a7ed878a070d4f6251['h00ed8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0076d] =  If409768b648a33a7ed878a070d4f6251['h00eda] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0076e] =  If409768b648a33a7ed878a070d4f6251['h00edc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0076f] =  If409768b648a33a7ed878a070d4f6251['h00ede] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00770] =  If409768b648a33a7ed878a070d4f6251['h00ee0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00771] =  If409768b648a33a7ed878a070d4f6251['h00ee2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00772] =  If409768b648a33a7ed878a070d4f6251['h00ee4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00773] =  If409768b648a33a7ed878a070d4f6251['h00ee6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00774] =  If409768b648a33a7ed878a070d4f6251['h00ee8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00775] =  If409768b648a33a7ed878a070d4f6251['h00eea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00776] =  If409768b648a33a7ed878a070d4f6251['h00eec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00777] =  If409768b648a33a7ed878a070d4f6251['h00eee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00778] =  If409768b648a33a7ed878a070d4f6251['h00ef0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00779] =  If409768b648a33a7ed878a070d4f6251['h00ef2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0077a] =  If409768b648a33a7ed878a070d4f6251['h00ef4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0077b] =  If409768b648a33a7ed878a070d4f6251['h00ef6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0077c] =  If409768b648a33a7ed878a070d4f6251['h00ef8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0077d] =  If409768b648a33a7ed878a070d4f6251['h00efa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0077e] =  If409768b648a33a7ed878a070d4f6251['h00efc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0077f] =  If409768b648a33a7ed878a070d4f6251['h00efe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00780] =  If409768b648a33a7ed878a070d4f6251['h00f00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00781] =  If409768b648a33a7ed878a070d4f6251['h00f02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00782] =  If409768b648a33a7ed878a070d4f6251['h00f04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00783] =  If409768b648a33a7ed878a070d4f6251['h00f06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00784] =  If409768b648a33a7ed878a070d4f6251['h00f08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00785] =  If409768b648a33a7ed878a070d4f6251['h00f0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00786] =  If409768b648a33a7ed878a070d4f6251['h00f0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00787] =  If409768b648a33a7ed878a070d4f6251['h00f0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00788] =  If409768b648a33a7ed878a070d4f6251['h00f10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00789] =  If409768b648a33a7ed878a070d4f6251['h00f12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0078a] =  If409768b648a33a7ed878a070d4f6251['h00f14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0078b] =  If409768b648a33a7ed878a070d4f6251['h00f16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0078c] =  If409768b648a33a7ed878a070d4f6251['h00f18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0078d] =  If409768b648a33a7ed878a070d4f6251['h00f1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0078e] =  If409768b648a33a7ed878a070d4f6251['h00f1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0078f] =  If409768b648a33a7ed878a070d4f6251['h00f1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00790] =  If409768b648a33a7ed878a070d4f6251['h00f20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00791] =  If409768b648a33a7ed878a070d4f6251['h00f22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00792] =  If409768b648a33a7ed878a070d4f6251['h00f24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00793] =  If409768b648a33a7ed878a070d4f6251['h00f26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00794] =  If409768b648a33a7ed878a070d4f6251['h00f28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00795] =  If409768b648a33a7ed878a070d4f6251['h00f2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00796] =  If409768b648a33a7ed878a070d4f6251['h00f2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00797] =  If409768b648a33a7ed878a070d4f6251['h00f2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00798] =  If409768b648a33a7ed878a070d4f6251['h00f30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00799] =  If409768b648a33a7ed878a070d4f6251['h00f32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0079a] =  If409768b648a33a7ed878a070d4f6251['h00f34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0079b] =  If409768b648a33a7ed878a070d4f6251['h00f36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0079c] =  If409768b648a33a7ed878a070d4f6251['h00f38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0079d] =  If409768b648a33a7ed878a070d4f6251['h00f3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0079e] =  If409768b648a33a7ed878a070d4f6251['h00f3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0079f] =  If409768b648a33a7ed878a070d4f6251['h00f3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007a0] =  If409768b648a33a7ed878a070d4f6251['h00f40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007a1] =  If409768b648a33a7ed878a070d4f6251['h00f42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007a2] =  If409768b648a33a7ed878a070d4f6251['h00f44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007a3] =  If409768b648a33a7ed878a070d4f6251['h00f46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007a4] =  If409768b648a33a7ed878a070d4f6251['h00f48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007a5] =  If409768b648a33a7ed878a070d4f6251['h00f4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007a6] =  If409768b648a33a7ed878a070d4f6251['h00f4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007a7] =  If409768b648a33a7ed878a070d4f6251['h00f4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007a8] =  If409768b648a33a7ed878a070d4f6251['h00f50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007a9] =  If409768b648a33a7ed878a070d4f6251['h00f52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007aa] =  If409768b648a33a7ed878a070d4f6251['h00f54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ab] =  If409768b648a33a7ed878a070d4f6251['h00f56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ac] =  If409768b648a33a7ed878a070d4f6251['h00f58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ad] =  If409768b648a33a7ed878a070d4f6251['h00f5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ae] =  If409768b648a33a7ed878a070d4f6251['h00f5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007af] =  If409768b648a33a7ed878a070d4f6251['h00f5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007b0] =  If409768b648a33a7ed878a070d4f6251['h00f60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007b1] =  If409768b648a33a7ed878a070d4f6251['h00f62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007b2] =  If409768b648a33a7ed878a070d4f6251['h00f64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007b3] =  If409768b648a33a7ed878a070d4f6251['h00f66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007b4] =  If409768b648a33a7ed878a070d4f6251['h00f68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007b5] =  If409768b648a33a7ed878a070d4f6251['h00f6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007b6] =  If409768b648a33a7ed878a070d4f6251['h00f6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007b7] =  If409768b648a33a7ed878a070d4f6251['h00f6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007b8] =  If409768b648a33a7ed878a070d4f6251['h00f70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007b9] =  If409768b648a33a7ed878a070d4f6251['h00f72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ba] =  If409768b648a33a7ed878a070d4f6251['h00f74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007bb] =  If409768b648a33a7ed878a070d4f6251['h00f76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007bc] =  If409768b648a33a7ed878a070d4f6251['h00f78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007bd] =  If409768b648a33a7ed878a070d4f6251['h00f7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007be] =  If409768b648a33a7ed878a070d4f6251['h00f7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007bf] =  If409768b648a33a7ed878a070d4f6251['h00f7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007c0] =  If409768b648a33a7ed878a070d4f6251['h00f80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007c1] =  If409768b648a33a7ed878a070d4f6251['h00f82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007c2] =  If409768b648a33a7ed878a070d4f6251['h00f84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007c3] =  If409768b648a33a7ed878a070d4f6251['h00f86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007c4] =  If409768b648a33a7ed878a070d4f6251['h00f88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007c5] =  If409768b648a33a7ed878a070d4f6251['h00f8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007c6] =  If409768b648a33a7ed878a070d4f6251['h00f8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007c7] =  If409768b648a33a7ed878a070d4f6251['h00f8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007c8] =  If409768b648a33a7ed878a070d4f6251['h00f90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007c9] =  If409768b648a33a7ed878a070d4f6251['h00f92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ca] =  If409768b648a33a7ed878a070d4f6251['h00f94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007cb] =  If409768b648a33a7ed878a070d4f6251['h00f96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007cc] =  If409768b648a33a7ed878a070d4f6251['h00f98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007cd] =  If409768b648a33a7ed878a070d4f6251['h00f9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ce] =  If409768b648a33a7ed878a070d4f6251['h00f9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007cf] =  If409768b648a33a7ed878a070d4f6251['h00f9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007d0] =  If409768b648a33a7ed878a070d4f6251['h00fa0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007d1] =  If409768b648a33a7ed878a070d4f6251['h00fa2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007d2] =  If409768b648a33a7ed878a070d4f6251['h00fa4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007d3] =  If409768b648a33a7ed878a070d4f6251['h00fa6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007d4] =  If409768b648a33a7ed878a070d4f6251['h00fa8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007d5] =  If409768b648a33a7ed878a070d4f6251['h00faa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007d6] =  If409768b648a33a7ed878a070d4f6251['h00fac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007d7] =  If409768b648a33a7ed878a070d4f6251['h00fae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007d8] =  If409768b648a33a7ed878a070d4f6251['h00fb0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007d9] =  If409768b648a33a7ed878a070d4f6251['h00fb2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007da] =  If409768b648a33a7ed878a070d4f6251['h00fb4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007db] =  If409768b648a33a7ed878a070d4f6251['h00fb6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007dc] =  If409768b648a33a7ed878a070d4f6251['h00fb8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007dd] =  If409768b648a33a7ed878a070d4f6251['h00fba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007de] =  If409768b648a33a7ed878a070d4f6251['h00fbc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007df] =  If409768b648a33a7ed878a070d4f6251['h00fbe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007e0] =  If409768b648a33a7ed878a070d4f6251['h00fc0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007e1] =  If409768b648a33a7ed878a070d4f6251['h00fc2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007e2] =  If409768b648a33a7ed878a070d4f6251['h00fc4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007e3] =  If409768b648a33a7ed878a070d4f6251['h00fc6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007e4] =  If409768b648a33a7ed878a070d4f6251['h00fc8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007e5] =  If409768b648a33a7ed878a070d4f6251['h00fca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007e6] =  If409768b648a33a7ed878a070d4f6251['h00fcc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007e7] =  If409768b648a33a7ed878a070d4f6251['h00fce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007e8] =  If409768b648a33a7ed878a070d4f6251['h00fd0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007e9] =  If409768b648a33a7ed878a070d4f6251['h00fd2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ea] =  If409768b648a33a7ed878a070d4f6251['h00fd4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007eb] =  If409768b648a33a7ed878a070d4f6251['h00fd6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ec] =  If409768b648a33a7ed878a070d4f6251['h00fd8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ed] =  If409768b648a33a7ed878a070d4f6251['h00fda] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ee] =  If409768b648a33a7ed878a070d4f6251['h00fdc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ef] =  If409768b648a33a7ed878a070d4f6251['h00fde] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007f0] =  If409768b648a33a7ed878a070d4f6251['h00fe0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007f1] =  If409768b648a33a7ed878a070d4f6251['h00fe2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007f2] =  If409768b648a33a7ed878a070d4f6251['h00fe4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007f3] =  If409768b648a33a7ed878a070d4f6251['h00fe6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007f4] =  If409768b648a33a7ed878a070d4f6251['h00fe8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007f5] =  If409768b648a33a7ed878a070d4f6251['h00fea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007f6] =  If409768b648a33a7ed878a070d4f6251['h00fec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007f7] =  If409768b648a33a7ed878a070d4f6251['h00fee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007f8] =  If409768b648a33a7ed878a070d4f6251['h00ff0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007f9] =  If409768b648a33a7ed878a070d4f6251['h00ff2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007fa] =  If409768b648a33a7ed878a070d4f6251['h00ff4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007fb] =  If409768b648a33a7ed878a070d4f6251['h00ff6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007fc] =  If409768b648a33a7ed878a070d4f6251['h00ff8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007fd] =  If409768b648a33a7ed878a070d4f6251['h00ffa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007fe] =  If409768b648a33a7ed878a070d4f6251['h00ffc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h007ff] =  If409768b648a33a7ed878a070d4f6251['h00ffe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00800] =  If409768b648a33a7ed878a070d4f6251['h01000] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00801] =  If409768b648a33a7ed878a070d4f6251['h01002] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00802] =  If409768b648a33a7ed878a070d4f6251['h01004] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00803] =  If409768b648a33a7ed878a070d4f6251['h01006] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00804] =  If409768b648a33a7ed878a070d4f6251['h01008] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00805] =  If409768b648a33a7ed878a070d4f6251['h0100a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00806] =  If409768b648a33a7ed878a070d4f6251['h0100c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00807] =  If409768b648a33a7ed878a070d4f6251['h0100e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00808] =  If409768b648a33a7ed878a070d4f6251['h01010] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00809] =  If409768b648a33a7ed878a070d4f6251['h01012] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0080a] =  If409768b648a33a7ed878a070d4f6251['h01014] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0080b] =  If409768b648a33a7ed878a070d4f6251['h01016] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0080c] =  If409768b648a33a7ed878a070d4f6251['h01018] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0080d] =  If409768b648a33a7ed878a070d4f6251['h0101a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0080e] =  If409768b648a33a7ed878a070d4f6251['h0101c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0080f] =  If409768b648a33a7ed878a070d4f6251['h0101e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00810] =  If409768b648a33a7ed878a070d4f6251['h01020] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00811] =  If409768b648a33a7ed878a070d4f6251['h01022] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00812] =  If409768b648a33a7ed878a070d4f6251['h01024] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00813] =  If409768b648a33a7ed878a070d4f6251['h01026] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00814] =  If409768b648a33a7ed878a070d4f6251['h01028] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00815] =  If409768b648a33a7ed878a070d4f6251['h0102a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00816] =  If409768b648a33a7ed878a070d4f6251['h0102c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00817] =  If409768b648a33a7ed878a070d4f6251['h0102e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00818] =  If409768b648a33a7ed878a070d4f6251['h01030] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00819] =  If409768b648a33a7ed878a070d4f6251['h01032] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0081a] =  If409768b648a33a7ed878a070d4f6251['h01034] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0081b] =  If409768b648a33a7ed878a070d4f6251['h01036] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0081c] =  If409768b648a33a7ed878a070d4f6251['h01038] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0081d] =  If409768b648a33a7ed878a070d4f6251['h0103a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0081e] =  If409768b648a33a7ed878a070d4f6251['h0103c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0081f] =  If409768b648a33a7ed878a070d4f6251['h0103e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00820] =  If409768b648a33a7ed878a070d4f6251['h01040] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00821] =  If409768b648a33a7ed878a070d4f6251['h01042] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00822] =  If409768b648a33a7ed878a070d4f6251['h01044] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00823] =  If409768b648a33a7ed878a070d4f6251['h01046] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00824] =  If409768b648a33a7ed878a070d4f6251['h01048] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00825] =  If409768b648a33a7ed878a070d4f6251['h0104a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00826] =  If409768b648a33a7ed878a070d4f6251['h0104c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00827] =  If409768b648a33a7ed878a070d4f6251['h0104e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00828] =  If409768b648a33a7ed878a070d4f6251['h01050] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00829] =  If409768b648a33a7ed878a070d4f6251['h01052] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0082a] =  If409768b648a33a7ed878a070d4f6251['h01054] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0082b] =  If409768b648a33a7ed878a070d4f6251['h01056] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0082c] =  If409768b648a33a7ed878a070d4f6251['h01058] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0082d] =  If409768b648a33a7ed878a070d4f6251['h0105a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0082e] =  If409768b648a33a7ed878a070d4f6251['h0105c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0082f] =  If409768b648a33a7ed878a070d4f6251['h0105e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00830] =  If409768b648a33a7ed878a070d4f6251['h01060] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00831] =  If409768b648a33a7ed878a070d4f6251['h01062] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00832] =  If409768b648a33a7ed878a070d4f6251['h01064] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00833] =  If409768b648a33a7ed878a070d4f6251['h01066] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00834] =  If409768b648a33a7ed878a070d4f6251['h01068] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00835] =  If409768b648a33a7ed878a070d4f6251['h0106a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00836] =  If409768b648a33a7ed878a070d4f6251['h0106c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00837] =  If409768b648a33a7ed878a070d4f6251['h0106e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00838] =  If409768b648a33a7ed878a070d4f6251['h01070] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00839] =  If409768b648a33a7ed878a070d4f6251['h01072] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0083a] =  If409768b648a33a7ed878a070d4f6251['h01074] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0083b] =  If409768b648a33a7ed878a070d4f6251['h01076] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0083c] =  If409768b648a33a7ed878a070d4f6251['h01078] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0083d] =  If409768b648a33a7ed878a070d4f6251['h0107a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0083e] =  If409768b648a33a7ed878a070d4f6251['h0107c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0083f] =  If409768b648a33a7ed878a070d4f6251['h0107e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00840] =  If409768b648a33a7ed878a070d4f6251['h01080] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00841] =  If409768b648a33a7ed878a070d4f6251['h01082] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00842] =  If409768b648a33a7ed878a070d4f6251['h01084] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00843] =  If409768b648a33a7ed878a070d4f6251['h01086] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00844] =  If409768b648a33a7ed878a070d4f6251['h01088] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00845] =  If409768b648a33a7ed878a070d4f6251['h0108a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00846] =  If409768b648a33a7ed878a070d4f6251['h0108c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00847] =  If409768b648a33a7ed878a070d4f6251['h0108e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00848] =  If409768b648a33a7ed878a070d4f6251['h01090] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00849] =  If409768b648a33a7ed878a070d4f6251['h01092] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0084a] =  If409768b648a33a7ed878a070d4f6251['h01094] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0084b] =  If409768b648a33a7ed878a070d4f6251['h01096] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0084c] =  If409768b648a33a7ed878a070d4f6251['h01098] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0084d] =  If409768b648a33a7ed878a070d4f6251['h0109a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0084e] =  If409768b648a33a7ed878a070d4f6251['h0109c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0084f] =  If409768b648a33a7ed878a070d4f6251['h0109e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00850] =  If409768b648a33a7ed878a070d4f6251['h010a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00851] =  If409768b648a33a7ed878a070d4f6251['h010a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00852] =  If409768b648a33a7ed878a070d4f6251['h010a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00853] =  If409768b648a33a7ed878a070d4f6251['h010a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00854] =  If409768b648a33a7ed878a070d4f6251['h010a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00855] =  If409768b648a33a7ed878a070d4f6251['h010aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00856] =  If409768b648a33a7ed878a070d4f6251['h010ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00857] =  If409768b648a33a7ed878a070d4f6251['h010ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00858] =  If409768b648a33a7ed878a070d4f6251['h010b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00859] =  If409768b648a33a7ed878a070d4f6251['h010b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0085a] =  If409768b648a33a7ed878a070d4f6251['h010b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0085b] =  If409768b648a33a7ed878a070d4f6251['h010b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0085c] =  If409768b648a33a7ed878a070d4f6251['h010b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0085d] =  If409768b648a33a7ed878a070d4f6251['h010ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0085e] =  If409768b648a33a7ed878a070d4f6251['h010bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0085f] =  If409768b648a33a7ed878a070d4f6251['h010be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00860] =  If409768b648a33a7ed878a070d4f6251['h010c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00861] =  If409768b648a33a7ed878a070d4f6251['h010c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00862] =  If409768b648a33a7ed878a070d4f6251['h010c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00863] =  If409768b648a33a7ed878a070d4f6251['h010c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00864] =  If409768b648a33a7ed878a070d4f6251['h010c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00865] =  If409768b648a33a7ed878a070d4f6251['h010ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00866] =  If409768b648a33a7ed878a070d4f6251['h010cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00867] =  If409768b648a33a7ed878a070d4f6251['h010ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00868] =  If409768b648a33a7ed878a070d4f6251['h010d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00869] =  If409768b648a33a7ed878a070d4f6251['h010d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0086a] =  If409768b648a33a7ed878a070d4f6251['h010d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0086b] =  If409768b648a33a7ed878a070d4f6251['h010d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0086c] =  If409768b648a33a7ed878a070d4f6251['h010d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0086d] =  If409768b648a33a7ed878a070d4f6251['h010da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0086e] =  If409768b648a33a7ed878a070d4f6251['h010dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0086f] =  If409768b648a33a7ed878a070d4f6251['h010de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00870] =  If409768b648a33a7ed878a070d4f6251['h010e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00871] =  If409768b648a33a7ed878a070d4f6251['h010e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00872] =  If409768b648a33a7ed878a070d4f6251['h010e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00873] =  If409768b648a33a7ed878a070d4f6251['h010e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00874] =  If409768b648a33a7ed878a070d4f6251['h010e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00875] =  If409768b648a33a7ed878a070d4f6251['h010ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00876] =  If409768b648a33a7ed878a070d4f6251['h010ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00877] =  If409768b648a33a7ed878a070d4f6251['h010ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00878] =  If409768b648a33a7ed878a070d4f6251['h010f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00879] =  If409768b648a33a7ed878a070d4f6251['h010f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0087a] =  If409768b648a33a7ed878a070d4f6251['h010f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0087b] =  If409768b648a33a7ed878a070d4f6251['h010f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0087c] =  If409768b648a33a7ed878a070d4f6251['h010f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0087d] =  If409768b648a33a7ed878a070d4f6251['h010fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0087e] =  If409768b648a33a7ed878a070d4f6251['h010fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0087f] =  If409768b648a33a7ed878a070d4f6251['h010fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00880] =  If409768b648a33a7ed878a070d4f6251['h01100] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00881] =  If409768b648a33a7ed878a070d4f6251['h01102] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00882] =  If409768b648a33a7ed878a070d4f6251['h01104] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00883] =  If409768b648a33a7ed878a070d4f6251['h01106] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00884] =  If409768b648a33a7ed878a070d4f6251['h01108] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00885] =  If409768b648a33a7ed878a070d4f6251['h0110a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00886] =  If409768b648a33a7ed878a070d4f6251['h0110c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00887] =  If409768b648a33a7ed878a070d4f6251['h0110e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00888] =  If409768b648a33a7ed878a070d4f6251['h01110] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00889] =  If409768b648a33a7ed878a070d4f6251['h01112] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0088a] =  If409768b648a33a7ed878a070d4f6251['h01114] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0088b] =  If409768b648a33a7ed878a070d4f6251['h01116] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0088c] =  If409768b648a33a7ed878a070d4f6251['h01118] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0088d] =  If409768b648a33a7ed878a070d4f6251['h0111a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0088e] =  If409768b648a33a7ed878a070d4f6251['h0111c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0088f] =  If409768b648a33a7ed878a070d4f6251['h0111e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00890] =  If409768b648a33a7ed878a070d4f6251['h01120] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00891] =  If409768b648a33a7ed878a070d4f6251['h01122] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00892] =  If409768b648a33a7ed878a070d4f6251['h01124] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00893] =  If409768b648a33a7ed878a070d4f6251['h01126] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00894] =  If409768b648a33a7ed878a070d4f6251['h01128] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00895] =  If409768b648a33a7ed878a070d4f6251['h0112a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00896] =  If409768b648a33a7ed878a070d4f6251['h0112c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00897] =  If409768b648a33a7ed878a070d4f6251['h0112e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00898] =  If409768b648a33a7ed878a070d4f6251['h01130] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00899] =  If409768b648a33a7ed878a070d4f6251['h01132] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0089a] =  If409768b648a33a7ed878a070d4f6251['h01134] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0089b] =  If409768b648a33a7ed878a070d4f6251['h01136] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0089c] =  If409768b648a33a7ed878a070d4f6251['h01138] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0089d] =  If409768b648a33a7ed878a070d4f6251['h0113a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0089e] =  If409768b648a33a7ed878a070d4f6251['h0113c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0089f] =  If409768b648a33a7ed878a070d4f6251['h0113e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008a0] =  If409768b648a33a7ed878a070d4f6251['h01140] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008a1] =  If409768b648a33a7ed878a070d4f6251['h01142] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008a2] =  If409768b648a33a7ed878a070d4f6251['h01144] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008a3] =  If409768b648a33a7ed878a070d4f6251['h01146] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008a4] =  If409768b648a33a7ed878a070d4f6251['h01148] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008a5] =  If409768b648a33a7ed878a070d4f6251['h0114a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008a6] =  If409768b648a33a7ed878a070d4f6251['h0114c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008a7] =  If409768b648a33a7ed878a070d4f6251['h0114e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008a8] =  If409768b648a33a7ed878a070d4f6251['h01150] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008a9] =  If409768b648a33a7ed878a070d4f6251['h01152] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008aa] =  If409768b648a33a7ed878a070d4f6251['h01154] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ab] =  If409768b648a33a7ed878a070d4f6251['h01156] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ac] =  If409768b648a33a7ed878a070d4f6251['h01158] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ad] =  If409768b648a33a7ed878a070d4f6251['h0115a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ae] =  If409768b648a33a7ed878a070d4f6251['h0115c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008af] =  If409768b648a33a7ed878a070d4f6251['h0115e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008b0] =  If409768b648a33a7ed878a070d4f6251['h01160] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008b1] =  If409768b648a33a7ed878a070d4f6251['h01162] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008b2] =  If409768b648a33a7ed878a070d4f6251['h01164] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008b3] =  If409768b648a33a7ed878a070d4f6251['h01166] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008b4] =  If409768b648a33a7ed878a070d4f6251['h01168] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008b5] =  If409768b648a33a7ed878a070d4f6251['h0116a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008b6] =  If409768b648a33a7ed878a070d4f6251['h0116c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008b7] =  If409768b648a33a7ed878a070d4f6251['h0116e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008b8] =  If409768b648a33a7ed878a070d4f6251['h01170] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008b9] =  If409768b648a33a7ed878a070d4f6251['h01172] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ba] =  If409768b648a33a7ed878a070d4f6251['h01174] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008bb] =  If409768b648a33a7ed878a070d4f6251['h01176] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008bc] =  If409768b648a33a7ed878a070d4f6251['h01178] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008bd] =  If409768b648a33a7ed878a070d4f6251['h0117a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008be] =  If409768b648a33a7ed878a070d4f6251['h0117c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008bf] =  If409768b648a33a7ed878a070d4f6251['h0117e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008c0] =  If409768b648a33a7ed878a070d4f6251['h01180] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008c1] =  If409768b648a33a7ed878a070d4f6251['h01182] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008c2] =  If409768b648a33a7ed878a070d4f6251['h01184] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008c3] =  If409768b648a33a7ed878a070d4f6251['h01186] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008c4] =  If409768b648a33a7ed878a070d4f6251['h01188] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008c5] =  If409768b648a33a7ed878a070d4f6251['h0118a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008c6] =  If409768b648a33a7ed878a070d4f6251['h0118c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008c7] =  If409768b648a33a7ed878a070d4f6251['h0118e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008c8] =  If409768b648a33a7ed878a070d4f6251['h01190] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008c9] =  If409768b648a33a7ed878a070d4f6251['h01192] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ca] =  If409768b648a33a7ed878a070d4f6251['h01194] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008cb] =  If409768b648a33a7ed878a070d4f6251['h01196] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008cc] =  If409768b648a33a7ed878a070d4f6251['h01198] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008cd] =  If409768b648a33a7ed878a070d4f6251['h0119a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ce] =  If409768b648a33a7ed878a070d4f6251['h0119c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008cf] =  If409768b648a33a7ed878a070d4f6251['h0119e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008d0] =  If409768b648a33a7ed878a070d4f6251['h011a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008d1] =  If409768b648a33a7ed878a070d4f6251['h011a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008d2] =  If409768b648a33a7ed878a070d4f6251['h011a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008d3] =  If409768b648a33a7ed878a070d4f6251['h011a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008d4] =  If409768b648a33a7ed878a070d4f6251['h011a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008d5] =  If409768b648a33a7ed878a070d4f6251['h011aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008d6] =  If409768b648a33a7ed878a070d4f6251['h011ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008d7] =  If409768b648a33a7ed878a070d4f6251['h011ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008d8] =  If409768b648a33a7ed878a070d4f6251['h011b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008d9] =  If409768b648a33a7ed878a070d4f6251['h011b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008da] =  If409768b648a33a7ed878a070d4f6251['h011b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008db] =  If409768b648a33a7ed878a070d4f6251['h011b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008dc] =  If409768b648a33a7ed878a070d4f6251['h011b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008dd] =  If409768b648a33a7ed878a070d4f6251['h011ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008de] =  If409768b648a33a7ed878a070d4f6251['h011bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008df] =  If409768b648a33a7ed878a070d4f6251['h011be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008e0] =  If409768b648a33a7ed878a070d4f6251['h011c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008e1] =  If409768b648a33a7ed878a070d4f6251['h011c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008e2] =  If409768b648a33a7ed878a070d4f6251['h011c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008e3] =  If409768b648a33a7ed878a070d4f6251['h011c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008e4] =  If409768b648a33a7ed878a070d4f6251['h011c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008e5] =  If409768b648a33a7ed878a070d4f6251['h011ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008e6] =  If409768b648a33a7ed878a070d4f6251['h011cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008e7] =  If409768b648a33a7ed878a070d4f6251['h011ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008e8] =  If409768b648a33a7ed878a070d4f6251['h011d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008e9] =  If409768b648a33a7ed878a070d4f6251['h011d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ea] =  If409768b648a33a7ed878a070d4f6251['h011d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008eb] =  If409768b648a33a7ed878a070d4f6251['h011d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ec] =  If409768b648a33a7ed878a070d4f6251['h011d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ed] =  If409768b648a33a7ed878a070d4f6251['h011da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ee] =  If409768b648a33a7ed878a070d4f6251['h011dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ef] =  If409768b648a33a7ed878a070d4f6251['h011de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008f0] =  If409768b648a33a7ed878a070d4f6251['h011e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008f1] =  If409768b648a33a7ed878a070d4f6251['h011e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008f2] =  If409768b648a33a7ed878a070d4f6251['h011e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008f3] =  If409768b648a33a7ed878a070d4f6251['h011e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008f4] =  If409768b648a33a7ed878a070d4f6251['h011e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008f5] =  If409768b648a33a7ed878a070d4f6251['h011ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008f6] =  If409768b648a33a7ed878a070d4f6251['h011ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008f7] =  If409768b648a33a7ed878a070d4f6251['h011ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008f8] =  If409768b648a33a7ed878a070d4f6251['h011f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008f9] =  If409768b648a33a7ed878a070d4f6251['h011f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008fa] =  If409768b648a33a7ed878a070d4f6251['h011f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008fb] =  If409768b648a33a7ed878a070d4f6251['h011f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008fc] =  If409768b648a33a7ed878a070d4f6251['h011f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008fd] =  If409768b648a33a7ed878a070d4f6251['h011fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008fe] =  If409768b648a33a7ed878a070d4f6251['h011fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h008ff] =  If409768b648a33a7ed878a070d4f6251['h011fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00900] =  If409768b648a33a7ed878a070d4f6251['h01200] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00901] =  If409768b648a33a7ed878a070d4f6251['h01202] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00902] =  If409768b648a33a7ed878a070d4f6251['h01204] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00903] =  If409768b648a33a7ed878a070d4f6251['h01206] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00904] =  If409768b648a33a7ed878a070d4f6251['h01208] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00905] =  If409768b648a33a7ed878a070d4f6251['h0120a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00906] =  If409768b648a33a7ed878a070d4f6251['h0120c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00907] =  If409768b648a33a7ed878a070d4f6251['h0120e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00908] =  If409768b648a33a7ed878a070d4f6251['h01210] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00909] =  If409768b648a33a7ed878a070d4f6251['h01212] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0090a] =  If409768b648a33a7ed878a070d4f6251['h01214] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0090b] =  If409768b648a33a7ed878a070d4f6251['h01216] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0090c] =  If409768b648a33a7ed878a070d4f6251['h01218] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0090d] =  If409768b648a33a7ed878a070d4f6251['h0121a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0090e] =  If409768b648a33a7ed878a070d4f6251['h0121c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0090f] =  If409768b648a33a7ed878a070d4f6251['h0121e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00910] =  If409768b648a33a7ed878a070d4f6251['h01220] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00911] =  If409768b648a33a7ed878a070d4f6251['h01222] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00912] =  If409768b648a33a7ed878a070d4f6251['h01224] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00913] =  If409768b648a33a7ed878a070d4f6251['h01226] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00914] =  If409768b648a33a7ed878a070d4f6251['h01228] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00915] =  If409768b648a33a7ed878a070d4f6251['h0122a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00916] =  If409768b648a33a7ed878a070d4f6251['h0122c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00917] =  If409768b648a33a7ed878a070d4f6251['h0122e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00918] =  If409768b648a33a7ed878a070d4f6251['h01230] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00919] =  If409768b648a33a7ed878a070d4f6251['h01232] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0091a] =  If409768b648a33a7ed878a070d4f6251['h01234] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0091b] =  If409768b648a33a7ed878a070d4f6251['h01236] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0091c] =  If409768b648a33a7ed878a070d4f6251['h01238] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0091d] =  If409768b648a33a7ed878a070d4f6251['h0123a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0091e] =  If409768b648a33a7ed878a070d4f6251['h0123c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0091f] =  If409768b648a33a7ed878a070d4f6251['h0123e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00920] =  If409768b648a33a7ed878a070d4f6251['h01240] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00921] =  If409768b648a33a7ed878a070d4f6251['h01242] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00922] =  If409768b648a33a7ed878a070d4f6251['h01244] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00923] =  If409768b648a33a7ed878a070d4f6251['h01246] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00924] =  If409768b648a33a7ed878a070d4f6251['h01248] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00925] =  If409768b648a33a7ed878a070d4f6251['h0124a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00926] =  If409768b648a33a7ed878a070d4f6251['h0124c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00927] =  If409768b648a33a7ed878a070d4f6251['h0124e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00928] =  If409768b648a33a7ed878a070d4f6251['h01250] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00929] =  If409768b648a33a7ed878a070d4f6251['h01252] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0092a] =  If409768b648a33a7ed878a070d4f6251['h01254] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0092b] =  If409768b648a33a7ed878a070d4f6251['h01256] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0092c] =  If409768b648a33a7ed878a070d4f6251['h01258] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0092d] =  If409768b648a33a7ed878a070d4f6251['h0125a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0092e] =  If409768b648a33a7ed878a070d4f6251['h0125c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0092f] =  If409768b648a33a7ed878a070d4f6251['h0125e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00930] =  If409768b648a33a7ed878a070d4f6251['h01260] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00931] =  If409768b648a33a7ed878a070d4f6251['h01262] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00932] =  If409768b648a33a7ed878a070d4f6251['h01264] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00933] =  If409768b648a33a7ed878a070d4f6251['h01266] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00934] =  If409768b648a33a7ed878a070d4f6251['h01268] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00935] =  If409768b648a33a7ed878a070d4f6251['h0126a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00936] =  If409768b648a33a7ed878a070d4f6251['h0126c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00937] =  If409768b648a33a7ed878a070d4f6251['h0126e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00938] =  If409768b648a33a7ed878a070d4f6251['h01270] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00939] =  If409768b648a33a7ed878a070d4f6251['h01272] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0093a] =  If409768b648a33a7ed878a070d4f6251['h01274] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0093b] =  If409768b648a33a7ed878a070d4f6251['h01276] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0093c] =  If409768b648a33a7ed878a070d4f6251['h01278] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0093d] =  If409768b648a33a7ed878a070d4f6251['h0127a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0093e] =  If409768b648a33a7ed878a070d4f6251['h0127c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0093f] =  If409768b648a33a7ed878a070d4f6251['h0127e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00940] =  If409768b648a33a7ed878a070d4f6251['h01280] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00941] =  If409768b648a33a7ed878a070d4f6251['h01282] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00942] =  If409768b648a33a7ed878a070d4f6251['h01284] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00943] =  If409768b648a33a7ed878a070d4f6251['h01286] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00944] =  If409768b648a33a7ed878a070d4f6251['h01288] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00945] =  If409768b648a33a7ed878a070d4f6251['h0128a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00946] =  If409768b648a33a7ed878a070d4f6251['h0128c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00947] =  If409768b648a33a7ed878a070d4f6251['h0128e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00948] =  If409768b648a33a7ed878a070d4f6251['h01290] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00949] =  If409768b648a33a7ed878a070d4f6251['h01292] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0094a] =  If409768b648a33a7ed878a070d4f6251['h01294] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0094b] =  If409768b648a33a7ed878a070d4f6251['h01296] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0094c] =  If409768b648a33a7ed878a070d4f6251['h01298] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0094d] =  If409768b648a33a7ed878a070d4f6251['h0129a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0094e] =  If409768b648a33a7ed878a070d4f6251['h0129c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0094f] =  If409768b648a33a7ed878a070d4f6251['h0129e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00950] =  If409768b648a33a7ed878a070d4f6251['h012a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00951] =  If409768b648a33a7ed878a070d4f6251['h012a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00952] =  If409768b648a33a7ed878a070d4f6251['h012a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00953] =  If409768b648a33a7ed878a070d4f6251['h012a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00954] =  If409768b648a33a7ed878a070d4f6251['h012a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00955] =  If409768b648a33a7ed878a070d4f6251['h012aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00956] =  If409768b648a33a7ed878a070d4f6251['h012ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00957] =  If409768b648a33a7ed878a070d4f6251['h012ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00958] =  If409768b648a33a7ed878a070d4f6251['h012b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00959] =  If409768b648a33a7ed878a070d4f6251['h012b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0095a] =  If409768b648a33a7ed878a070d4f6251['h012b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0095b] =  If409768b648a33a7ed878a070d4f6251['h012b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0095c] =  If409768b648a33a7ed878a070d4f6251['h012b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0095d] =  If409768b648a33a7ed878a070d4f6251['h012ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0095e] =  If409768b648a33a7ed878a070d4f6251['h012bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0095f] =  If409768b648a33a7ed878a070d4f6251['h012be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00960] =  If409768b648a33a7ed878a070d4f6251['h012c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00961] =  If409768b648a33a7ed878a070d4f6251['h012c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00962] =  If409768b648a33a7ed878a070d4f6251['h012c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00963] =  If409768b648a33a7ed878a070d4f6251['h012c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00964] =  If409768b648a33a7ed878a070d4f6251['h012c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00965] =  If409768b648a33a7ed878a070d4f6251['h012ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00966] =  If409768b648a33a7ed878a070d4f6251['h012cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00967] =  If409768b648a33a7ed878a070d4f6251['h012ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00968] =  If409768b648a33a7ed878a070d4f6251['h012d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00969] =  If409768b648a33a7ed878a070d4f6251['h012d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0096a] =  If409768b648a33a7ed878a070d4f6251['h012d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0096b] =  If409768b648a33a7ed878a070d4f6251['h012d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0096c] =  If409768b648a33a7ed878a070d4f6251['h012d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0096d] =  If409768b648a33a7ed878a070d4f6251['h012da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0096e] =  If409768b648a33a7ed878a070d4f6251['h012dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0096f] =  If409768b648a33a7ed878a070d4f6251['h012de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00970] =  If409768b648a33a7ed878a070d4f6251['h012e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00971] =  If409768b648a33a7ed878a070d4f6251['h012e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00972] =  If409768b648a33a7ed878a070d4f6251['h012e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00973] =  If409768b648a33a7ed878a070d4f6251['h012e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00974] =  If409768b648a33a7ed878a070d4f6251['h012e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00975] =  If409768b648a33a7ed878a070d4f6251['h012ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00976] =  If409768b648a33a7ed878a070d4f6251['h012ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00977] =  If409768b648a33a7ed878a070d4f6251['h012ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00978] =  If409768b648a33a7ed878a070d4f6251['h012f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00979] =  If409768b648a33a7ed878a070d4f6251['h012f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0097a] =  If409768b648a33a7ed878a070d4f6251['h012f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0097b] =  If409768b648a33a7ed878a070d4f6251['h012f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0097c] =  If409768b648a33a7ed878a070d4f6251['h012f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0097d] =  If409768b648a33a7ed878a070d4f6251['h012fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0097e] =  If409768b648a33a7ed878a070d4f6251['h012fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0097f] =  If409768b648a33a7ed878a070d4f6251['h012fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00980] =  If409768b648a33a7ed878a070d4f6251['h01300] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00981] =  If409768b648a33a7ed878a070d4f6251['h01302] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00982] =  If409768b648a33a7ed878a070d4f6251['h01304] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00983] =  If409768b648a33a7ed878a070d4f6251['h01306] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00984] =  If409768b648a33a7ed878a070d4f6251['h01308] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00985] =  If409768b648a33a7ed878a070d4f6251['h0130a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00986] =  If409768b648a33a7ed878a070d4f6251['h0130c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00987] =  If409768b648a33a7ed878a070d4f6251['h0130e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00988] =  If409768b648a33a7ed878a070d4f6251['h01310] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00989] =  If409768b648a33a7ed878a070d4f6251['h01312] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0098a] =  If409768b648a33a7ed878a070d4f6251['h01314] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0098b] =  If409768b648a33a7ed878a070d4f6251['h01316] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0098c] =  If409768b648a33a7ed878a070d4f6251['h01318] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0098d] =  If409768b648a33a7ed878a070d4f6251['h0131a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0098e] =  If409768b648a33a7ed878a070d4f6251['h0131c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0098f] =  If409768b648a33a7ed878a070d4f6251['h0131e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00990] =  If409768b648a33a7ed878a070d4f6251['h01320] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00991] =  If409768b648a33a7ed878a070d4f6251['h01322] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00992] =  If409768b648a33a7ed878a070d4f6251['h01324] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00993] =  If409768b648a33a7ed878a070d4f6251['h01326] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00994] =  If409768b648a33a7ed878a070d4f6251['h01328] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00995] =  If409768b648a33a7ed878a070d4f6251['h0132a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00996] =  If409768b648a33a7ed878a070d4f6251['h0132c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00997] =  If409768b648a33a7ed878a070d4f6251['h0132e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00998] =  If409768b648a33a7ed878a070d4f6251['h01330] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00999] =  If409768b648a33a7ed878a070d4f6251['h01332] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0099a] =  If409768b648a33a7ed878a070d4f6251['h01334] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0099b] =  If409768b648a33a7ed878a070d4f6251['h01336] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0099c] =  If409768b648a33a7ed878a070d4f6251['h01338] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0099d] =  If409768b648a33a7ed878a070d4f6251['h0133a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0099e] =  If409768b648a33a7ed878a070d4f6251['h0133c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h0099f] =  If409768b648a33a7ed878a070d4f6251['h0133e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009a0] =  If409768b648a33a7ed878a070d4f6251['h01340] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009a1] =  If409768b648a33a7ed878a070d4f6251['h01342] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009a2] =  If409768b648a33a7ed878a070d4f6251['h01344] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009a3] =  If409768b648a33a7ed878a070d4f6251['h01346] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009a4] =  If409768b648a33a7ed878a070d4f6251['h01348] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009a5] =  If409768b648a33a7ed878a070d4f6251['h0134a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009a6] =  If409768b648a33a7ed878a070d4f6251['h0134c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009a7] =  If409768b648a33a7ed878a070d4f6251['h0134e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009a8] =  If409768b648a33a7ed878a070d4f6251['h01350] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009a9] =  If409768b648a33a7ed878a070d4f6251['h01352] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009aa] =  If409768b648a33a7ed878a070d4f6251['h01354] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ab] =  If409768b648a33a7ed878a070d4f6251['h01356] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ac] =  If409768b648a33a7ed878a070d4f6251['h01358] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ad] =  If409768b648a33a7ed878a070d4f6251['h0135a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ae] =  If409768b648a33a7ed878a070d4f6251['h0135c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009af] =  If409768b648a33a7ed878a070d4f6251['h0135e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009b0] =  If409768b648a33a7ed878a070d4f6251['h01360] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009b1] =  If409768b648a33a7ed878a070d4f6251['h01362] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009b2] =  If409768b648a33a7ed878a070d4f6251['h01364] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009b3] =  If409768b648a33a7ed878a070d4f6251['h01366] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009b4] =  If409768b648a33a7ed878a070d4f6251['h01368] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009b5] =  If409768b648a33a7ed878a070d4f6251['h0136a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009b6] =  If409768b648a33a7ed878a070d4f6251['h0136c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009b7] =  If409768b648a33a7ed878a070d4f6251['h0136e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009b8] =  If409768b648a33a7ed878a070d4f6251['h01370] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009b9] =  If409768b648a33a7ed878a070d4f6251['h01372] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ba] =  If409768b648a33a7ed878a070d4f6251['h01374] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009bb] =  If409768b648a33a7ed878a070d4f6251['h01376] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009bc] =  If409768b648a33a7ed878a070d4f6251['h01378] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009bd] =  If409768b648a33a7ed878a070d4f6251['h0137a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009be] =  If409768b648a33a7ed878a070d4f6251['h0137c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009bf] =  If409768b648a33a7ed878a070d4f6251['h0137e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009c0] =  If409768b648a33a7ed878a070d4f6251['h01380] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009c1] =  If409768b648a33a7ed878a070d4f6251['h01382] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009c2] =  If409768b648a33a7ed878a070d4f6251['h01384] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009c3] =  If409768b648a33a7ed878a070d4f6251['h01386] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009c4] =  If409768b648a33a7ed878a070d4f6251['h01388] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009c5] =  If409768b648a33a7ed878a070d4f6251['h0138a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009c6] =  If409768b648a33a7ed878a070d4f6251['h0138c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009c7] =  If409768b648a33a7ed878a070d4f6251['h0138e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009c8] =  If409768b648a33a7ed878a070d4f6251['h01390] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009c9] =  If409768b648a33a7ed878a070d4f6251['h01392] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ca] =  If409768b648a33a7ed878a070d4f6251['h01394] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009cb] =  If409768b648a33a7ed878a070d4f6251['h01396] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009cc] =  If409768b648a33a7ed878a070d4f6251['h01398] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009cd] =  If409768b648a33a7ed878a070d4f6251['h0139a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ce] =  If409768b648a33a7ed878a070d4f6251['h0139c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009cf] =  If409768b648a33a7ed878a070d4f6251['h0139e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009d0] =  If409768b648a33a7ed878a070d4f6251['h013a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009d1] =  If409768b648a33a7ed878a070d4f6251['h013a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009d2] =  If409768b648a33a7ed878a070d4f6251['h013a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009d3] =  If409768b648a33a7ed878a070d4f6251['h013a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009d4] =  If409768b648a33a7ed878a070d4f6251['h013a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009d5] =  If409768b648a33a7ed878a070d4f6251['h013aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009d6] =  If409768b648a33a7ed878a070d4f6251['h013ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009d7] =  If409768b648a33a7ed878a070d4f6251['h013ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009d8] =  If409768b648a33a7ed878a070d4f6251['h013b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009d9] =  If409768b648a33a7ed878a070d4f6251['h013b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009da] =  If409768b648a33a7ed878a070d4f6251['h013b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009db] =  If409768b648a33a7ed878a070d4f6251['h013b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009dc] =  If409768b648a33a7ed878a070d4f6251['h013b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009dd] =  If409768b648a33a7ed878a070d4f6251['h013ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009de] =  If409768b648a33a7ed878a070d4f6251['h013bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009df] =  If409768b648a33a7ed878a070d4f6251['h013be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009e0] =  If409768b648a33a7ed878a070d4f6251['h013c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009e1] =  If409768b648a33a7ed878a070d4f6251['h013c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009e2] =  If409768b648a33a7ed878a070d4f6251['h013c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009e3] =  If409768b648a33a7ed878a070d4f6251['h013c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009e4] =  If409768b648a33a7ed878a070d4f6251['h013c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009e5] =  If409768b648a33a7ed878a070d4f6251['h013ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009e6] =  If409768b648a33a7ed878a070d4f6251['h013cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009e7] =  If409768b648a33a7ed878a070d4f6251['h013ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009e8] =  If409768b648a33a7ed878a070d4f6251['h013d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009e9] =  If409768b648a33a7ed878a070d4f6251['h013d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ea] =  If409768b648a33a7ed878a070d4f6251['h013d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009eb] =  If409768b648a33a7ed878a070d4f6251['h013d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ec] =  If409768b648a33a7ed878a070d4f6251['h013d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ed] =  If409768b648a33a7ed878a070d4f6251['h013da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ee] =  If409768b648a33a7ed878a070d4f6251['h013dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ef] =  If409768b648a33a7ed878a070d4f6251['h013de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009f0] =  If409768b648a33a7ed878a070d4f6251['h013e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009f1] =  If409768b648a33a7ed878a070d4f6251['h013e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009f2] =  If409768b648a33a7ed878a070d4f6251['h013e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009f3] =  If409768b648a33a7ed878a070d4f6251['h013e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009f4] =  If409768b648a33a7ed878a070d4f6251['h013e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009f5] =  If409768b648a33a7ed878a070d4f6251['h013ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009f6] =  If409768b648a33a7ed878a070d4f6251['h013ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009f7] =  If409768b648a33a7ed878a070d4f6251['h013ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009f8] =  If409768b648a33a7ed878a070d4f6251['h013f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009f9] =  If409768b648a33a7ed878a070d4f6251['h013f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009fa] =  If409768b648a33a7ed878a070d4f6251['h013f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009fb] =  If409768b648a33a7ed878a070d4f6251['h013f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009fc] =  If409768b648a33a7ed878a070d4f6251['h013f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009fd] =  If409768b648a33a7ed878a070d4f6251['h013fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009fe] =  If409768b648a33a7ed878a070d4f6251['h013fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h009ff] =  If409768b648a33a7ed878a070d4f6251['h013fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a00] =  If409768b648a33a7ed878a070d4f6251['h01400] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a01] =  If409768b648a33a7ed878a070d4f6251['h01402] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a02] =  If409768b648a33a7ed878a070d4f6251['h01404] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a03] =  If409768b648a33a7ed878a070d4f6251['h01406] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a04] =  If409768b648a33a7ed878a070d4f6251['h01408] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a05] =  If409768b648a33a7ed878a070d4f6251['h0140a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a06] =  If409768b648a33a7ed878a070d4f6251['h0140c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a07] =  If409768b648a33a7ed878a070d4f6251['h0140e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a08] =  If409768b648a33a7ed878a070d4f6251['h01410] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a09] =  If409768b648a33a7ed878a070d4f6251['h01412] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a0a] =  If409768b648a33a7ed878a070d4f6251['h01414] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a0b] =  If409768b648a33a7ed878a070d4f6251['h01416] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a0c] =  If409768b648a33a7ed878a070d4f6251['h01418] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a0d] =  If409768b648a33a7ed878a070d4f6251['h0141a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a0e] =  If409768b648a33a7ed878a070d4f6251['h0141c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a0f] =  If409768b648a33a7ed878a070d4f6251['h0141e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a10] =  If409768b648a33a7ed878a070d4f6251['h01420] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a11] =  If409768b648a33a7ed878a070d4f6251['h01422] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a12] =  If409768b648a33a7ed878a070d4f6251['h01424] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a13] =  If409768b648a33a7ed878a070d4f6251['h01426] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a14] =  If409768b648a33a7ed878a070d4f6251['h01428] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a15] =  If409768b648a33a7ed878a070d4f6251['h0142a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a16] =  If409768b648a33a7ed878a070d4f6251['h0142c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a17] =  If409768b648a33a7ed878a070d4f6251['h0142e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a18] =  If409768b648a33a7ed878a070d4f6251['h01430] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a19] =  If409768b648a33a7ed878a070d4f6251['h01432] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a1a] =  If409768b648a33a7ed878a070d4f6251['h01434] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a1b] =  If409768b648a33a7ed878a070d4f6251['h01436] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a1c] =  If409768b648a33a7ed878a070d4f6251['h01438] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a1d] =  If409768b648a33a7ed878a070d4f6251['h0143a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a1e] =  If409768b648a33a7ed878a070d4f6251['h0143c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a1f] =  If409768b648a33a7ed878a070d4f6251['h0143e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a20] =  If409768b648a33a7ed878a070d4f6251['h01440] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a21] =  If409768b648a33a7ed878a070d4f6251['h01442] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a22] =  If409768b648a33a7ed878a070d4f6251['h01444] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a23] =  If409768b648a33a7ed878a070d4f6251['h01446] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a24] =  If409768b648a33a7ed878a070d4f6251['h01448] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a25] =  If409768b648a33a7ed878a070d4f6251['h0144a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a26] =  If409768b648a33a7ed878a070d4f6251['h0144c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a27] =  If409768b648a33a7ed878a070d4f6251['h0144e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a28] =  If409768b648a33a7ed878a070d4f6251['h01450] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a29] =  If409768b648a33a7ed878a070d4f6251['h01452] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a2a] =  If409768b648a33a7ed878a070d4f6251['h01454] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a2b] =  If409768b648a33a7ed878a070d4f6251['h01456] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a2c] =  If409768b648a33a7ed878a070d4f6251['h01458] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a2d] =  If409768b648a33a7ed878a070d4f6251['h0145a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a2e] =  If409768b648a33a7ed878a070d4f6251['h0145c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a2f] =  If409768b648a33a7ed878a070d4f6251['h0145e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a30] =  If409768b648a33a7ed878a070d4f6251['h01460] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a31] =  If409768b648a33a7ed878a070d4f6251['h01462] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a32] =  If409768b648a33a7ed878a070d4f6251['h01464] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a33] =  If409768b648a33a7ed878a070d4f6251['h01466] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a34] =  If409768b648a33a7ed878a070d4f6251['h01468] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a35] =  If409768b648a33a7ed878a070d4f6251['h0146a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a36] =  If409768b648a33a7ed878a070d4f6251['h0146c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a37] =  If409768b648a33a7ed878a070d4f6251['h0146e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a38] =  If409768b648a33a7ed878a070d4f6251['h01470] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a39] =  If409768b648a33a7ed878a070d4f6251['h01472] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a3a] =  If409768b648a33a7ed878a070d4f6251['h01474] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a3b] =  If409768b648a33a7ed878a070d4f6251['h01476] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a3c] =  If409768b648a33a7ed878a070d4f6251['h01478] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a3d] =  If409768b648a33a7ed878a070d4f6251['h0147a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a3e] =  If409768b648a33a7ed878a070d4f6251['h0147c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a3f] =  If409768b648a33a7ed878a070d4f6251['h0147e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a40] =  If409768b648a33a7ed878a070d4f6251['h01480] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a41] =  If409768b648a33a7ed878a070d4f6251['h01482] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a42] =  If409768b648a33a7ed878a070d4f6251['h01484] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a43] =  If409768b648a33a7ed878a070d4f6251['h01486] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a44] =  If409768b648a33a7ed878a070d4f6251['h01488] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a45] =  If409768b648a33a7ed878a070d4f6251['h0148a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a46] =  If409768b648a33a7ed878a070d4f6251['h0148c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a47] =  If409768b648a33a7ed878a070d4f6251['h0148e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a48] =  If409768b648a33a7ed878a070d4f6251['h01490] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a49] =  If409768b648a33a7ed878a070d4f6251['h01492] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a4a] =  If409768b648a33a7ed878a070d4f6251['h01494] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a4b] =  If409768b648a33a7ed878a070d4f6251['h01496] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a4c] =  If409768b648a33a7ed878a070d4f6251['h01498] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a4d] =  If409768b648a33a7ed878a070d4f6251['h0149a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a4e] =  If409768b648a33a7ed878a070d4f6251['h0149c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a4f] =  If409768b648a33a7ed878a070d4f6251['h0149e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a50] =  If409768b648a33a7ed878a070d4f6251['h014a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a51] =  If409768b648a33a7ed878a070d4f6251['h014a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a52] =  If409768b648a33a7ed878a070d4f6251['h014a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a53] =  If409768b648a33a7ed878a070d4f6251['h014a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a54] =  If409768b648a33a7ed878a070d4f6251['h014a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a55] =  If409768b648a33a7ed878a070d4f6251['h014aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a56] =  If409768b648a33a7ed878a070d4f6251['h014ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a57] =  If409768b648a33a7ed878a070d4f6251['h014ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a58] =  If409768b648a33a7ed878a070d4f6251['h014b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a59] =  If409768b648a33a7ed878a070d4f6251['h014b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a5a] =  If409768b648a33a7ed878a070d4f6251['h014b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a5b] =  If409768b648a33a7ed878a070d4f6251['h014b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a5c] =  If409768b648a33a7ed878a070d4f6251['h014b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a5d] =  If409768b648a33a7ed878a070d4f6251['h014ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a5e] =  If409768b648a33a7ed878a070d4f6251['h014bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a5f] =  If409768b648a33a7ed878a070d4f6251['h014be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a60] =  If409768b648a33a7ed878a070d4f6251['h014c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a61] =  If409768b648a33a7ed878a070d4f6251['h014c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a62] =  If409768b648a33a7ed878a070d4f6251['h014c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a63] =  If409768b648a33a7ed878a070d4f6251['h014c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a64] =  If409768b648a33a7ed878a070d4f6251['h014c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a65] =  If409768b648a33a7ed878a070d4f6251['h014ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a66] =  If409768b648a33a7ed878a070d4f6251['h014cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a67] =  If409768b648a33a7ed878a070d4f6251['h014ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a68] =  If409768b648a33a7ed878a070d4f6251['h014d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a69] =  If409768b648a33a7ed878a070d4f6251['h014d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a6a] =  If409768b648a33a7ed878a070d4f6251['h014d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a6b] =  If409768b648a33a7ed878a070d4f6251['h014d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a6c] =  If409768b648a33a7ed878a070d4f6251['h014d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a6d] =  If409768b648a33a7ed878a070d4f6251['h014da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a6e] =  If409768b648a33a7ed878a070d4f6251['h014dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a6f] =  If409768b648a33a7ed878a070d4f6251['h014de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a70] =  If409768b648a33a7ed878a070d4f6251['h014e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a71] =  If409768b648a33a7ed878a070d4f6251['h014e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a72] =  If409768b648a33a7ed878a070d4f6251['h014e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a73] =  If409768b648a33a7ed878a070d4f6251['h014e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a74] =  If409768b648a33a7ed878a070d4f6251['h014e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a75] =  If409768b648a33a7ed878a070d4f6251['h014ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a76] =  If409768b648a33a7ed878a070d4f6251['h014ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a77] =  If409768b648a33a7ed878a070d4f6251['h014ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a78] =  If409768b648a33a7ed878a070d4f6251['h014f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a79] =  If409768b648a33a7ed878a070d4f6251['h014f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a7a] =  If409768b648a33a7ed878a070d4f6251['h014f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a7b] =  If409768b648a33a7ed878a070d4f6251['h014f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a7c] =  If409768b648a33a7ed878a070d4f6251['h014f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a7d] =  If409768b648a33a7ed878a070d4f6251['h014fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a7e] =  If409768b648a33a7ed878a070d4f6251['h014fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a7f] =  If409768b648a33a7ed878a070d4f6251['h014fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a80] =  If409768b648a33a7ed878a070d4f6251['h01500] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a81] =  If409768b648a33a7ed878a070d4f6251['h01502] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a82] =  If409768b648a33a7ed878a070d4f6251['h01504] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a83] =  If409768b648a33a7ed878a070d4f6251['h01506] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a84] =  If409768b648a33a7ed878a070d4f6251['h01508] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a85] =  If409768b648a33a7ed878a070d4f6251['h0150a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a86] =  If409768b648a33a7ed878a070d4f6251['h0150c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a87] =  If409768b648a33a7ed878a070d4f6251['h0150e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a88] =  If409768b648a33a7ed878a070d4f6251['h01510] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a89] =  If409768b648a33a7ed878a070d4f6251['h01512] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a8a] =  If409768b648a33a7ed878a070d4f6251['h01514] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a8b] =  If409768b648a33a7ed878a070d4f6251['h01516] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a8c] =  If409768b648a33a7ed878a070d4f6251['h01518] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a8d] =  If409768b648a33a7ed878a070d4f6251['h0151a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a8e] =  If409768b648a33a7ed878a070d4f6251['h0151c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a8f] =  If409768b648a33a7ed878a070d4f6251['h0151e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a90] =  If409768b648a33a7ed878a070d4f6251['h01520] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a91] =  If409768b648a33a7ed878a070d4f6251['h01522] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a92] =  If409768b648a33a7ed878a070d4f6251['h01524] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a93] =  If409768b648a33a7ed878a070d4f6251['h01526] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a94] =  If409768b648a33a7ed878a070d4f6251['h01528] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a95] =  If409768b648a33a7ed878a070d4f6251['h0152a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a96] =  If409768b648a33a7ed878a070d4f6251['h0152c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a97] =  If409768b648a33a7ed878a070d4f6251['h0152e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a98] =  If409768b648a33a7ed878a070d4f6251['h01530] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a99] =  If409768b648a33a7ed878a070d4f6251['h01532] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a9a] =  If409768b648a33a7ed878a070d4f6251['h01534] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a9b] =  If409768b648a33a7ed878a070d4f6251['h01536] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a9c] =  If409768b648a33a7ed878a070d4f6251['h01538] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a9d] =  If409768b648a33a7ed878a070d4f6251['h0153a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a9e] =  If409768b648a33a7ed878a070d4f6251['h0153c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00a9f] =  If409768b648a33a7ed878a070d4f6251['h0153e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aa0] =  If409768b648a33a7ed878a070d4f6251['h01540] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aa1] =  If409768b648a33a7ed878a070d4f6251['h01542] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aa2] =  If409768b648a33a7ed878a070d4f6251['h01544] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aa3] =  If409768b648a33a7ed878a070d4f6251['h01546] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aa4] =  If409768b648a33a7ed878a070d4f6251['h01548] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aa5] =  If409768b648a33a7ed878a070d4f6251['h0154a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aa6] =  If409768b648a33a7ed878a070d4f6251['h0154c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aa7] =  If409768b648a33a7ed878a070d4f6251['h0154e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aa8] =  If409768b648a33a7ed878a070d4f6251['h01550] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aa9] =  If409768b648a33a7ed878a070d4f6251['h01552] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aaa] =  If409768b648a33a7ed878a070d4f6251['h01554] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aab] =  If409768b648a33a7ed878a070d4f6251['h01556] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aac] =  If409768b648a33a7ed878a070d4f6251['h01558] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aad] =  If409768b648a33a7ed878a070d4f6251['h0155a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aae] =  If409768b648a33a7ed878a070d4f6251['h0155c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aaf] =  If409768b648a33a7ed878a070d4f6251['h0155e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ab0] =  If409768b648a33a7ed878a070d4f6251['h01560] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ab1] =  If409768b648a33a7ed878a070d4f6251['h01562] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ab2] =  If409768b648a33a7ed878a070d4f6251['h01564] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ab3] =  If409768b648a33a7ed878a070d4f6251['h01566] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ab4] =  If409768b648a33a7ed878a070d4f6251['h01568] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ab5] =  If409768b648a33a7ed878a070d4f6251['h0156a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ab6] =  If409768b648a33a7ed878a070d4f6251['h0156c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ab7] =  If409768b648a33a7ed878a070d4f6251['h0156e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ab8] =  If409768b648a33a7ed878a070d4f6251['h01570] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ab9] =  If409768b648a33a7ed878a070d4f6251['h01572] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aba] =  If409768b648a33a7ed878a070d4f6251['h01574] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00abb] =  If409768b648a33a7ed878a070d4f6251['h01576] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00abc] =  If409768b648a33a7ed878a070d4f6251['h01578] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00abd] =  If409768b648a33a7ed878a070d4f6251['h0157a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00abe] =  If409768b648a33a7ed878a070d4f6251['h0157c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00abf] =  If409768b648a33a7ed878a070d4f6251['h0157e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ac0] =  If409768b648a33a7ed878a070d4f6251['h01580] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ac1] =  If409768b648a33a7ed878a070d4f6251['h01582] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ac2] =  If409768b648a33a7ed878a070d4f6251['h01584] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ac3] =  If409768b648a33a7ed878a070d4f6251['h01586] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ac4] =  If409768b648a33a7ed878a070d4f6251['h01588] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ac5] =  If409768b648a33a7ed878a070d4f6251['h0158a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ac6] =  If409768b648a33a7ed878a070d4f6251['h0158c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ac7] =  If409768b648a33a7ed878a070d4f6251['h0158e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ac8] =  If409768b648a33a7ed878a070d4f6251['h01590] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ac9] =  If409768b648a33a7ed878a070d4f6251['h01592] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aca] =  If409768b648a33a7ed878a070d4f6251['h01594] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00acb] =  If409768b648a33a7ed878a070d4f6251['h01596] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00acc] =  If409768b648a33a7ed878a070d4f6251['h01598] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00acd] =  If409768b648a33a7ed878a070d4f6251['h0159a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ace] =  If409768b648a33a7ed878a070d4f6251['h0159c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00acf] =  If409768b648a33a7ed878a070d4f6251['h0159e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ad0] =  If409768b648a33a7ed878a070d4f6251['h015a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ad1] =  If409768b648a33a7ed878a070d4f6251['h015a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ad2] =  If409768b648a33a7ed878a070d4f6251['h015a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ad3] =  If409768b648a33a7ed878a070d4f6251['h015a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ad4] =  If409768b648a33a7ed878a070d4f6251['h015a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ad5] =  If409768b648a33a7ed878a070d4f6251['h015aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ad6] =  If409768b648a33a7ed878a070d4f6251['h015ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ad7] =  If409768b648a33a7ed878a070d4f6251['h015ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ad8] =  If409768b648a33a7ed878a070d4f6251['h015b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ad9] =  If409768b648a33a7ed878a070d4f6251['h015b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ada] =  If409768b648a33a7ed878a070d4f6251['h015b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00adb] =  If409768b648a33a7ed878a070d4f6251['h015b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00adc] =  If409768b648a33a7ed878a070d4f6251['h015b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00add] =  If409768b648a33a7ed878a070d4f6251['h015ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ade] =  If409768b648a33a7ed878a070d4f6251['h015bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00adf] =  If409768b648a33a7ed878a070d4f6251['h015be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ae0] =  If409768b648a33a7ed878a070d4f6251['h015c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ae1] =  If409768b648a33a7ed878a070d4f6251['h015c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ae2] =  If409768b648a33a7ed878a070d4f6251['h015c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ae3] =  If409768b648a33a7ed878a070d4f6251['h015c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ae4] =  If409768b648a33a7ed878a070d4f6251['h015c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ae5] =  If409768b648a33a7ed878a070d4f6251['h015ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ae6] =  If409768b648a33a7ed878a070d4f6251['h015cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ae7] =  If409768b648a33a7ed878a070d4f6251['h015ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ae8] =  If409768b648a33a7ed878a070d4f6251['h015d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ae9] =  If409768b648a33a7ed878a070d4f6251['h015d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aea] =  If409768b648a33a7ed878a070d4f6251['h015d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aeb] =  If409768b648a33a7ed878a070d4f6251['h015d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aec] =  If409768b648a33a7ed878a070d4f6251['h015d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aed] =  If409768b648a33a7ed878a070d4f6251['h015da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aee] =  If409768b648a33a7ed878a070d4f6251['h015dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aef] =  If409768b648a33a7ed878a070d4f6251['h015de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00af0] =  If409768b648a33a7ed878a070d4f6251['h015e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00af1] =  If409768b648a33a7ed878a070d4f6251['h015e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00af2] =  If409768b648a33a7ed878a070d4f6251['h015e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00af3] =  If409768b648a33a7ed878a070d4f6251['h015e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00af4] =  If409768b648a33a7ed878a070d4f6251['h015e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00af5] =  If409768b648a33a7ed878a070d4f6251['h015ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00af6] =  If409768b648a33a7ed878a070d4f6251['h015ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00af7] =  If409768b648a33a7ed878a070d4f6251['h015ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00af8] =  If409768b648a33a7ed878a070d4f6251['h015f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00af9] =  If409768b648a33a7ed878a070d4f6251['h015f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00afa] =  If409768b648a33a7ed878a070d4f6251['h015f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00afb] =  If409768b648a33a7ed878a070d4f6251['h015f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00afc] =  If409768b648a33a7ed878a070d4f6251['h015f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00afd] =  If409768b648a33a7ed878a070d4f6251['h015fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00afe] =  If409768b648a33a7ed878a070d4f6251['h015fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00aff] =  If409768b648a33a7ed878a070d4f6251['h015fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b00] =  If409768b648a33a7ed878a070d4f6251['h01600] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b01] =  If409768b648a33a7ed878a070d4f6251['h01602] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b02] =  If409768b648a33a7ed878a070d4f6251['h01604] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b03] =  If409768b648a33a7ed878a070d4f6251['h01606] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b04] =  If409768b648a33a7ed878a070d4f6251['h01608] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b05] =  If409768b648a33a7ed878a070d4f6251['h0160a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b06] =  If409768b648a33a7ed878a070d4f6251['h0160c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b07] =  If409768b648a33a7ed878a070d4f6251['h0160e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b08] =  If409768b648a33a7ed878a070d4f6251['h01610] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b09] =  If409768b648a33a7ed878a070d4f6251['h01612] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b0a] =  If409768b648a33a7ed878a070d4f6251['h01614] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b0b] =  If409768b648a33a7ed878a070d4f6251['h01616] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b0c] =  If409768b648a33a7ed878a070d4f6251['h01618] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b0d] =  If409768b648a33a7ed878a070d4f6251['h0161a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b0e] =  If409768b648a33a7ed878a070d4f6251['h0161c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b0f] =  If409768b648a33a7ed878a070d4f6251['h0161e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b10] =  If409768b648a33a7ed878a070d4f6251['h01620] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b11] =  If409768b648a33a7ed878a070d4f6251['h01622] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b12] =  If409768b648a33a7ed878a070d4f6251['h01624] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b13] =  If409768b648a33a7ed878a070d4f6251['h01626] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b14] =  If409768b648a33a7ed878a070d4f6251['h01628] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b15] =  If409768b648a33a7ed878a070d4f6251['h0162a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b16] =  If409768b648a33a7ed878a070d4f6251['h0162c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b17] =  If409768b648a33a7ed878a070d4f6251['h0162e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b18] =  If409768b648a33a7ed878a070d4f6251['h01630] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b19] =  If409768b648a33a7ed878a070d4f6251['h01632] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b1a] =  If409768b648a33a7ed878a070d4f6251['h01634] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b1b] =  If409768b648a33a7ed878a070d4f6251['h01636] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b1c] =  If409768b648a33a7ed878a070d4f6251['h01638] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b1d] =  If409768b648a33a7ed878a070d4f6251['h0163a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b1e] =  If409768b648a33a7ed878a070d4f6251['h0163c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b1f] =  If409768b648a33a7ed878a070d4f6251['h0163e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b20] =  If409768b648a33a7ed878a070d4f6251['h01640] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b21] =  If409768b648a33a7ed878a070d4f6251['h01642] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b22] =  If409768b648a33a7ed878a070d4f6251['h01644] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b23] =  If409768b648a33a7ed878a070d4f6251['h01646] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b24] =  If409768b648a33a7ed878a070d4f6251['h01648] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b25] =  If409768b648a33a7ed878a070d4f6251['h0164a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b26] =  If409768b648a33a7ed878a070d4f6251['h0164c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b27] =  If409768b648a33a7ed878a070d4f6251['h0164e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b28] =  If409768b648a33a7ed878a070d4f6251['h01650] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b29] =  If409768b648a33a7ed878a070d4f6251['h01652] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b2a] =  If409768b648a33a7ed878a070d4f6251['h01654] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b2b] =  If409768b648a33a7ed878a070d4f6251['h01656] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b2c] =  If409768b648a33a7ed878a070d4f6251['h01658] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b2d] =  If409768b648a33a7ed878a070d4f6251['h0165a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b2e] =  If409768b648a33a7ed878a070d4f6251['h0165c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b2f] =  If409768b648a33a7ed878a070d4f6251['h0165e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b30] =  If409768b648a33a7ed878a070d4f6251['h01660] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b31] =  If409768b648a33a7ed878a070d4f6251['h01662] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b32] =  If409768b648a33a7ed878a070d4f6251['h01664] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b33] =  If409768b648a33a7ed878a070d4f6251['h01666] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b34] =  If409768b648a33a7ed878a070d4f6251['h01668] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b35] =  If409768b648a33a7ed878a070d4f6251['h0166a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b36] =  If409768b648a33a7ed878a070d4f6251['h0166c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b37] =  If409768b648a33a7ed878a070d4f6251['h0166e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b38] =  If409768b648a33a7ed878a070d4f6251['h01670] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b39] =  If409768b648a33a7ed878a070d4f6251['h01672] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b3a] =  If409768b648a33a7ed878a070d4f6251['h01674] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b3b] =  If409768b648a33a7ed878a070d4f6251['h01676] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b3c] =  If409768b648a33a7ed878a070d4f6251['h01678] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b3d] =  If409768b648a33a7ed878a070d4f6251['h0167a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b3e] =  If409768b648a33a7ed878a070d4f6251['h0167c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b3f] =  If409768b648a33a7ed878a070d4f6251['h0167e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b40] =  If409768b648a33a7ed878a070d4f6251['h01680] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b41] =  If409768b648a33a7ed878a070d4f6251['h01682] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b42] =  If409768b648a33a7ed878a070d4f6251['h01684] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b43] =  If409768b648a33a7ed878a070d4f6251['h01686] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b44] =  If409768b648a33a7ed878a070d4f6251['h01688] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b45] =  If409768b648a33a7ed878a070d4f6251['h0168a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b46] =  If409768b648a33a7ed878a070d4f6251['h0168c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b47] =  If409768b648a33a7ed878a070d4f6251['h0168e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b48] =  If409768b648a33a7ed878a070d4f6251['h01690] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b49] =  If409768b648a33a7ed878a070d4f6251['h01692] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b4a] =  If409768b648a33a7ed878a070d4f6251['h01694] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b4b] =  If409768b648a33a7ed878a070d4f6251['h01696] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b4c] =  If409768b648a33a7ed878a070d4f6251['h01698] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b4d] =  If409768b648a33a7ed878a070d4f6251['h0169a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b4e] =  If409768b648a33a7ed878a070d4f6251['h0169c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b4f] =  If409768b648a33a7ed878a070d4f6251['h0169e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b50] =  If409768b648a33a7ed878a070d4f6251['h016a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b51] =  If409768b648a33a7ed878a070d4f6251['h016a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b52] =  If409768b648a33a7ed878a070d4f6251['h016a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b53] =  If409768b648a33a7ed878a070d4f6251['h016a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b54] =  If409768b648a33a7ed878a070d4f6251['h016a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b55] =  If409768b648a33a7ed878a070d4f6251['h016aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b56] =  If409768b648a33a7ed878a070d4f6251['h016ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b57] =  If409768b648a33a7ed878a070d4f6251['h016ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b58] =  If409768b648a33a7ed878a070d4f6251['h016b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b59] =  If409768b648a33a7ed878a070d4f6251['h016b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b5a] =  If409768b648a33a7ed878a070d4f6251['h016b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b5b] =  If409768b648a33a7ed878a070d4f6251['h016b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b5c] =  If409768b648a33a7ed878a070d4f6251['h016b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b5d] =  If409768b648a33a7ed878a070d4f6251['h016ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b5e] =  If409768b648a33a7ed878a070d4f6251['h016bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b5f] =  If409768b648a33a7ed878a070d4f6251['h016be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b60] =  If409768b648a33a7ed878a070d4f6251['h016c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b61] =  If409768b648a33a7ed878a070d4f6251['h016c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b62] =  If409768b648a33a7ed878a070d4f6251['h016c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b63] =  If409768b648a33a7ed878a070d4f6251['h016c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b64] =  If409768b648a33a7ed878a070d4f6251['h016c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b65] =  If409768b648a33a7ed878a070d4f6251['h016ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b66] =  If409768b648a33a7ed878a070d4f6251['h016cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b67] =  If409768b648a33a7ed878a070d4f6251['h016ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b68] =  If409768b648a33a7ed878a070d4f6251['h016d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b69] =  If409768b648a33a7ed878a070d4f6251['h016d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b6a] =  If409768b648a33a7ed878a070d4f6251['h016d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b6b] =  If409768b648a33a7ed878a070d4f6251['h016d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b6c] =  If409768b648a33a7ed878a070d4f6251['h016d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b6d] =  If409768b648a33a7ed878a070d4f6251['h016da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b6e] =  If409768b648a33a7ed878a070d4f6251['h016dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b6f] =  If409768b648a33a7ed878a070d4f6251['h016de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b70] =  If409768b648a33a7ed878a070d4f6251['h016e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b71] =  If409768b648a33a7ed878a070d4f6251['h016e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b72] =  If409768b648a33a7ed878a070d4f6251['h016e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b73] =  If409768b648a33a7ed878a070d4f6251['h016e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b74] =  If409768b648a33a7ed878a070d4f6251['h016e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b75] =  If409768b648a33a7ed878a070d4f6251['h016ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b76] =  If409768b648a33a7ed878a070d4f6251['h016ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b77] =  If409768b648a33a7ed878a070d4f6251['h016ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b78] =  If409768b648a33a7ed878a070d4f6251['h016f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b79] =  If409768b648a33a7ed878a070d4f6251['h016f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b7a] =  If409768b648a33a7ed878a070d4f6251['h016f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b7b] =  If409768b648a33a7ed878a070d4f6251['h016f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b7c] =  If409768b648a33a7ed878a070d4f6251['h016f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b7d] =  If409768b648a33a7ed878a070d4f6251['h016fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b7e] =  If409768b648a33a7ed878a070d4f6251['h016fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b7f] =  If409768b648a33a7ed878a070d4f6251['h016fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b80] =  If409768b648a33a7ed878a070d4f6251['h01700] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b81] =  If409768b648a33a7ed878a070d4f6251['h01702] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b82] =  If409768b648a33a7ed878a070d4f6251['h01704] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b83] =  If409768b648a33a7ed878a070d4f6251['h01706] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b84] =  If409768b648a33a7ed878a070d4f6251['h01708] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b85] =  If409768b648a33a7ed878a070d4f6251['h0170a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b86] =  If409768b648a33a7ed878a070d4f6251['h0170c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b87] =  If409768b648a33a7ed878a070d4f6251['h0170e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b88] =  If409768b648a33a7ed878a070d4f6251['h01710] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b89] =  If409768b648a33a7ed878a070d4f6251['h01712] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b8a] =  If409768b648a33a7ed878a070d4f6251['h01714] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b8b] =  If409768b648a33a7ed878a070d4f6251['h01716] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b8c] =  If409768b648a33a7ed878a070d4f6251['h01718] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b8d] =  If409768b648a33a7ed878a070d4f6251['h0171a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b8e] =  If409768b648a33a7ed878a070d4f6251['h0171c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b8f] =  If409768b648a33a7ed878a070d4f6251['h0171e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b90] =  If409768b648a33a7ed878a070d4f6251['h01720] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b91] =  If409768b648a33a7ed878a070d4f6251['h01722] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b92] =  If409768b648a33a7ed878a070d4f6251['h01724] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b93] =  If409768b648a33a7ed878a070d4f6251['h01726] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b94] =  If409768b648a33a7ed878a070d4f6251['h01728] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b95] =  If409768b648a33a7ed878a070d4f6251['h0172a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b96] =  If409768b648a33a7ed878a070d4f6251['h0172c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b97] =  If409768b648a33a7ed878a070d4f6251['h0172e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b98] =  If409768b648a33a7ed878a070d4f6251['h01730] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b99] =  If409768b648a33a7ed878a070d4f6251['h01732] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b9a] =  If409768b648a33a7ed878a070d4f6251['h01734] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b9b] =  If409768b648a33a7ed878a070d4f6251['h01736] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b9c] =  If409768b648a33a7ed878a070d4f6251['h01738] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b9d] =  If409768b648a33a7ed878a070d4f6251['h0173a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b9e] =  If409768b648a33a7ed878a070d4f6251['h0173c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00b9f] =  If409768b648a33a7ed878a070d4f6251['h0173e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ba0] =  If409768b648a33a7ed878a070d4f6251['h01740] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ba1] =  If409768b648a33a7ed878a070d4f6251['h01742] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ba2] =  If409768b648a33a7ed878a070d4f6251['h01744] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ba3] =  If409768b648a33a7ed878a070d4f6251['h01746] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ba4] =  If409768b648a33a7ed878a070d4f6251['h01748] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ba5] =  If409768b648a33a7ed878a070d4f6251['h0174a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ba6] =  If409768b648a33a7ed878a070d4f6251['h0174c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ba7] =  If409768b648a33a7ed878a070d4f6251['h0174e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ba8] =  If409768b648a33a7ed878a070d4f6251['h01750] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ba9] =  If409768b648a33a7ed878a070d4f6251['h01752] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00baa] =  If409768b648a33a7ed878a070d4f6251['h01754] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bab] =  If409768b648a33a7ed878a070d4f6251['h01756] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bac] =  If409768b648a33a7ed878a070d4f6251['h01758] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bad] =  If409768b648a33a7ed878a070d4f6251['h0175a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bae] =  If409768b648a33a7ed878a070d4f6251['h0175c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00baf] =  If409768b648a33a7ed878a070d4f6251['h0175e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bb0] =  If409768b648a33a7ed878a070d4f6251['h01760] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bb1] =  If409768b648a33a7ed878a070d4f6251['h01762] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bb2] =  If409768b648a33a7ed878a070d4f6251['h01764] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bb3] =  If409768b648a33a7ed878a070d4f6251['h01766] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bb4] =  If409768b648a33a7ed878a070d4f6251['h01768] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bb5] =  If409768b648a33a7ed878a070d4f6251['h0176a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bb6] =  If409768b648a33a7ed878a070d4f6251['h0176c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bb7] =  If409768b648a33a7ed878a070d4f6251['h0176e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bb8] =  If409768b648a33a7ed878a070d4f6251['h01770] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bb9] =  If409768b648a33a7ed878a070d4f6251['h01772] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bba] =  If409768b648a33a7ed878a070d4f6251['h01774] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bbb] =  If409768b648a33a7ed878a070d4f6251['h01776] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bbc] =  If409768b648a33a7ed878a070d4f6251['h01778] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bbd] =  If409768b648a33a7ed878a070d4f6251['h0177a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bbe] =  If409768b648a33a7ed878a070d4f6251['h0177c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bbf] =  If409768b648a33a7ed878a070d4f6251['h0177e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bc0] =  If409768b648a33a7ed878a070d4f6251['h01780] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bc1] =  If409768b648a33a7ed878a070d4f6251['h01782] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bc2] =  If409768b648a33a7ed878a070d4f6251['h01784] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bc3] =  If409768b648a33a7ed878a070d4f6251['h01786] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bc4] =  If409768b648a33a7ed878a070d4f6251['h01788] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bc5] =  If409768b648a33a7ed878a070d4f6251['h0178a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bc6] =  If409768b648a33a7ed878a070d4f6251['h0178c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bc7] =  If409768b648a33a7ed878a070d4f6251['h0178e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bc8] =  If409768b648a33a7ed878a070d4f6251['h01790] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bc9] =  If409768b648a33a7ed878a070d4f6251['h01792] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bca] =  If409768b648a33a7ed878a070d4f6251['h01794] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bcb] =  If409768b648a33a7ed878a070d4f6251['h01796] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bcc] =  If409768b648a33a7ed878a070d4f6251['h01798] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bcd] =  If409768b648a33a7ed878a070d4f6251['h0179a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bce] =  If409768b648a33a7ed878a070d4f6251['h0179c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bcf] =  If409768b648a33a7ed878a070d4f6251['h0179e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bd0] =  If409768b648a33a7ed878a070d4f6251['h017a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bd1] =  If409768b648a33a7ed878a070d4f6251['h017a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bd2] =  If409768b648a33a7ed878a070d4f6251['h017a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bd3] =  If409768b648a33a7ed878a070d4f6251['h017a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bd4] =  If409768b648a33a7ed878a070d4f6251['h017a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bd5] =  If409768b648a33a7ed878a070d4f6251['h017aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bd6] =  If409768b648a33a7ed878a070d4f6251['h017ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bd7] =  If409768b648a33a7ed878a070d4f6251['h017ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bd8] =  If409768b648a33a7ed878a070d4f6251['h017b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bd9] =  If409768b648a33a7ed878a070d4f6251['h017b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bda] =  If409768b648a33a7ed878a070d4f6251['h017b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bdb] =  If409768b648a33a7ed878a070d4f6251['h017b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bdc] =  If409768b648a33a7ed878a070d4f6251['h017b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bdd] =  If409768b648a33a7ed878a070d4f6251['h017ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bde] =  If409768b648a33a7ed878a070d4f6251['h017bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bdf] =  If409768b648a33a7ed878a070d4f6251['h017be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00be0] =  If409768b648a33a7ed878a070d4f6251['h017c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00be1] =  If409768b648a33a7ed878a070d4f6251['h017c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00be2] =  If409768b648a33a7ed878a070d4f6251['h017c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00be3] =  If409768b648a33a7ed878a070d4f6251['h017c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00be4] =  If409768b648a33a7ed878a070d4f6251['h017c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00be5] =  If409768b648a33a7ed878a070d4f6251['h017ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00be6] =  If409768b648a33a7ed878a070d4f6251['h017cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00be7] =  If409768b648a33a7ed878a070d4f6251['h017ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00be8] =  If409768b648a33a7ed878a070d4f6251['h017d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00be9] =  If409768b648a33a7ed878a070d4f6251['h017d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bea] =  If409768b648a33a7ed878a070d4f6251['h017d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00beb] =  If409768b648a33a7ed878a070d4f6251['h017d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bec] =  If409768b648a33a7ed878a070d4f6251['h017d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bed] =  If409768b648a33a7ed878a070d4f6251['h017da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bee] =  If409768b648a33a7ed878a070d4f6251['h017dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bef] =  If409768b648a33a7ed878a070d4f6251['h017de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bf0] =  If409768b648a33a7ed878a070d4f6251['h017e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bf1] =  If409768b648a33a7ed878a070d4f6251['h017e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bf2] =  If409768b648a33a7ed878a070d4f6251['h017e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bf3] =  If409768b648a33a7ed878a070d4f6251['h017e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bf4] =  If409768b648a33a7ed878a070d4f6251['h017e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bf5] =  If409768b648a33a7ed878a070d4f6251['h017ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bf6] =  If409768b648a33a7ed878a070d4f6251['h017ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bf7] =  If409768b648a33a7ed878a070d4f6251['h017ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bf8] =  If409768b648a33a7ed878a070d4f6251['h017f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bf9] =  If409768b648a33a7ed878a070d4f6251['h017f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bfa] =  If409768b648a33a7ed878a070d4f6251['h017f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bfb] =  If409768b648a33a7ed878a070d4f6251['h017f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bfc] =  If409768b648a33a7ed878a070d4f6251['h017f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bfd] =  If409768b648a33a7ed878a070d4f6251['h017fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bfe] =  If409768b648a33a7ed878a070d4f6251['h017fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00bff] =  If409768b648a33a7ed878a070d4f6251['h017fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c00] =  If409768b648a33a7ed878a070d4f6251['h01800] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c01] =  If409768b648a33a7ed878a070d4f6251['h01802] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c02] =  If409768b648a33a7ed878a070d4f6251['h01804] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c03] =  If409768b648a33a7ed878a070d4f6251['h01806] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c04] =  If409768b648a33a7ed878a070d4f6251['h01808] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c05] =  If409768b648a33a7ed878a070d4f6251['h0180a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c06] =  If409768b648a33a7ed878a070d4f6251['h0180c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c07] =  If409768b648a33a7ed878a070d4f6251['h0180e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c08] =  If409768b648a33a7ed878a070d4f6251['h01810] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c09] =  If409768b648a33a7ed878a070d4f6251['h01812] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c0a] =  If409768b648a33a7ed878a070d4f6251['h01814] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c0b] =  If409768b648a33a7ed878a070d4f6251['h01816] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c0c] =  If409768b648a33a7ed878a070d4f6251['h01818] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c0d] =  If409768b648a33a7ed878a070d4f6251['h0181a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c0e] =  If409768b648a33a7ed878a070d4f6251['h0181c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c0f] =  If409768b648a33a7ed878a070d4f6251['h0181e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c10] =  If409768b648a33a7ed878a070d4f6251['h01820] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c11] =  If409768b648a33a7ed878a070d4f6251['h01822] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c12] =  If409768b648a33a7ed878a070d4f6251['h01824] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c13] =  If409768b648a33a7ed878a070d4f6251['h01826] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c14] =  If409768b648a33a7ed878a070d4f6251['h01828] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c15] =  If409768b648a33a7ed878a070d4f6251['h0182a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c16] =  If409768b648a33a7ed878a070d4f6251['h0182c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c17] =  If409768b648a33a7ed878a070d4f6251['h0182e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c18] =  If409768b648a33a7ed878a070d4f6251['h01830] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c19] =  If409768b648a33a7ed878a070d4f6251['h01832] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c1a] =  If409768b648a33a7ed878a070d4f6251['h01834] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c1b] =  If409768b648a33a7ed878a070d4f6251['h01836] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c1c] =  If409768b648a33a7ed878a070d4f6251['h01838] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c1d] =  If409768b648a33a7ed878a070d4f6251['h0183a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c1e] =  If409768b648a33a7ed878a070d4f6251['h0183c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c1f] =  If409768b648a33a7ed878a070d4f6251['h0183e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c20] =  If409768b648a33a7ed878a070d4f6251['h01840] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c21] =  If409768b648a33a7ed878a070d4f6251['h01842] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c22] =  If409768b648a33a7ed878a070d4f6251['h01844] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c23] =  If409768b648a33a7ed878a070d4f6251['h01846] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c24] =  If409768b648a33a7ed878a070d4f6251['h01848] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c25] =  If409768b648a33a7ed878a070d4f6251['h0184a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c26] =  If409768b648a33a7ed878a070d4f6251['h0184c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c27] =  If409768b648a33a7ed878a070d4f6251['h0184e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c28] =  If409768b648a33a7ed878a070d4f6251['h01850] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c29] =  If409768b648a33a7ed878a070d4f6251['h01852] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c2a] =  If409768b648a33a7ed878a070d4f6251['h01854] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c2b] =  If409768b648a33a7ed878a070d4f6251['h01856] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c2c] =  If409768b648a33a7ed878a070d4f6251['h01858] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c2d] =  If409768b648a33a7ed878a070d4f6251['h0185a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c2e] =  If409768b648a33a7ed878a070d4f6251['h0185c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c2f] =  If409768b648a33a7ed878a070d4f6251['h0185e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c30] =  If409768b648a33a7ed878a070d4f6251['h01860] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c31] =  If409768b648a33a7ed878a070d4f6251['h01862] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c32] =  If409768b648a33a7ed878a070d4f6251['h01864] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c33] =  If409768b648a33a7ed878a070d4f6251['h01866] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c34] =  If409768b648a33a7ed878a070d4f6251['h01868] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c35] =  If409768b648a33a7ed878a070d4f6251['h0186a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c36] =  If409768b648a33a7ed878a070d4f6251['h0186c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c37] =  If409768b648a33a7ed878a070d4f6251['h0186e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c38] =  If409768b648a33a7ed878a070d4f6251['h01870] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c39] =  If409768b648a33a7ed878a070d4f6251['h01872] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c3a] =  If409768b648a33a7ed878a070d4f6251['h01874] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c3b] =  If409768b648a33a7ed878a070d4f6251['h01876] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c3c] =  If409768b648a33a7ed878a070d4f6251['h01878] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c3d] =  If409768b648a33a7ed878a070d4f6251['h0187a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c3e] =  If409768b648a33a7ed878a070d4f6251['h0187c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c3f] =  If409768b648a33a7ed878a070d4f6251['h0187e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c40] =  If409768b648a33a7ed878a070d4f6251['h01880] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c41] =  If409768b648a33a7ed878a070d4f6251['h01882] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c42] =  If409768b648a33a7ed878a070d4f6251['h01884] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c43] =  If409768b648a33a7ed878a070d4f6251['h01886] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c44] =  If409768b648a33a7ed878a070d4f6251['h01888] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c45] =  If409768b648a33a7ed878a070d4f6251['h0188a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c46] =  If409768b648a33a7ed878a070d4f6251['h0188c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c47] =  If409768b648a33a7ed878a070d4f6251['h0188e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c48] =  If409768b648a33a7ed878a070d4f6251['h01890] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c49] =  If409768b648a33a7ed878a070d4f6251['h01892] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c4a] =  If409768b648a33a7ed878a070d4f6251['h01894] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c4b] =  If409768b648a33a7ed878a070d4f6251['h01896] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c4c] =  If409768b648a33a7ed878a070d4f6251['h01898] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c4d] =  If409768b648a33a7ed878a070d4f6251['h0189a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c4e] =  If409768b648a33a7ed878a070d4f6251['h0189c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c4f] =  If409768b648a33a7ed878a070d4f6251['h0189e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c50] =  If409768b648a33a7ed878a070d4f6251['h018a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c51] =  If409768b648a33a7ed878a070d4f6251['h018a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c52] =  If409768b648a33a7ed878a070d4f6251['h018a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c53] =  If409768b648a33a7ed878a070d4f6251['h018a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c54] =  If409768b648a33a7ed878a070d4f6251['h018a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c55] =  If409768b648a33a7ed878a070d4f6251['h018aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c56] =  If409768b648a33a7ed878a070d4f6251['h018ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c57] =  If409768b648a33a7ed878a070d4f6251['h018ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c58] =  If409768b648a33a7ed878a070d4f6251['h018b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c59] =  If409768b648a33a7ed878a070d4f6251['h018b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c5a] =  If409768b648a33a7ed878a070d4f6251['h018b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c5b] =  If409768b648a33a7ed878a070d4f6251['h018b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c5c] =  If409768b648a33a7ed878a070d4f6251['h018b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c5d] =  If409768b648a33a7ed878a070d4f6251['h018ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c5e] =  If409768b648a33a7ed878a070d4f6251['h018bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c5f] =  If409768b648a33a7ed878a070d4f6251['h018be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c60] =  If409768b648a33a7ed878a070d4f6251['h018c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c61] =  If409768b648a33a7ed878a070d4f6251['h018c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c62] =  If409768b648a33a7ed878a070d4f6251['h018c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c63] =  If409768b648a33a7ed878a070d4f6251['h018c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c64] =  If409768b648a33a7ed878a070d4f6251['h018c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c65] =  If409768b648a33a7ed878a070d4f6251['h018ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c66] =  If409768b648a33a7ed878a070d4f6251['h018cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c67] =  If409768b648a33a7ed878a070d4f6251['h018ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c68] =  If409768b648a33a7ed878a070d4f6251['h018d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c69] =  If409768b648a33a7ed878a070d4f6251['h018d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c6a] =  If409768b648a33a7ed878a070d4f6251['h018d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c6b] =  If409768b648a33a7ed878a070d4f6251['h018d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c6c] =  If409768b648a33a7ed878a070d4f6251['h018d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c6d] =  If409768b648a33a7ed878a070d4f6251['h018da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c6e] =  If409768b648a33a7ed878a070d4f6251['h018dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c6f] =  If409768b648a33a7ed878a070d4f6251['h018de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c70] =  If409768b648a33a7ed878a070d4f6251['h018e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c71] =  If409768b648a33a7ed878a070d4f6251['h018e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c72] =  If409768b648a33a7ed878a070d4f6251['h018e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c73] =  If409768b648a33a7ed878a070d4f6251['h018e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c74] =  If409768b648a33a7ed878a070d4f6251['h018e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c75] =  If409768b648a33a7ed878a070d4f6251['h018ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c76] =  If409768b648a33a7ed878a070d4f6251['h018ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c77] =  If409768b648a33a7ed878a070d4f6251['h018ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c78] =  If409768b648a33a7ed878a070d4f6251['h018f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c79] =  If409768b648a33a7ed878a070d4f6251['h018f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c7a] =  If409768b648a33a7ed878a070d4f6251['h018f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c7b] =  If409768b648a33a7ed878a070d4f6251['h018f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c7c] =  If409768b648a33a7ed878a070d4f6251['h018f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c7d] =  If409768b648a33a7ed878a070d4f6251['h018fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c7e] =  If409768b648a33a7ed878a070d4f6251['h018fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c7f] =  If409768b648a33a7ed878a070d4f6251['h018fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c80] =  If409768b648a33a7ed878a070d4f6251['h01900] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c81] =  If409768b648a33a7ed878a070d4f6251['h01902] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c82] =  If409768b648a33a7ed878a070d4f6251['h01904] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c83] =  If409768b648a33a7ed878a070d4f6251['h01906] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c84] =  If409768b648a33a7ed878a070d4f6251['h01908] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c85] =  If409768b648a33a7ed878a070d4f6251['h0190a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c86] =  If409768b648a33a7ed878a070d4f6251['h0190c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c87] =  If409768b648a33a7ed878a070d4f6251['h0190e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c88] =  If409768b648a33a7ed878a070d4f6251['h01910] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c89] =  If409768b648a33a7ed878a070d4f6251['h01912] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c8a] =  If409768b648a33a7ed878a070d4f6251['h01914] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c8b] =  If409768b648a33a7ed878a070d4f6251['h01916] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c8c] =  If409768b648a33a7ed878a070d4f6251['h01918] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c8d] =  If409768b648a33a7ed878a070d4f6251['h0191a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c8e] =  If409768b648a33a7ed878a070d4f6251['h0191c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c8f] =  If409768b648a33a7ed878a070d4f6251['h0191e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c90] =  If409768b648a33a7ed878a070d4f6251['h01920] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c91] =  If409768b648a33a7ed878a070d4f6251['h01922] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c92] =  If409768b648a33a7ed878a070d4f6251['h01924] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c93] =  If409768b648a33a7ed878a070d4f6251['h01926] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c94] =  If409768b648a33a7ed878a070d4f6251['h01928] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c95] =  If409768b648a33a7ed878a070d4f6251['h0192a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c96] =  If409768b648a33a7ed878a070d4f6251['h0192c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c97] =  If409768b648a33a7ed878a070d4f6251['h0192e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c98] =  If409768b648a33a7ed878a070d4f6251['h01930] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c99] =  If409768b648a33a7ed878a070d4f6251['h01932] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c9a] =  If409768b648a33a7ed878a070d4f6251['h01934] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c9b] =  If409768b648a33a7ed878a070d4f6251['h01936] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c9c] =  If409768b648a33a7ed878a070d4f6251['h01938] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c9d] =  If409768b648a33a7ed878a070d4f6251['h0193a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c9e] =  If409768b648a33a7ed878a070d4f6251['h0193c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00c9f] =  If409768b648a33a7ed878a070d4f6251['h0193e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ca0] =  If409768b648a33a7ed878a070d4f6251['h01940] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ca1] =  If409768b648a33a7ed878a070d4f6251['h01942] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ca2] =  If409768b648a33a7ed878a070d4f6251['h01944] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ca3] =  If409768b648a33a7ed878a070d4f6251['h01946] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ca4] =  If409768b648a33a7ed878a070d4f6251['h01948] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ca5] =  If409768b648a33a7ed878a070d4f6251['h0194a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ca6] =  If409768b648a33a7ed878a070d4f6251['h0194c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ca7] =  If409768b648a33a7ed878a070d4f6251['h0194e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ca8] =  If409768b648a33a7ed878a070d4f6251['h01950] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ca9] =  If409768b648a33a7ed878a070d4f6251['h01952] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00caa] =  If409768b648a33a7ed878a070d4f6251['h01954] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cab] =  If409768b648a33a7ed878a070d4f6251['h01956] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cac] =  If409768b648a33a7ed878a070d4f6251['h01958] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cad] =  If409768b648a33a7ed878a070d4f6251['h0195a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cae] =  If409768b648a33a7ed878a070d4f6251['h0195c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00caf] =  If409768b648a33a7ed878a070d4f6251['h0195e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cb0] =  If409768b648a33a7ed878a070d4f6251['h01960] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cb1] =  If409768b648a33a7ed878a070d4f6251['h01962] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cb2] =  If409768b648a33a7ed878a070d4f6251['h01964] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cb3] =  If409768b648a33a7ed878a070d4f6251['h01966] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cb4] =  If409768b648a33a7ed878a070d4f6251['h01968] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cb5] =  If409768b648a33a7ed878a070d4f6251['h0196a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cb6] =  If409768b648a33a7ed878a070d4f6251['h0196c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cb7] =  If409768b648a33a7ed878a070d4f6251['h0196e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cb8] =  If409768b648a33a7ed878a070d4f6251['h01970] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cb9] =  If409768b648a33a7ed878a070d4f6251['h01972] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cba] =  If409768b648a33a7ed878a070d4f6251['h01974] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cbb] =  If409768b648a33a7ed878a070d4f6251['h01976] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cbc] =  If409768b648a33a7ed878a070d4f6251['h01978] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cbd] =  If409768b648a33a7ed878a070d4f6251['h0197a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cbe] =  If409768b648a33a7ed878a070d4f6251['h0197c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cbf] =  If409768b648a33a7ed878a070d4f6251['h0197e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cc0] =  If409768b648a33a7ed878a070d4f6251['h01980] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cc1] =  If409768b648a33a7ed878a070d4f6251['h01982] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cc2] =  If409768b648a33a7ed878a070d4f6251['h01984] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cc3] =  If409768b648a33a7ed878a070d4f6251['h01986] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cc4] =  If409768b648a33a7ed878a070d4f6251['h01988] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cc5] =  If409768b648a33a7ed878a070d4f6251['h0198a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cc6] =  If409768b648a33a7ed878a070d4f6251['h0198c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cc7] =  If409768b648a33a7ed878a070d4f6251['h0198e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cc8] =  If409768b648a33a7ed878a070d4f6251['h01990] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cc9] =  If409768b648a33a7ed878a070d4f6251['h01992] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cca] =  If409768b648a33a7ed878a070d4f6251['h01994] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ccb] =  If409768b648a33a7ed878a070d4f6251['h01996] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ccc] =  If409768b648a33a7ed878a070d4f6251['h01998] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ccd] =  If409768b648a33a7ed878a070d4f6251['h0199a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cce] =  If409768b648a33a7ed878a070d4f6251['h0199c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ccf] =  If409768b648a33a7ed878a070d4f6251['h0199e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cd0] =  If409768b648a33a7ed878a070d4f6251['h019a0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cd1] =  If409768b648a33a7ed878a070d4f6251['h019a2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cd2] =  If409768b648a33a7ed878a070d4f6251['h019a4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cd3] =  If409768b648a33a7ed878a070d4f6251['h019a6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cd4] =  If409768b648a33a7ed878a070d4f6251['h019a8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cd5] =  If409768b648a33a7ed878a070d4f6251['h019aa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cd6] =  If409768b648a33a7ed878a070d4f6251['h019ac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cd7] =  If409768b648a33a7ed878a070d4f6251['h019ae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cd8] =  If409768b648a33a7ed878a070d4f6251['h019b0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cd9] =  If409768b648a33a7ed878a070d4f6251['h019b2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cda] =  If409768b648a33a7ed878a070d4f6251['h019b4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cdb] =  If409768b648a33a7ed878a070d4f6251['h019b6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cdc] =  If409768b648a33a7ed878a070d4f6251['h019b8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cdd] =  If409768b648a33a7ed878a070d4f6251['h019ba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cde] =  If409768b648a33a7ed878a070d4f6251['h019bc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cdf] =  If409768b648a33a7ed878a070d4f6251['h019be] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ce0] =  If409768b648a33a7ed878a070d4f6251['h019c0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ce1] =  If409768b648a33a7ed878a070d4f6251['h019c2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ce2] =  If409768b648a33a7ed878a070d4f6251['h019c4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ce3] =  If409768b648a33a7ed878a070d4f6251['h019c6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ce4] =  If409768b648a33a7ed878a070d4f6251['h019c8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ce5] =  If409768b648a33a7ed878a070d4f6251['h019ca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ce6] =  If409768b648a33a7ed878a070d4f6251['h019cc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ce7] =  If409768b648a33a7ed878a070d4f6251['h019ce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ce8] =  If409768b648a33a7ed878a070d4f6251['h019d0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ce9] =  If409768b648a33a7ed878a070d4f6251['h019d2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cea] =  If409768b648a33a7ed878a070d4f6251['h019d4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ceb] =  If409768b648a33a7ed878a070d4f6251['h019d6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cec] =  If409768b648a33a7ed878a070d4f6251['h019d8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ced] =  If409768b648a33a7ed878a070d4f6251['h019da] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cee] =  If409768b648a33a7ed878a070d4f6251['h019dc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cef] =  If409768b648a33a7ed878a070d4f6251['h019de] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cf0] =  If409768b648a33a7ed878a070d4f6251['h019e0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cf1] =  If409768b648a33a7ed878a070d4f6251['h019e2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cf2] =  If409768b648a33a7ed878a070d4f6251['h019e4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cf3] =  If409768b648a33a7ed878a070d4f6251['h019e6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cf4] =  If409768b648a33a7ed878a070d4f6251['h019e8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cf5] =  If409768b648a33a7ed878a070d4f6251['h019ea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cf6] =  If409768b648a33a7ed878a070d4f6251['h019ec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cf7] =  If409768b648a33a7ed878a070d4f6251['h019ee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cf8] =  If409768b648a33a7ed878a070d4f6251['h019f0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cf9] =  If409768b648a33a7ed878a070d4f6251['h019f2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cfa] =  If409768b648a33a7ed878a070d4f6251['h019f4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cfb] =  If409768b648a33a7ed878a070d4f6251['h019f6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cfc] =  If409768b648a33a7ed878a070d4f6251['h019f8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cfd] =  If409768b648a33a7ed878a070d4f6251['h019fa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cfe] =  If409768b648a33a7ed878a070d4f6251['h019fc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00cff] =  If409768b648a33a7ed878a070d4f6251['h019fe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d00] =  If409768b648a33a7ed878a070d4f6251['h01a00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d01] =  If409768b648a33a7ed878a070d4f6251['h01a02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d02] =  If409768b648a33a7ed878a070d4f6251['h01a04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d03] =  If409768b648a33a7ed878a070d4f6251['h01a06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d04] =  If409768b648a33a7ed878a070d4f6251['h01a08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d05] =  If409768b648a33a7ed878a070d4f6251['h01a0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d06] =  If409768b648a33a7ed878a070d4f6251['h01a0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d07] =  If409768b648a33a7ed878a070d4f6251['h01a0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d08] =  If409768b648a33a7ed878a070d4f6251['h01a10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d09] =  If409768b648a33a7ed878a070d4f6251['h01a12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d0a] =  If409768b648a33a7ed878a070d4f6251['h01a14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d0b] =  If409768b648a33a7ed878a070d4f6251['h01a16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d0c] =  If409768b648a33a7ed878a070d4f6251['h01a18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d0d] =  If409768b648a33a7ed878a070d4f6251['h01a1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d0e] =  If409768b648a33a7ed878a070d4f6251['h01a1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d0f] =  If409768b648a33a7ed878a070d4f6251['h01a1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d10] =  If409768b648a33a7ed878a070d4f6251['h01a20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d11] =  If409768b648a33a7ed878a070d4f6251['h01a22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d12] =  If409768b648a33a7ed878a070d4f6251['h01a24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d13] =  If409768b648a33a7ed878a070d4f6251['h01a26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d14] =  If409768b648a33a7ed878a070d4f6251['h01a28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d15] =  If409768b648a33a7ed878a070d4f6251['h01a2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d16] =  If409768b648a33a7ed878a070d4f6251['h01a2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d17] =  If409768b648a33a7ed878a070d4f6251['h01a2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d18] =  If409768b648a33a7ed878a070d4f6251['h01a30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d19] =  If409768b648a33a7ed878a070d4f6251['h01a32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d1a] =  If409768b648a33a7ed878a070d4f6251['h01a34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d1b] =  If409768b648a33a7ed878a070d4f6251['h01a36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d1c] =  If409768b648a33a7ed878a070d4f6251['h01a38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d1d] =  If409768b648a33a7ed878a070d4f6251['h01a3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d1e] =  If409768b648a33a7ed878a070d4f6251['h01a3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d1f] =  If409768b648a33a7ed878a070d4f6251['h01a3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d20] =  If409768b648a33a7ed878a070d4f6251['h01a40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d21] =  If409768b648a33a7ed878a070d4f6251['h01a42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d22] =  If409768b648a33a7ed878a070d4f6251['h01a44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d23] =  If409768b648a33a7ed878a070d4f6251['h01a46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d24] =  If409768b648a33a7ed878a070d4f6251['h01a48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d25] =  If409768b648a33a7ed878a070d4f6251['h01a4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d26] =  If409768b648a33a7ed878a070d4f6251['h01a4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d27] =  If409768b648a33a7ed878a070d4f6251['h01a4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d28] =  If409768b648a33a7ed878a070d4f6251['h01a50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d29] =  If409768b648a33a7ed878a070d4f6251['h01a52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d2a] =  If409768b648a33a7ed878a070d4f6251['h01a54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d2b] =  If409768b648a33a7ed878a070d4f6251['h01a56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d2c] =  If409768b648a33a7ed878a070d4f6251['h01a58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d2d] =  If409768b648a33a7ed878a070d4f6251['h01a5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d2e] =  If409768b648a33a7ed878a070d4f6251['h01a5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d2f] =  If409768b648a33a7ed878a070d4f6251['h01a5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d30] =  If409768b648a33a7ed878a070d4f6251['h01a60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d31] =  If409768b648a33a7ed878a070d4f6251['h01a62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d32] =  If409768b648a33a7ed878a070d4f6251['h01a64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d33] =  If409768b648a33a7ed878a070d4f6251['h01a66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d34] =  If409768b648a33a7ed878a070d4f6251['h01a68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d35] =  If409768b648a33a7ed878a070d4f6251['h01a6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d36] =  If409768b648a33a7ed878a070d4f6251['h01a6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d37] =  If409768b648a33a7ed878a070d4f6251['h01a6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d38] =  If409768b648a33a7ed878a070d4f6251['h01a70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d39] =  If409768b648a33a7ed878a070d4f6251['h01a72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d3a] =  If409768b648a33a7ed878a070d4f6251['h01a74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d3b] =  If409768b648a33a7ed878a070d4f6251['h01a76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d3c] =  If409768b648a33a7ed878a070d4f6251['h01a78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d3d] =  If409768b648a33a7ed878a070d4f6251['h01a7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d3e] =  If409768b648a33a7ed878a070d4f6251['h01a7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d3f] =  If409768b648a33a7ed878a070d4f6251['h01a7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d40] =  If409768b648a33a7ed878a070d4f6251['h01a80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d41] =  If409768b648a33a7ed878a070d4f6251['h01a82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d42] =  If409768b648a33a7ed878a070d4f6251['h01a84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d43] =  If409768b648a33a7ed878a070d4f6251['h01a86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d44] =  If409768b648a33a7ed878a070d4f6251['h01a88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d45] =  If409768b648a33a7ed878a070d4f6251['h01a8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d46] =  If409768b648a33a7ed878a070d4f6251['h01a8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d47] =  If409768b648a33a7ed878a070d4f6251['h01a8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d48] =  If409768b648a33a7ed878a070d4f6251['h01a90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d49] =  If409768b648a33a7ed878a070d4f6251['h01a92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d4a] =  If409768b648a33a7ed878a070d4f6251['h01a94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d4b] =  If409768b648a33a7ed878a070d4f6251['h01a96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d4c] =  If409768b648a33a7ed878a070d4f6251['h01a98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d4d] =  If409768b648a33a7ed878a070d4f6251['h01a9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d4e] =  If409768b648a33a7ed878a070d4f6251['h01a9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d4f] =  If409768b648a33a7ed878a070d4f6251['h01a9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d50] =  If409768b648a33a7ed878a070d4f6251['h01aa0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d51] =  If409768b648a33a7ed878a070d4f6251['h01aa2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d52] =  If409768b648a33a7ed878a070d4f6251['h01aa4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d53] =  If409768b648a33a7ed878a070d4f6251['h01aa6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d54] =  If409768b648a33a7ed878a070d4f6251['h01aa8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d55] =  If409768b648a33a7ed878a070d4f6251['h01aaa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d56] =  If409768b648a33a7ed878a070d4f6251['h01aac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d57] =  If409768b648a33a7ed878a070d4f6251['h01aae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d58] =  If409768b648a33a7ed878a070d4f6251['h01ab0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d59] =  If409768b648a33a7ed878a070d4f6251['h01ab2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d5a] =  If409768b648a33a7ed878a070d4f6251['h01ab4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d5b] =  If409768b648a33a7ed878a070d4f6251['h01ab6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d5c] =  If409768b648a33a7ed878a070d4f6251['h01ab8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d5d] =  If409768b648a33a7ed878a070d4f6251['h01aba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d5e] =  If409768b648a33a7ed878a070d4f6251['h01abc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d5f] =  If409768b648a33a7ed878a070d4f6251['h01abe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d60] =  If409768b648a33a7ed878a070d4f6251['h01ac0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d61] =  If409768b648a33a7ed878a070d4f6251['h01ac2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d62] =  If409768b648a33a7ed878a070d4f6251['h01ac4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d63] =  If409768b648a33a7ed878a070d4f6251['h01ac6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d64] =  If409768b648a33a7ed878a070d4f6251['h01ac8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d65] =  If409768b648a33a7ed878a070d4f6251['h01aca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d66] =  If409768b648a33a7ed878a070d4f6251['h01acc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d67] =  If409768b648a33a7ed878a070d4f6251['h01ace] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d68] =  If409768b648a33a7ed878a070d4f6251['h01ad0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d69] =  If409768b648a33a7ed878a070d4f6251['h01ad2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d6a] =  If409768b648a33a7ed878a070d4f6251['h01ad4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d6b] =  If409768b648a33a7ed878a070d4f6251['h01ad6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d6c] =  If409768b648a33a7ed878a070d4f6251['h01ad8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d6d] =  If409768b648a33a7ed878a070d4f6251['h01ada] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d6e] =  If409768b648a33a7ed878a070d4f6251['h01adc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d6f] =  If409768b648a33a7ed878a070d4f6251['h01ade] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d70] =  If409768b648a33a7ed878a070d4f6251['h01ae0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d71] =  If409768b648a33a7ed878a070d4f6251['h01ae2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d72] =  If409768b648a33a7ed878a070d4f6251['h01ae4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d73] =  If409768b648a33a7ed878a070d4f6251['h01ae6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d74] =  If409768b648a33a7ed878a070d4f6251['h01ae8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d75] =  If409768b648a33a7ed878a070d4f6251['h01aea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d76] =  If409768b648a33a7ed878a070d4f6251['h01aec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d77] =  If409768b648a33a7ed878a070d4f6251['h01aee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d78] =  If409768b648a33a7ed878a070d4f6251['h01af0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d79] =  If409768b648a33a7ed878a070d4f6251['h01af2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d7a] =  If409768b648a33a7ed878a070d4f6251['h01af4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d7b] =  If409768b648a33a7ed878a070d4f6251['h01af6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d7c] =  If409768b648a33a7ed878a070d4f6251['h01af8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d7d] =  If409768b648a33a7ed878a070d4f6251['h01afa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d7e] =  If409768b648a33a7ed878a070d4f6251['h01afc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d7f] =  If409768b648a33a7ed878a070d4f6251['h01afe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d80] =  If409768b648a33a7ed878a070d4f6251['h01b00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d81] =  If409768b648a33a7ed878a070d4f6251['h01b02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d82] =  If409768b648a33a7ed878a070d4f6251['h01b04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d83] =  If409768b648a33a7ed878a070d4f6251['h01b06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d84] =  If409768b648a33a7ed878a070d4f6251['h01b08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d85] =  If409768b648a33a7ed878a070d4f6251['h01b0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d86] =  If409768b648a33a7ed878a070d4f6251['h01b0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d87] =  If409768b648a33a7ed878a070d4f6251['h01b0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d88] =  If409768b648a33a7ed878a070d4f6251['h01b10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d89] =  If409768b648a33a7ed878a070d4f6251['h01b12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d8a] =  If409768b648a33a7ed878a070d4f6251['h01b14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d8b] =  If409768b648a33a7ed878a070d4f6251['h01b16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d8c] =  If409768b648a33a7ed878a070d4f6251['h01b18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d8d] =  If409768b648a33a7ed878a070d4f6251['h01b1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d8e] =  If409768b648a33a7ed878a070d4f6251['h01b1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d8f] =  If409768b648a33a7ed878a070d4f6251['h01b1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d90] =  If409768b648a33a7ed878a070d4f6251['h01b20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d91] =  If409768b648a33a7ed878a070d4f6251['h01b22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d92] =  If409768b648a33a7ed878a070d4f6251['h01b24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d93] =  If409768b648a33a7ed878a070d4f6251['h01b26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d94] =  If409768b648a33a7ed878a070d4f6251['h01b28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d95] =  If409768b648a33a7ed878a070d4f6251['h01b2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d96] =  If409768b648a33a7ed878a070d4f6251['h01b2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d97] =  If409768b648a33a7ed878a070d4f6251['h01b2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d98] =  If409768b648a33a7ed878a070d4f6251['h01b30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d99] =  If409768b648a33a7ed878a070d4f6251['h01b32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d9a] =  If409768b648a33a7ed878a070d4f6251['h01b34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d9b] =  If409768b648a33a7ed878a070d4f6251['h01b36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d9c] =  If409768b648a33a7ed878a070d4f6251['h01b38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d9d] =  If409768b648a33a7ed878a070d4f6251['h01b3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d9e] =  If409768b648a33a7ed878a070d4f6251['h01b3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00d9f] =  If409768b648a33a7ed878a070d4f6251['h01b3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00da0] =  If409768b648a33a7ed878a070d4f6251['h01b40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00da1] =  If409768b648a33a7ed878a070d4f6251['h01b42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00da2] =  If409768b648a33a7ed878a070d4f6251['h01b44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00da3] =  If409768b648a33a7ed878a070d4f6251['h01b46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00da4] =  If409768b648a33a7ed878a070d4f6251['h01b48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00da5] =  If409768b648a33a7ed878a070d4f6251['h01b4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00da6] =  If409768b648a33a7ed878a070d4f6251['h01b4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00da7] =  If409768b648a33a7ed878a070d4f6251['h01b4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00da8] =  If409768b648a33a7ed878a070d4f6251['h01b50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00da9] =  If409768b648a33a7ed878a070d4f6251['h01b52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00daa] =  If409768b648a33a7ed878a070d4f6251['h01b54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dab] =  If409768b648a33a7ed878a070d4f6251['h01b56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dac] =  If409768b648a33a7ed878a070d4f6251['h01b58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dad] =  If409768b648a33a7ed878a070d4f6251['h01b5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dae] =  If409768b648a33a7ed878a070d4f6251['h01b5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00daf] =  If409768b648a33a7ed878a070d4f6251['h01b5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00db0] =  If409768b648a33a7ed878a070d4f6251['h01b60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00db1] =  If409768b648a33a7ed878a070d4f6251['h01b62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00db2] =  If409768b648a33a7ed878a070d4f6251['h01b64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00db3] =  If409768b648a33a7ed878a070d4f6251['h01b66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00db4] =  If409768b648a33a7ed878a070d4f6251['h01b68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00db5] =  If409768b648a33a7ed878a070d4f6251['h01b6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00db6] =  If409768b648a33a7ed878a070d4f6251['h01b6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00db7] =  If409768b648a33a7ed878a070d4f6251['h01b6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00db8] =  If409768b648a33a7ed878a070d4f6251['h01b70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00db9] =  If409768b648a33a7ed878a070d4f6251['h01b72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dba] =  If409768b648a33a7ed878a070d4f6251['h01b74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dbb] =  If409768b648a33a7ed878a070d4f6251['h01b76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dbc] =  If409768b648a33a7ed878a070d4f6251['h01b78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dbd] =  If409768b648a33a7ed878a070d4f6251['h01b7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dbe] =  If409768b648a33a7ed878a070d4f6251['h01b7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dbf] =  If409768b648a33a7ed878a070d4f6251['h01b7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dc0] =  If409768b648a33a7ed878a070d4f6251['h01b80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dc1] =  If409768b648a33a7ed878a070d4f6251['h01b82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dc2] =  If409768b648a33a7ed878a070d4f6251['h01b84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dc3] =  If409768b648a33a7ed878a070d4f6251['h01b86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dc4] =  If409768b648a33a7ed878a070d4f6251['h01b88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dc5] =  If409768b648a33a7ed878a070d4f6251['h01b8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dc6] =  If409768b648a33a7ed878a070d4f6251['h01b8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dc7] =  If409768b648a33a7ed878a070d4f6251['h01b8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dc8] =  If409768b648a33a7ed878a070d4f6251['h01b90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dc9] =  If409768b648a33a7ed878a070d4f6251['h01b92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dca] =  If409768b648a33a7ed878a070d4f6251['h01b94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dcb] =  If409768b648a33a7ed878a070d4f6251['h01b96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dcc] =  If409768b648a33a7ed878a070d4f6251['h01b98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dcd] =  If409768b648a33a7ed878a070d4f6251['h01b9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dce] =  If409768b648a33a7ed878a070d4f6251['h01b9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dcf] =  If409768b648a33a7ed878a070d4f6251['h01b9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dd0] =  If409768b648a33a7ed878a070d4f6251['h01ba0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dd1] =  If409768b648a33a7ed878a070d4f6251['h01ba2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dd2] =  If409768b648a33a7ed878a070d4f6251['h01ba4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dd3] =  If409768b648a33a7ed878a070d4f6251['h01ba6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dd4] =  If409768b648a33a7ed878a070d4f6251['h01ba8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dd5] =  If409768b648a33a7ed878a070d4f6251['h01baa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dd6] =  If409768b648a33a7ed878a070d4f6251['h01bac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dd7] =  If409768b648a33a7ed878a070d4f6251['h01bae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dd8] =  If409768b648a33a7ed878a070d4f6251['h01bb0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dd9] =  If409768b648a33a7ed878a070d4f6251['h01bb2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dda] =  If409768b648a33a7ed878a070d4f6251['h01bb4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ddb] =  If409768b648a33a7ed878a070d4f6251['h01bb6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ddc] =  If409768b648a33a7ed878a070d4f6251['h01bb8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ddd] =  If409768b648a33a7ed878a070d4f6251['h01bba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dde] =  If409768b648a33a7ed878a070d4f6251['h01bbc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ddf] =  If409768b648a33a7ed878a070d4f6251['h01bbe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00de0] =  If409768b648a33a7ed878a070d4f6251['h01bc0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00de1] =  If409768b648a33a7ed878a070d4f6251['h01bc2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00de2] =  If409768b648a33a7ed878a070d4f6251['h01bc4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00de3] =  If409768b648a33a7ed878a070d4f6251['h01bc6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00de4] =  If409768b648a33a7ed878a070d4f6251['h01bc8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00de5] =  If409768b648a33a7ed878a070d4f6251['h01bca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00de6] =  If409768b648a33a7ed878a070d4f6251['h01bcc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00de7] =  If409768b648a33a7ed878a070d4f6251['h01bce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00de8] =  If409768b648a33a7ed878a070d4f6251['h01bd0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00de9] =  If409768b648a33a7ed878a070d4f6251['h01bd2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dea] =  If409768b648a33a7ed878a070d4f6251['h01bd4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00deb] =  If409768b648a33a7ed878a070d4f6251['h01bd6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dec] =  If409768b648a33a7ed878a070d4f6251['h01bd8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ded] =  If409768b648a33a7ed878a070d4f6251['h01bda] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dee] =  If409768b648a33a7ed878a070d4f6251['h01bdc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00def] =  If409768b648a33a7ed878a070d4f6251['h01bde] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00df0] =  If409768b648a33a7ed878a070d4f6251['h01be0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00df1] =  If409768b648a33a7ed878a070d4f6251['h01be2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00df2] =  If409768b648a33a7ed878a070d4f6251['h01be4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00df3] =  If409768b648a33a7ed878a070d4f6251['h01be6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00df4] =  If409768b648a33a7ed878a070d4f6251['h01be8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00df5] =  If409768b648a33a7ed878a070d4f6251['h01bea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00df6] =  If409768b648a33a7ed878a070d4f6251['h01bec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00df7] =  If409768b648a33a7ed878a070d4f6251['h01bee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00df8] =  If409768b648a33a7ed878a070d4f6251['h01bf0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00df9] =  If409768b648a33a7ed878a070d4f6251['h01bf2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dfa] =  If409768b648a33a7ed878a070d4f6251['h01bf4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dfb] =  If409768b648a33a7ed878a070d4f6251['h01bf6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dfc] =  If409768b648a33a7ed878a070d4f6251['h01bf8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dfd] =  If409768b648a33a7ed878a070d4f6251['h01bfa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dfe] =  If409768b648a33a7ed878a070d4f6251['h01bfc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00dff] =  If409768b648a33a7ed878a070d4f6251['h01bfe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e00] =  If409768b648a33a7ed878a070d4f6251['h01c00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e01] =  If409768b648a33a7ed878a070d4f6251['h01c02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e02] =  If409768b648a33a7ed878a070d4f6251['h01c04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e03] =  If409768b648a33a7ed878a070d4f6251['h01c06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e04] =  If409768b648a33a7ed878a070d4f6251['h01c08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e05] =  If409768b648a33a7ed878a070d4f6251['h01c0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e06] =  If409768b648a33a7ed878a070d4f6251['h01c0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e07] =  If409768b648a33a7ed878a070d4f6251['h01c0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e08] =  If409768b648a33a7ed878a070d4f6251['h01c10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e09] =  If409768b648a33a7ed878a070d4f6251['h01c12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e0a] =  If409768b648a33a7ed878a070d4f6251['h01c14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e0b] =  If409768b648a33a7ed878a070d4f6251['h01c16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e0c] =  If409768b648a33a7ed878a070d4f6251['h01c18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e0d] =  If409768b648a33a7ed878a070d4f6251['h01c1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e0e] =  If409768b648a33a7ed878a070d4f6251['h01c1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e0f] =  If409768b648a33a7ed878a070d4f6251['h01c1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e10] =  If409768b648a33a7ed878a070d4f6251['h01c20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e11] =  If409768b648a33a7ed878a070d4f6251['h01c22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e12] =  If409768b648a33a7ed878a070d4f6251['h01c24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e13] =  If409768b648a33a7ed878a070d4f6251['h01c26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e14] =  If409768b648a33a7ed878a070d4f6251['h01c28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e15] =  If409768b648a33a7ed878a070d4f6251['h01c2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e16] =  If409768b648a33a7ed878a070d4f6251['h01c2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e17] =  If409768b648a33a7ed878a070d4f6251['h01c2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e18] =  If409768b648a33a7ed878a070d4f6251['h01c30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e19] =  If409768b648a33a7ed878a070d4f6251['h01c32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e1a] =  If409768b648a33a7ed878a070d4f6251['h01c34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e1b] =  If409768b648a33a7ed878a070d4f6251['h01c36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e1c] =  If409768b648a33a7ed878a070d4f6251['h01c38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e1d] =  If409768b648a33a7ed878a070d4f6251['h01c3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e1e] =  If409768b648a33a7ed878a070d4f6251['h01c3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e1f] =  If409768b648a33a7ed878a070d4f6251['h01c3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e20] =  If409768b648a33a7ed878a070d4f6251['h01c40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e21] =  If409768b648a33a7ed878a070d4f6251['h01c42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e22] =  If409768b648a33a7ed878a070d4f6251['h01c44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e23] =  If409768b648a33a7ed878a070d4f6251['h01c46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e24] =  If409768b648a33a7ed878a070d4f6251['h01c48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e25] =  If409768b648a33a7ed878a070d4f6251['h01c4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e26] =  If409768b648a33a7ed878a070d4f6251['h01c4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e27] =  If409768b648a33a7ed878a070d4f6251['h01c4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e28] =  If409768b648a33a7ed878a070d4f6251['h01c50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e29] =  If409768b648a33a7ed878a070d4f6251['h01c52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e2a] =  If409768b648a33a7ed878a070d4f6251['h01c54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e2b] =  If409768b648a33a7ed878a070d4f6251['h01c56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e2c] =  If409768b648a33a7ed878a070d4f6251['h01c58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e2d] =  If409768b648a33a7ed878a070d4f6251['h01c5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e2e] =  If409768b648a33a7ed878a070d4f6251['h01c5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e2f] =  If409768b648a33a7ed878a070d4f6251['h01c5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e30] =  If409768b648a33a7ed878a070d4f6251['h01c60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e31] =  If409768b648a33a7ed878a070d4f6251['h01c62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e32] =  If409768b648a33a7ed878a070d4f6251['h01c64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e33] =  If409768b648a33a7ed878a070d4f6251['h01c66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e34] =  If409768b648a33a7ed878a070d4f6251['h01c68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e35] =  If409768b648a33a7ed878a070d4f6251['h01c6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e36] =  If409768b648a33a7ed878a070d4f6251['h01c6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e37] =  If409768b648a33a7ed878a070d4f6251['h01c6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e38] =  If409768b648a33a7ed878a070d4f6251['h01c70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e39] =  If409768b648a33a7ed878a070d4f6251['h01c72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e3a] =  If409768b648a33a7ed878a070d4f6251['h01c74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e3b] =  If409768b648a33a7ed878a070d4f6251['h01c76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e3c] =  If409768b648a33a7ed878a070d4f6251['h01c78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e3d] =  If409768b648a33a7ed878a070d4f6251['h01c7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e3e] =  If409768b648a33a7ed878a070d4f6251['h01c7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e3f] =  If409768b648a33a7ed878a070d4f6251['h01c7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e40] =  If409768b648a33a7ed878a070d4f6251['h01c80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e41] =  If409768b648a33a7ed878a070d4f6251['h01c82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e42] =  If409768b648a33a7ed878a070d4f6251['h01c84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e43] =  If409768b648a33a7ed878a070d4f6251['h01c86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e44] =  If409768b648a33a7ed878a070d4f6251['h01c88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e45] =  If409768b648a33a7ed878a070d4f6251['h01c8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e46] =  If409768b648a33a7ed878a070d4f6251['h01c8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e47] =  If409768b648a33a7ed878a070d4f6251['h01c8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e48] =  If409768b648a33a7ed878a070d4f6251['h01c90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e49] =  If409768b648a33a7ed878a070d4f6251['h01c92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e4a] =  If409768b648a33a7ed878a070d4f6251['h01c94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e4b] =  If409768b648a33a7ed878a070d4f6251['h01c96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e4c] =  If409768b648a33a7ed878a070d4f6251['h01c98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e4d] =  If409768b648a33a7ed878a070d4f6251['h01c9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e4e] =  If409768b648a33a7ed878a070d4f6251['h01c9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e4f] =  If409768b648a33a7ed878a070d4f6251['h01c9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e50] =  If409768b648a33a7ed878a070d4f6251['h01ca0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e51] =  If409768b648a33a7ed878a070d4f6251['h01ca2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e52] =  If409768b648a33a7ed878a070d4f6251['h01ca4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e53] =  If409768b648a33a7ed878a070d4f6251['h01ca6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e54] =  If409768b648a33a7ed878a070d4f6251['h01ca8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e55] =  If409768b648a33a7ed878a070d4f6251['h01caa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e56] =  If409768b648a33a7ed878a070d4f6251['h01cac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e57] =  If409768b648a33a7ed878a070d4f6251['h01cae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e58] =  If409768b648a33a7ed878a070d4f6251['h01cb0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e59] =  If409768b648a33a7ed878a070d4f6251['h01cb2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e5a] =  If409768b648a33a7ed878a070d4f6251['h01cb4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e5b] =  If409768b648a33a7ed878a070d4f6251['h01cb6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e5c] =  If409768b648a33a7ed878a070d4f6251['h01cb8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e5d] =  If409768b648a33a7ed878a070d4f6251['h01cba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e5e] =  If409768b648a33a7ed878a070d4f6251['h01cbc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e5f] =  If409768b648a33a7ed878a070d4f6251['h01cbe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e60] =  If409768b648a33a7ed878a070d4f6251['h01cc0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e61] =  If409768b648a33a7ed878a070d4f6251['h01cc2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e62] =  If409768b648a33a7ed878a070d4f6251['h01cc4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e63] =  If409768b648a33a7ed878a070d4f6251['h01cc6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e64] =  If409768b648a33a7ed878a070d4f6251['h01cc8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e65] =  If409768b648a33a7ed878a070d4f6251['h01cca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e66] =  If409768b648a33a7ed878a070d4f6251['h01ccc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e67] =  If409768b648a33a7ed878a070d4f6251['h01cce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e68] =  If409768b648a33a7ed878a070d4f6251['h01cd0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e69] =  If409768b648a33a7ed878a070d4f6251['h01cd2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e6a] =  If409768b648a33a7ed878a070d4f6251['h01cd4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e6b] =  If409768b648a33a7ed878a070d4f6251['h01cd6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e6c] =  If409768b648a33a7ed878a070d4f6251['h01cd8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e6d] =  If409768b648a33a7ed878a070d4f6251['h01cda] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e6e] =  If409768b648a33a7ed878a070d4f6251['h01cdc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e6f] =  If409768b648a33a7ed878a070d4f6251['h01cde] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e70] =  If409768b648a33a7ed878a070d4f6251['h01ce0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e71] =  If409768b648a33a7ed878a070d4f6251['h01ce2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e72] =  If409768b648a33a7ed878a070d4f6251['h01ce4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e73] =  If409768b648a33a7ed878a070d4f6251['h01ce6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e74] =  If409768b648a33a7ed878a070d4f6251['h01ce8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e75] =  If409768b648a33a7ed878a070d4f6251['h01cea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e76] =  If409768b648a33a7ed878a070d4f6251['h01cec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e77] =  If409768b648a33a7ed878a070d4f6251['h01cee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e78] =  If409768b648a33a7ed878a070d4f6251['h01cf0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e79] =  If409768b648a33a7ed878a070d4f6251['h01cf2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e7a] =  If409768b648a33a7ed878a070d4f6251['h01cf4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e7b] =  If409768b648a33a7ed878a070d4f6251['h01cf6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e7c] =  If409768b648a33a7ed878a070d4f6251['h01cf8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e7d] =  If409768b648a33a7ed878a070d4f6251['h01cfa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e7e] =  If409768b648a33a7ed878a070d4f6251['h01cfc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e7f] =  If409768b648a33a7ed878a070d4f6251['h01cfe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e80] =  If409768b648a33a7ed878a070d4f6251['h01d00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e81] =  If409768b648a33a7ed878a070d4f6251['h01d02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e82] =  If409768b648a33a7ed878a070d4f6251['h01d04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e83] =  If409768b648a33a7ed878a070d4f6251['h01d06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e84] =  If409768b648a33a7ed878a070d4f6251['h01d08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e85] =  If409768b648a33a7ed878a070d4f6251['h01d0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e86] =  If409768b648a33a7ed878a070d4f6251['h01d0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e87] =  If409768b648a33a7ed878a070d4f6251['h01d0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e88] =  If409768b648a33a7ed878a070d4f6251['h01d10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e89] =  If409768b648a33a7ed878a070d4f6251['h01d12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e8a] =  If409768b648a33a7ed878a070d4f6251['h01d14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e8b] =  If409768b648a33a7ed878a070d4f6251['h01d16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e8c] =  If409768b648a33a7ed878a070d4f6251['h01d18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e8d] =  If409768b648a33a7ed878a070d4f6251['h01d1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e8e] =  If409768b648a33a7ed878a070d4f6251['h01d1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e8f] =  If409768b648a33a7ed878a070d4f6251['h01d1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e90] =  If409768b648a33a7ed878a070d4f6251['h01d20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e91] =  If409768b648a33a7ed878a070d4f6251['h01d22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e92] =  If409768b648a33a7ed878a070d4f6251['h01d24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e93] =  If409768b648a33a7ed878a070d4f6251['h01d26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e94] =  If409768b648a33a7ed878a070d4f6251['h01d28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e95] =  If409768b648a33a7ed878a070d4f6251['h01d2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e96] =  If409768b648a33a7ed878a070d4f6251['h01d2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e97] =  If409768b648a33a7ed878a070d4f6251['h01d2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e98] =  If409768b648a33a7ed878a070d4f6251['h01d30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e99] =  If409768b648a33a7ed878a070d4f6251['h01d32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e9a] =  If409768b648a33a7ed878a070d4f6251['h01d34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e9b] =  If409768b648a33a7ed878a070d4f6251['h01d36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e9c] =  If409768b648a33a7ed878a070d4f6251['h01d38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e9d] =  If409768b648a33a7ed878a070d4f6251['h01d3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e9e] =  If409768b648a33a7ed878a070d4f6251['h01d3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00e9f] =  If409768b648a33a7ed878a070d4f6251['h01d3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ea0] =  If409768b648a33a7ed878a070d4f6251['h01d40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ea1] =  If409768b648a33a7ed878a070d4f6251['h01d42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ea2] =  If409768b648a33a7ed878a070d4f6251['h01d44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ea3] =  If409768b648a33a7ed878a070d4f6251['h01d46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ea4] =  If409768b648a33a7ed878a070d4f6251['h01d48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ea5] =  If409768b648a33a7ed878a070d4f6251['h01d4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ea6] =  If409768b648a33a7ed878a070d4f6251['h01d4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ea7] =  If409768b648a33a7ed878a070d4f6251['h01d4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ea8] =  If409768b648a33a7ed878a070d4f6251['h01d50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ea9] =  If409768b648a33a7ed878a070d4f6251['h01d52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eaa] =  If409768b648a33a7ed878a070d4f6251['h01d54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eab] =  If409768b648a33a7ed878a070d4f6251['h01d56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eac] =  If409768b648a33a7ed878a070d4f6251['h01d58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ead] =  If409768b648a33a7ed878a070d4f6251['h01d5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eae] =  If409768b648a33a7ed878a070d4f6251['h01d5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eaf] =  If409768b648a33a7ed878a070d4f6251['h01d5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eb0] =  If409768b648a33a7ed878a070d4f6251['h01d60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eb1] =  If409768b648a33a7ed878a070d4f6251['h01d62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eb2] =  If409768b648a33a7ed878a070d4f6251['h01d64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eb3] =  If409768b648a33a7ed878a070d4f6251['h01d66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eb4] =  If409768b648a33a7ed878a070d4f6251['h01d68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eb5] =  If409768b648a33a7ed878a070d4f6251['h01d6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eb6] =  If409768b648a33a7ed878a070d4f6251['h01d6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eb7] =  If409768b648a33a7ed878a070d4f6251['h01d6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eb8] =  If409768b648a33a7ed878a070d4f6251['h01d70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eb9] =  If409768b648a33a7ed878a070d4f6251['h01d72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eba] =  If409768b648a33a7ed878a070d4f6251['h01d74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ebb] =  If409768b648a33a7ed878a070d4f6251['h01d76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ebc] =  If409768b648a33a7ed878a070d4f6251['h01d78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ebd] =  If409768b648a33a7ed878a070d4f6251['h01d7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ebe] =  If409768b648a33a7ed878a070d4f6251['h01d7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ebf] =  If409768b648a33a7ed878a070d4f6251['h01d7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ec0] =  If409768b648a33a7ed878a070d4f6251['h01d80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ec1] =  If409768b648a33a7ed878a070d4f6251['h01d82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ec2] =  If409768b648a33a7ed878a070d4f6251['h01d84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ec3] =  If409768b648a33a7ed878a070d4f6251['h01d86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ec4] =  If409768b648a33a7ed878a070d4f6251['h01d88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ec5] =  If409768b648a33a7ed878a070d4f6251['h01d8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ec6] =  If409768b648a33a7ed878a070d4f6251['h01d8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ec7] =  If409768b648a33a7ed878a070d4f6251['h01d8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ec8] =  If409768b648a33a7ed878a070d4f6251['h01d90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ec9] =  If409768b648a33a7ed878a070d4f6251['h01d92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eca] =  If409768b648a33a7ed878a070d4f6251['h01d94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ecb] =  If409768b648a33a7ed878a070d4f6251['h01d96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ecc] =  If409768b648a33a7ed878a070d4f6251['h01d98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ecd] =  If409768b648a33a7ed878a070d4f6251['h01d9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ece] =  If409768b648a33a7ed878a070d4f6251['h01d9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ecf] =  If409768b648a33a7ed878a070d4f6251['h01d9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ed0] =  If409768b648a33a7ed878a070d4f6251['h01da0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ed1] =  If409768b648a33a7ed878a070d4f6251['h01da2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ed2] =  If409768b648a33a7ed878a070d4f6251['h01da4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ed3] =  If409768b648a33a7ed878a070d4f6251['h01da6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ed4] =  If409768b648a33a7ed878a070d4f6251['h01da8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ed5] =  If409768b648a33a7ed878a070d4f6251['h01daa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ed6] =  If409768b648a33a7ed878a070d4f6251['h01dac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ed7] =  If409768b648a33a7ed878a070d4f6251['h01dae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ed8] =  If409768b648a33a7ed878a070d4f6251['h01db0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ed9] =  If409768b648a33a7ed878a070d4f6251['h01db2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eda] =  If409768b648a33a7ed878a070d4f6251['h01db4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00edb] =  If409768b648a33a7ed878a070d4f6251['h01db6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00edc] =  If409768b648a33a7ed878a070d4f6251['h01db8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00edd] =  If409768b648a33a7ed878a070d4f6251['h01dba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ede] =  If409768b648a33a7ed878a070d4f6251['h01dbc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00edf] =  If409768b648a33a7ed878a070d4f6251['h01dbe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ee0] =  If409768b648a33a7ed878a070d4f6251['h01dc0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ee1] =  If409768b648a33a7ed878a070d4f6251['h01dc2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ee2] =  If409768b648a33a7ed878a070d4f6251['h01dc4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ee3] =  If409768b648a33a7ed878a070d4f6251['h01dc6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ee4] =  If409768b648a33a7ed878a070d4f6251['h01dc8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ee5] =  If409768b648a33a7ed878a070d4f6251['h01dca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ee6] =  If409768b648a33a7ed878a070d4f6251['h01dcc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ee7] =  If409768b648a33a7ed878a070d4f6251['h01dce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ee8] =  If409768b648a33a7ed878a070d4f6251['h01dd0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ee9] =  If409768b648a33a7ed878a070d4f6251['h01dd2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eea] =  If409768b648a33a7ed878a070d4f6251['h01dd4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eeb] =  If409768b648a33a7ed878a070d4f6251['h01dd6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eec] =  If409768b648a33a7ed878a070d4f6251['h01dd8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eed] =  If409768b648a33a7ed878a070d4f6251['h01dda] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eee] =  If409768b648a33a7ed878a070d4f6251['h01ddc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eef] =  If409768b648a33a7ed878a070d4f6251['h01dde] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ef0] =  If409768b648a33a7ed878a070d4f6251['h01de0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ef1] =  If409768b648a33a7ed878a070d4f6251['h01de2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ef2] =  If409768b648a33a7ed878a070d4f6251['h01de4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ef3] =  If409768b648a33a7ed878a070d4f6251['h01de6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ef4] =  If409768b648a33a7ed878a070d4f6251['h01de8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ef5] =  If409768b648a33a7ed878a070d4f6251['h01dea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ef6] =  If409768b648a33a7ed878a070d4f6251['h01dec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ef7] =  If409768b648a33a7ed878a070d4f6251['h01dee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ef8] =  If409768b648a33a7ed878a070d4f6251['h01df0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ef9] =  If409768b648a33a7ed878a070d4f6251['h01df2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00efa] =  If409768b648a33a7ed878a070d4f6251['h01df4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00efb] =  If409768b648a33a7ed878a070d4f6251['h01df6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00efc] =  If409768b648a33a7ed878a070d4f6251['h01df8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00efd] =  If409768b648a33a7ed878a070d4f6251['h01dfa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00efe] =  If409768b648a33a7ed878a070d4f6251['h01dfc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00eff] =  If409768b648a33a7ed878a070d4f6251['h01dfe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f00] =  If409768b648a33a7ed878a070d4f6251['h01e00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f01] =  If409768b648a33a7ed878a070d4f6251['h01e02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f02] =  If409768b648a33a7ed878a070d4f6251['h01e04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f03] =  If409768b648a33a7ed878a070d4f6251['h01e06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f04] =  If409768b648a33a7ed878a070d4f6251['h01e08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f05] =  If409768b648a33a7ed878a070d4f6251['h01e0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f06] =  If409768b648a33a7ed878a070d4f6251['h01e0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f07] =  If409768b648a33a7ed878a070d4f6251['h01e0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f08] =  If409768b648a33a7ed878a070d4f6251['h01e10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f09] =  If409768b648a33a7ed878a070d4f6251['h01e12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f0a] =  If409768b648a33a7ed878a070d4f6251['h01e14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f0b] =  If409768b648a33a7ed878a070d4f6251['h01e16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f0c] =  If409768b648a33a7ed878a070d4f6251['h01e18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f0d] =  If409768b648a33a7ed878a070d4f6251['h01e1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f0e] =  If409768b648a33a7ed878a070d4f6251['h01e1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f0f] =  If409768b648a33a7ed878a070d4f6251['h01e1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f10] =  If409768b648a33a7ed878a070d4f6251['h01e20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f11] =  If409768b648a33a7ed878a070d4f6251['h01e22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f12] =  If409768b648a33a7ed878a070d4f6251['h01e24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f13] =  If409768b648a33a7ed878a070d4f6251['h01e26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f14] =  If409768b648a33a7ed878a070d4f6251['h01e28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f15] =  If409768b648a33a7ed878a070d4f6251['h01e2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f16] =  If409768b648a33a7ed878a070d4f6251['h01e2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f17] =  If409768b648a33a7ed878a070d4f6251['h01e2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f18] =  If409768b648a33a7ed878a070d4f6251['h01e30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f19] =  If409768b648a33a7ed878a070d4f6251['h01e32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f1a] =  If409768b648a33a7ed878a070d4f6251['h01e34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f1b] =  If409768b648a33a7ed878a070d4f6251['h01e36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f1c] =  If409768b648a33a7ed878a070d4f6251['h01e38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f1d] =  If409768b648a33a7ed878a070d4f6251['h01e3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f1e] =  If409768b648a33a7ed878a070d4f6251['h01e3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f1f] =  If409768b648a33a7ed878a070d4f6251['h01e3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f20] =  If409768b648a33a7ed878a070d4f6251['h01e40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f21] =  If409768b648a33a7ed878a070d4f6251['h01e42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f22] =  If409768b648a33a7ed878a070d4f6251['h01e44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f23] =  If409768b648a33a7ed878a070d4f6251['h01e46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f24] =  If409768b648a33a7ed878a070d4f6251['h01e48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f25] =  If409768b648a33a7ed878a070d4f6251['h01e4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f26] =  If409768b648a33a7ed878a070d4f6251['h01e4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f27] =  If409768b648a33a7ed878a070d4f6251['h01e4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f28] =  If409768b648a33a7ed878a070d4f6251['h01e50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f29] =  If409768b648a33a7ed878a070d4f6251['h01e52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f2a] =  If409768b648a33a7ed878a070d4f6251['h01e54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f2b] =  If409768b648a33a7ed878a070d4f6251['h01e56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f2c] =  If409768b648a33a7ed878a070d4f6251['h01e58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f2d] =  If409768b648a33a7ed878a070d4f6251['h01e5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f2e] =  If409768b648a33a7ed878a070d4f6251['h01e5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f2f] =  If409768b648a33a7ed878a070d4f6251['h01e5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f30] =  If409768b648a33a7ed878a070d4f6251['h01e60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f31] =  If409768b648a33a7ed878a070d4f6251['h01e62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f32] =  If409768b648a33a7ed878a070d4f6251['h01e64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f33] =  If409768b648a33a7ed878a070d4f6251['h01e66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f34] =  If409768b648a33a7ed878a070d4f6251['h01e68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f35] =  If409768b648a33a7ed878a070d4f6251['h01e6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f36] =  If409768b648a33a7ed878a070d4f6251['h01e6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f37] =  If409768b648a33a7ed878a070d4f6251['h01e6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f38] =  If409768b648a33a7ed878a070d4f6251['h01e70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f39] =  If409768b648a33a7ed878a070d4f6251['h01e72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f3a] =  If409768b648a33a7ed878a070d4f6251['h01e74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f3b] =  If409768b648a33a7ed878a070d4f6251['h01e76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f3c] =  If409768b648a33a7ed878a070d4f6251['h01e78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f3d] =  If409768b648a33a7ed878a070d4f6251['h01e7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f3e] =  If409768b648a33a7ed878a070d4f6251['h01e7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f3f] =  If409768b648a33a7ed878a070d4f6251['h01e7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f40] =  If409768b648a33a7ed878a070d4f6251['h01e80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f41] =  If409768b648a33a7ed878a070d4f6251['h01e82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f42] =  If409768b648a33a7ed878a070d4f6251['h01e84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f43] =  If409768b648a33a7ed878a070d4f6251['h01e86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f44] =  If409768b648a33a7ed878a070d4f6251['h01e88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f45] =  If409768b648a33a7ed878a070d4f6251['h01e8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f46] =  If409768b648a33a7ed878a070d4f6251['h01e8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f47] =  If409768b648a33a7ed878a070d4f6251['h01e8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f48] =  If409768b648a33a7ed878a070d4f6251['h01e90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f49] =  If409768b648a33a7ed878a070d4f6251['h01e92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f4a] =  If409768b648a33a7ed878a070d4f6251['h01e94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f4b] =  If409768b648a33a7ed878a070d4f6251['h01e96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f4c] =  If409768b648a33a7ed878a070d4f6251['h01e98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f4d] =  If409768b648a33a7ed878a070d4f6251['h01e9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f4e] =  If409768b648a33a7ed878a070d4f6251['h01e9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f4f] =  If409768b648a33a7ed878a070d4f6251['h01e9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f50] =  If409768b648a33a7ed878a070d4f6251['h01ea0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f51] =  If409768b648a33a7ed878a070d4f6251['h01ea2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f52] =  If409768b648a33a7ed878a070d4f6251['h01ea4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f53] =  If409768b648a33a7ed878a070d4f6251['h01ea6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f54] =  If409768b648a33a7ed878a070d4f6251['h01ea8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f55] =  If409768b648a33a7ed878a070d4f6251['h01eaa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f56] =  If409768b648a33a7ed878a070d4f6251['h01eac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f57] =  If409768b648a33a7ed878a070d4f6251['h01eae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f58] =  If409768b648a33a7ed878a070d4f6251['h01eb0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f59] =  If409768b648a33a7ed878a070d4f6251['h01eb2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f5a] =  If409768b648a33a7ed878a070d4f6251['h01eb4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f5b] =  If409768b648a33a7ed878a070d4f6251['h01eb6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f5c] =  If409768b648a33a7ed878a070d4f6251['h01eb8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f5d] =  If409768b648a33a7ed878a070d4f6251['h01eba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f5e] =  If409768b648a33a7ed878a070d4f6251['h01ebc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f5f] =  If409768b648a33a7ed878a070d4f6251['h01ebe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f60] =  If409768b648a33a7ed878a070d4f6251['h01ec0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f61] =  If409768b648a33a7ed878a070d4f6251['h01ec2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f62] =  If409768b648a33a7ed878a070d4f6251['h01ec4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f63] =  If409768b648a33a7ed878a070d4f6251['h01ec6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f64] =  If409768b648a33a7ed878a070d4f6251['h01ec8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f65] =  If409768b648a33a7ed878a070d4f6251['h01eca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f66] =  If409768b648a33a7ed878a070d4f6251['h01ecc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f67] =  If409768b648a33a7ed878a070d4f6251['h01ece] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f68] =  If409768b648a33a7ed878a070d4f6251['h01ed0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f69] =  If409768b648a33a7ed878a070d4f6251['h01ed2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f6a] =  If409768b648a33a7ed878a070d4f6251['h01ed4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f6b] =  If409768b648a33a7ed878a070d4f6251['h01ed6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f6c] =  If409768b648a33a7ed878a070d4f6251['h01ed8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f6d] =  If409768b648a33a7ed878a070d4f6251['h01eda] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f6e] =  If409768b648a33a7ed878a070d4f6251['h01edc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f6f] =  If409768b648a33a7ed878a070d4f6251['h01ede] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f70] =  If409768b648a33a7ed878a070d4f6251['h01ee0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f71] =  If409768b648a33a7ed878a070d4f6251['h01ee2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f72] =  If409768b648a33a7ed878a070d4f6251['h01ee4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f73] =  If409768b648a33a7ed878a070d4f6251['h01ee6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f74] =  If409768b648a33a7ed878a070d4f6251['h01ee8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f75] =  If409768b648a33a7ed878a070d4f6251['h01eea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f76] =  If409768b648a33a7ed878a070d4f6251['h01eec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f77] =  If409768b648a33a7ed878a070d4f6251['h01eee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f78] =  If409768b648a33a7ed878a070d4f6251['h01ef0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f79] =  If409768b648a33a7ed878a070d4f6251['h01ef2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f7a] =  If409768b648a33a7ed878a070d4f6251['h01ef4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f7b] =  If409768b648a33a7ed878a070d4f6251['h01ef6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f7c] =  If409768b648a33a7ed878a070d4f6251['h01ef8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f7d] =  If409768b648a33a7ed878a070d4f6251['h01efa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f7e] =  If409768b648a33a7ed878a070d4f6251['h01efc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f7f] =  If409768b648a33a7ed878a070d4f6251['h01efe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f80] =  If409768b648a33a7ed878a070d4f6251['h01f00] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f81] =  If409768b648a33a7ed878a070d4f6251['h01f02] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f82] =  If409768b648a33a7ed878a070d4f6251['h01f04] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f83] =  If409768b648a33a7ed878a070d4f6251['h01f06] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f84] =  If409768b648a33a7ed878a070d4f6251['h01f08] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f85] =  If409768b648a33a7ed878a070d4f6251['h01f0a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f86] =  If409768b648a33a7ed878a070d4f6251['h01f0c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f87] =  If409768b648a33a7ed878a070d4f6251['h01f0e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f88] =  If409768b648a33a7ed878a070d4f6251['h01f10] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f89] =  If409768b648a33a7ed878a070d4f6251['h01f12] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f8a] =  If409768b648a33a7ed878a070d4f6251['h01f14] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f8b] =  If409768b648a33a7ed878a070d4f6251['h01f16] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f8c] =  If409768b648a33a7ed878a070d4f6251['h01f18] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f8d] =  If409768b648a33a7ed878a070d4f6251['h01f1a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f8e] =  If409768b648a33a7ed878a070d4f6251['h01f1c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f8f] =  If409768b648a33a7ed878a070d4f6251['h01f1e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f90] =  If409768b648a33a7ed878a070d4f6251['h01f20] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f91] =  If409768b648a33a7ed878a070d4f6251['h01f22] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f92] =  If409768b648a33a7ed878a070d4f6251['h01f24] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f93] =  If409768b648a33a7ed878a070d4f6251['h01f26] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f94] =  If409768b648a33a7ed878a070d4f6251['h01f28] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f95] =  If409768b648a33a7ed878a070d4f6251['h01f2a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f96] =  If409768b648a33a7ed878a070d4f6251['h01f2c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f97] =  If409768b648a33a7ed878a070d4f6251['h01f2e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f98] =  If409768b648a33a7ed878a070d4f6251['h01f30] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f99] =  If409768b648a33a7ed878a070d4f6251['h01f32] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f9a] =  If409768b648a33a7ed878a070d4f6251['h01f34] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f9b] =  If409768b648a33a7ed878a070d4f6251['h01f36] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f9c] =  If409768b648a33a7ed878a070d4f6251['h01f38] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f9d] =  If409768b648a33a7ed878a070d4f6251['h01f3a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f9e] =  If409768b648a33a7ed878a070d4f6251['h01f3c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00f9f] =  If409768b648a33a7ed878a070d4f6251['h01f3e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fa0] =  If409768b648a33a7ed878a070d4f6251['h01f40] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fa1] =  If409768b648a33a7ed878a070d4f6251['h01f42] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fa2] =  If409768b648a33a7ed878a070d4f6251['h01f44] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fa3] =  If409768b648a33a7ed878a070d4f6251['h01f46] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fa4] =  If409768b648a33a7ed878a070d4f6251['h01f48] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fa5] =  If409768b648a33a7ed878a070d4f6251['h01f4a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fa6] =  If409768b648a33a7ed878a070d4f6251['h01f4c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fa7] =  If409768b648a33a7ed878a070d4f6251['h01f4e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fa8] =  If409768b648a33a7ed878a070d4f6251['h01f50] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fa9] =  If409768b648a33a7ed878a070d4f6251['h01f52] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00faa] =  If409768b648a33a7ed878a070d4f6251['h01f54] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fab] =  If409768b648a33a7ed878a070d4f6251['h01f56] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fac] =  If409768b648a33a7ed878a070d4f6251['h01f58] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fad] =  If409768b648a33a7ed878a070d4f6251['h01f5a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fae] =  If409768b648a33a7ed878a070d4f6251['h01f5c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00faf] =  If409768b648a33a7ed878a070d4f6251['h01f5e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fb0] =  If409768b648a33a7ed878a070d4f6251['h01f60] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fb1] =  If409768b648a33a7ed878a070d4f6251['h01f62] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fb2] =  If409768b648a33a7ed878a070d4f6251['h01f64] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fb3] =  If409768b648a33a7ed878a070d4f6251['h01f66] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fb4] =  If409768b648a33a7ed878a070d4f6251['h01f68] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fb5] =  If409768b648a33a7ed878a070d4f6251['h01f6a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fb6] =  If409768b648a33a7ed878a070d4f6251['h01f6c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fb7] =  If409768b648a33a7ed878a070d4f6251['h01f6e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fb8] =  If409768b648a33a7ed878a070d4f6251['h01f70] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fb9] =  If409768b648a33a7ed878a070d4f6251['h01f72] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fba] =  If409768b648a33a7ed878a070d4f6251['h01f74] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fbb] =  If409768b648a33a7ed878a070d4f6251['h01f76] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fbc] =  If409768b648a33a7ed878a070d4f6251['h01f78] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fbd] =  If409768b648a33a7ed878a070d4f6251['h01f7a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fbe] =  If409768b648a33a7ed878a070d4f6251['h01f7c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fbf] =  If409768b648a33a7ed878a070d4f6251['h01f7e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fc0] =  If409768b648a33a7ed878a070d4f6251['h01f80] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fc1] =  If409768b648a33a7ed878a070d4f6251['h01f82] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fc2] =  If409768b648a33a7ed878a070d4f6251['h01f84] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fc3] =  If409768b648a33a7ed878a070d4f6251['h01f86] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fc4] =  If409768b648a33a7ed878a070d4f6251['h01f88] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fc5] =  If409768b648a33a7ed878a070d4f6251['h01f8a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fc6] =  If409768b648a33a7ed878a070d4f6251['h01f8c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fc7] =  If409768b648a33a7ed878a070d4f6251['h01f8e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fc8] =  If409768b648a33a7ed878a070d4f6251['h01f90] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fc9] =  If409768b648a33a7ed878a070d4f6251['h01f92] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fca] =  If409768b648a33a7ed878a070d4f6251['h01f94] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fcb] =  If409768b648a33a7ed878a070d4f6251['h01f96] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fcc] =  If409768b648a33a7ed878a070d4f6251['h01f98] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fcd] =  If409768b648a33a7ed878a070d4f6251['h01f9a] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fce] =  If409768b648a33a7ed878a070d4f6251['h01f9c] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fcf] =  If409768b648a33a7ed878a070d4f6251['h01f9e] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fd0] =  If409768b648a33a7ed878a070d4f6251['h01fa0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fd1] =  If409768b648a33a7ed878a070d4f6251['h01fa2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fd2] =  If409768b648a33a7ed878a070d4f6251['h01fa4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fd3] =  If409768b648a33a7ed878a070d4f6251['h01fa6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fd4] =  If409768b648a33a7ed878a070d4f6251['h01fa8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fd5] =  If409768b648a33a7ed878a070d4f6251['h01faa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fd6] =  If409768b648a33a7ed878a070d4f6251['h01fac] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fd7] =  If409768b648a33a7ed878a070d4f6251['h01fae] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fd8] =  If409768b648a33a7ed878a070d4f6251['h01fb0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fd9] =  If409768b648a33a7ed878a070d4f6251['h01fb2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fda] =  If409768b648a33a7ed878a070d4f6251['h01fb4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fdb] =  If409768b648a33a7ed878a070d4f6251['h01fb6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fdc] =  If409768b648a33a7ed878a070d4f6251['h01fb8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fdd] =  If409768b648a33a7ed878a070d4f6251['h01fba] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fde] =  If409768b648a33a7ed878a070d4f6251['h01fbc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fdf] =  If409768b648a33a7ed878a070d4f6251['h01fbe] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fe0] =  If409768b648a33a7ed878a070d4f6251['h01fc0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fe1] =  If409768b648a33a7ed878a070d4f6251['h01fc2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fe2] =  If409768b648a33a7ed878a070d4f6251['h01fc4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fe3] =  If409768b648a33a7ed878a070d4f6251['h01fc6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fe4] =  If409768b648a33a7ed878a070d4f6251['h01fc8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fe5] =  If409768b648a33a7ed878a070d4f6251['h01fca] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fe6] =  If409768b648a33a7ed878a070d4f6251['h01fcc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fe7] =  If409768b648a33a7ed878a070d4f6251['h01fce] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fe8] =  If409768b648a33a7ed878a070d4f6251['h01fd0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fe9] =  If409768b648a33a7ed878a070d4f6251['h01fd2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fea] =  If409768b648a33a7ed878a070d4f6251['h01fd4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00feb] =  If409768b648a33a7ed878a070d4f6251['h01fd6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fec] =  If409768b648a33a7ed878a070d4f6251['h01fd8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fed] =  If409768b648a33a7ed878a070d4f6251['h01fda] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fee] =  If409768b648a33a7ed878a070d4f6251['h01fdc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fef] =  If409768b648a33a7ed878a070d4f6251['h01fde] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ff0] =  If409768b648a33a7ed878a070d4f6251['h01fe0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ff1] =  If409768b648a33a7ed878a070d4f6251['h01fe2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ff2] =  If409768b648a33a7ed878a070d4f6251['h01fe4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ff3] =  If409768b648a33a7ed878a070d4f6251['h01fe6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ff4] =  If409768b648a33a7ed878a070d4f6251['h01fe8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ff5] =  If409768b648a33a7ed878a070d4f6251['h01fea] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ff6] =  If409768b648a33a7ed878a070d4f6251['h01fec] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ff7] =  If409768b648a33a7ed878a070d4f6251['h01fee] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ff8] =  If409768b648a33a7ed878a070d4f6251['h01ff0] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ff9] =  If409768b648a33a7ed878a070d4f6251['h01ff2] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ffa] =  If409768b648a33a7ed878a070d4f6251['h01ff4] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ffb] =  If409768b648a33a7ed878a070d4f6251['h01ff6] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ffc] =  If409768b648a33a7ed878a070d4f6251['h01ff8] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ffd] =  If409768b648a33a7ed878a070d4f6251['h01ffa] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00ffe] =  If409768b648a33a7ed878a070d4f6251['h01ffc] ;
//end
//always_comb begin // 
               Ic8a4ab93493bd6cdd4939054e46d2247['h00fff] =  If409768b648a33a7ed878a070d4f6251['h01ffe] ;
//end
