 reg  ['h0:0] [$clog2('h7000+1)-1:0] I5edb7954620e8b8032a9ad41b528b90c9fbed81d94a9becd64145bb694902376 ;
